
-- Copyright (C) 2010 David E. Roberts <davee dot roberts at fsmail dot net>

-- This file is part of AGCNORM (Apollo Guidance Computer NOR eMulator).
--
-- AGCNORM is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- AGCNORM is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with AGCNORM. If not, see <http://www.gnu.org/licenses/>.

-- Functional description.
-- =======================
--
-- This file implements the NOR gate logic of the Block II Apollo Guidance Computer (AGC)
-- as published at <http://klabs.org/history/ech/agc_schematics> with some
-- minor modifications by the author to enable the logic to operate within the hardware of
-- a Field Programmable Gate Array (FPGA). The logic is implemented as a VHDL description
-- for a Xilinx Spartan 3E device (XC3S500E-FG320-4) using release 11.1 of the ISE WebPACK tools.

-- Modification History.
-- =====================
--
-- Version : 
--    Date : 
--  Author : 
--  Reason : 
--
-- Version : 2.06
--    Date : 14th August 2010
--  Author : David E. Roberts
--  Reason : Change from LED/SWITCH debug of the Hydra-XC to a VGA debug for the Spartan 3E Starter Kit.
--         : Small changes to the signals used for debugging.
--         : Remove NHALGA hack from CH77.
--
-- Version : 2.03
--    Date : 11th April 2010
--  Author : David E. Roberts
--  Reason : Add FS01..FS33 to the DEBUG LEDS. FS01..FS20 assigned to X08 and FS21..FS33 assigned to X09.
--
-- Version : 2.02
--    Date : 10th April 2010
--  Author : David E. Roberts
--  Reason : Increase the number of DEBUG LEDS from 16 to 20 and increase the number of
--           DEBUG SWITCHES from 4 to 8.
--
-- Version : 2.01
--    Date : 20th March 2010
--  Author : David E. Roberts
--  Reason : Add DEBSWS.
--
-- Version : 2.00
--    Date : 18th March 2010
--  Author : David E. Roberts
--  Reason : Major re-write using instantiations of LUT4_L and FDRSE elements.
--
-- Version : 1.08
--    Date : 14th February 2010
--  Author : David E. Roberts
--  Reason : Remove combinatorial loop formed on A2/3 from 37343 -> 37346 -> 37348. Resolve by making
--           gates 37345 and 37346 into latches (NORX) with an initial value of '0'.
--
-- Version : 1.07
--    Date : 13th February 2010
--  Author : David E. Roberts
--  Reason : Add DEBLEDS. Convert some more NORX/NORX flip-flops to NORX/NORY.
--
-- Version : 1.06
--    Date : 27th January 2010
--  Author : David E. Roberts
--  Reason : Change A23/1 gate 48258 from T7PH??? to T7PHS4 and remove PULLU150 from CH77. I believe
--           the expander gate 48258 on A23/1 is an inhibit for T7PHS4 on A23/2. It doesn't make sense
--           for 48258 to be T7PHS4/ as this will leave T7PHS4 clocking away whilst stopping the inverse
--           clock - not sensible to me.
--         : Don't forget to keep changing the NORX/NORX flip-flops to NORX/NORY ones as in the comment
--           associated with Version 1.05...
--
-- Version : 1.05
--    Date : 27th January 2010
--  Author : David E. Roberts
--  Reason : Problem found with CH77 RESTART MONITOR logic. My cross-coupled NOR flip flops consisted
--           of cross-coupled latches to overcome the problem with the VHDL synthesis of trying to
--           resolve closed loop feedback paths - which the tool didn't like! I have a one-SYSCLOCK
--           wide pulse on MPAL/ (for some reason) which is causing my F/F implementation to oscillate.
--           Checking this by hand seems to indicate that this behaviour is correct - but not desired!
--           To overcome this problem, I am replacing the two cross-coupled latches (NORX, NORX) with a
--           latch (NORX) and a gate (NORY). I have tested this with CH77 and found it to work fine. This
--           needs replicating throughout the entire design... The choice of which latch is turned into
--           a gate is a little arbitary at the moment - but I am going with the CLEAR/RESET side as the
--           gate (NORY) with the SET side as the latch (NORX) element.
--
-- Version : 1.04
--    Date : 23rd January 2010
--  Author : David E. Roberts
--  Reason : Change the way I/O is handled. Revert back to a record structure passed from/to
--           the parent module.
--
-- Version : 1.03
--    Date : 22nd January 2010
--  Author : David E. Roberts
--  Reason : Resolve mess up with deriving SYSERROR from channel 77 alarms.
--
-- Version : 1.02
--    Date : 14th January 2010
--  Author : David E. Roberts
--  Reason : Gates 37139, 37140 and 37142 on A2/1 changed from sequential to combinatorial logic.
--           The DAS instruction was trying to test for overflow/underflow using the control
--           pulse TOV/ to latch UNF/ and OVF/ into BR1 and BR2 respectively on diagram A4/1.
--           Unfortunately, UNF/ and OVF/ are only valid when OVFSTB/ is active (A2/3).
--           OVFSTB/ is generated on A2/1 from CT/ which is in turn derived from the four-phase
--           clock generator. I suspect that delaying the clock signal through the identified
--           gates delays CT/ which in turn delays OVFSTB/ too much so that it is active once
--           TOV/ has become inactive! I suspect that these three gates were included in the
--           original design to delay signal CT/ to compensate for the delays through the
--           STAGE BRANCH DECODER and CROSS POINT GENERATOR which doesn't happen much in the
--           FPGA design. Removing these three effective gate delays will (hopefully) cause
--           OVFSTB/ to validly occur within the TOV/ window and will not cause any unforseen
--           problems to occur.
--
-- Version : 1.01
--    Date : 1st January 2010
--  Author : David E. Roberts
--  Reason : Changed input #1 of gates 41125 and 41126 of A13/1 from F10A to F10A/.
--           I believe this is necessary to stop the error MTCAL/ (TC Trap) from occuring.
--           I suspect that the original used F10A/ or used F10A with an on-board inverter
--           gate which has not been shown.
--
-- Version : 1.00
--    Date : 29th December 2009
--  Author : David E. Roberts
--  Reason : First creation

-- Known issues.
-- =============
--
-- There are some connector names that have been difficult to read from the schematic diagrams.
-- I have made my 'best guess'.
--
-- SYSERROR is raised because of a problem with signal MSCDBL/.

-- Automatically generated at 14:28:39 on 14/08/2010 

-- Error count was 0 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.AGCPACK.all;

package AGCIO is

  -- **********************************
  -- ***                            ***
  -- ***  INPUT record descriptor.  ***
  -- ***                            ***
  -- **********************************

  type t_INPUTS is
  record
    \NHVFAL\    : AGCBIT;
    \MAINRS\    : AGCBIT;
    \SBYBUT\    : AGCBIT;
    \IN3212\    : AGCBIT;
    \CAURST\    : AGCBIT;
    \IN3213\    : AGCBIT;
    \NKEY1\     : AGCBIT;
    \IN3214\    : AGCBIT;
    \NKEY2\     : AGCBIT;
    \MKEY1\     : AGCBIT;
    \NKEY3\     : AGCBIT;
    \MKEY2\     : AGCBIT;
    \NKEY4\     : AGCBIT;
    \MKEY3\     : AGCBIT;
    \NKEY5\     : AGCBIT;
    \MKEY4\     : AGCBIT;
    \NAVRST\    : AGCBIT;
    \MKEY5\     : AGCBIT;
    \IN3216\    : AGCBIT;
    \GATEX/\    : AGCBIT;
    \GATEY/\    : AGCBIT;
    \GATEZ/\    : AGCBIT;
    \SIGNX\     : AGCBIT;
    \SIGNY\     : AGCBIT;
    \SIGNZ\     : AGCBIT;
    \BMGXP\     : AGCBIT;
    \CDUXM\     : AGCBIT;
    \DKSTRT\    : AGCBIT;
    \BMGXM\     : AGCBIT;
    \CDUYP\     : AGCBIT;
    \DKEND\     : AGCBIT;
    \BMGYP\     : AGCBIT;
    \CDUYM\     : AGCBIT;
    \DKBSNC\    : AGCBIT;
    \BMGYM\     : AGCBIT;
    \CDUZP\     : AGCBIT;
    \UPL0\      : AGCBIT;
    \BMGZP\     : AGCBIT;
    \CDUZM\     : AGCBIT;
    \UPL1\      : AGCBIT;
    \BMGZM\     : AGCBIT;
    \PIPAX+\    : AGCBIT;
    \RRIN0\     : AGCBIT;
    \SHAFTP\    : AGCBIT;
    \PIPAX-\    : AGCBIT;
    \RRIN1\     : AGCBIT;
    \SHAFTM\    : AGCBIT;
    \PIPAY+\    : AGCBIT;
    \LRIN0\     : AGCBIT;
    \TRNP\      : AGCBIT;
    \PIPAY-\    : AGCBIT;
    \LRIN1\     : AGCBIT;
    \TRNM\      : AGCBIT;
    \PIPAZ+\    : AGCBIT;
    \XLNK0\     : AGCBIT;
    \CDUXP\     : AGCBIT;
    \PIPAZ-\    : AGCBIT;
    \XLNK1\     : AGCBIT;
    \ULLTHR\    : AGCBIT;
    \MNIM+Y\    : AGCBIT;
    \RRPONA\    : AGCBIT;
    \LFTOFF\    : AGCBIT;
    \MNIM-Y\    : AGCBIT;
    \RRRLSC\    : AGCBIT;
    \GUIREL\    : AGCBIT;
    \MNIM+R\    : AGCBIT;
    \MANR+P\    : AGCBIT;
    \TRAN+X\    : AGCBIT;
    \MNIM-R\    : AGCBIT;
    \MANR-P\    : AGCBIT;
    \TRAN-X\    : AGCBIT;
    \TRST9\     : AGCBIT;
    \MANR+Y\    : AGCBIT;
    \TRAN+Y\    : AGCBIT;
    \TRST10\    : AGCBIT;
    \MANR-Y\    : AGCBIT;
    \TRAN-Y\    : AGCBIT;
    \HOLFUN\    : AGCBIT;
    \MANR+R\    : AGCBIT;
    \TRAN+Z\    : AGCBIT;
    \FREFUN\    : AGCBIT;
    \MANR-R\    : AGCBIT;
    \TRAN-Z\    : AGCBIT;
    \S4BSAB\    : AGCBIT;
    \ISSTOR\    : AGCBIT;
    \OPCDFL\    : AGCBIT;
    \SMSEPR\    : AGCBIT;
    \OPCDEL\    : AGCBIT;
    \MRKRST\    : AGCBIT;
    \IN3008\    : AGCBIT;
    \CDUFAL\    : AGCBIT;
    \ZEROP\     : AGCBIT;
    \BLKUPL/\   : AGCBIT;
    \TEMPIN\    : AGCBIT;
    \MARK\      : AGCBIT;
    \SPSRDY\    : AGCBIT;
    \IMUFAL\    : AGCBIT;
    \OPMSW3\    : AGCBIT;
    \GCAPCL\    : AGCBIT;
    \LEMATT\    : AGCBIT;
    \MRKREJ\    : AGCBIT;
    \ROLGOF\    : AGCBIT;
    \IMUOPR\    : AGCBIT;
    \STRPRS\    : AGCBIT;
    \PCHGOF\    : AGCBIT;
    \IMUCAG\    : AGCBIT;
    \MNIM+P\    : AGCBIT;
    \LVDAGD\    : AGCBIT;
    \IN3301\    : AGCBIT;
    \MNIM-P\    : AGCBIT;
    \LRRLSC\    : AGCBIT;
    \CTLSAT\    : AGCBIT;
    \2FSFAL\    : AGCBIT;
    \FLTOUT\    : AGCBIT;
    \OPMSW2\    : AGCBIT;
    \SCAFAL\    : AGCBIT;
    \STRT2\     : AGCBIT;
    \VFAIL\     : AGCBIT;
  end record; -- t_INPUTS

  -- ***********************************
  -- ***                             ***
  -- ***  OUTPUT record descriptor.  ***
  -- ***                             ***
  -- ***********************************

  type t_OUTPUTS is
  record
    \3200A\     : AGCBIT;
    \CDUXDP\    : AGCBIT;
    \3200B\     : AGCBIT;
    \CDUXDM\    : AGCBIT;
    \3200C\     : AGCBIT;
    \CDUYDP\    : AGCBIT;
    \3200D\     : AGCBIT;
    \CDUYDM\    : AGCBIT;
    \25KPPS\    : AGCBIT;
    \CDUCLK\    : AGCBIT;
    \12KPPS\    : AGCBIT;
    \PIPINT\    : AGCBIT;
    \800SET\    : AGCBIT;
    \PIPASW\    : AGCBIT;
    \800RST\    : AGCBIT;
    \PIPDAT\    : AGCBIT;
    \GYENAB\    : AGCBIT;
    \CLK\       : AGCBIT;
    \CDUZDP\    : AGCBIT;
    \RRRST\     : AGCBIT;
    \CDUZDM\    : AGCBIT;
    \LRRST\     : AGCBIT;
    \OT1114\    : AGCBIT;
    \RC-X+P\    : AGCBIT;
    \OT1113\    : AGCBIT;
    \RC+X-Y\    : AGCBIT;
    \OT1112\    : AGCBIT;
    \RC+X+Y\    : AGCBIT;
    \OT1111\    : AGCBIT;
    \RC+X-P\    : AGCBIT;
    \OT1110\    : AGCBIT;
    \RC+X+P\    : AGCBIT;
    \OT1108\    : AGCBIT;
    \TMPCAU\    : AGCBIT;
    \OPEROR\    : AGCBIT;
    \ISSTDC\    : AGCBIT;
    \ELSNCM\    : AGCBIT;
    \OT1116\    : AGCBIT;
    \VNFLSH\    : AGCBIT;
    \ENERIM\    : AGCBIT;
    \CGCWAR\    : AGCBIT;
    \ZIMCDU\    : AGCBIT;
    \KYRLS\     : AGCBIT;
    \COARSE\    : AGCBIT;
    \UPLACT\    : AGCBIT;
    \ENEROP\    : AGCBIT;
    \S4BOFF\    : AGCBIT;
    \ZEROPT\    : AGCBIT;
    \S4BSEQ\    : AGCBIT;
    \MROLGT\    : AGCBIT;
    \RESTRT\    : AGCBIT;
    \ZOPCDU\    : AGCBIT;
    \SBYLIT\    : AGCBIT;
    \ALTSNC\    : AGCBIT;
    \COMACT\    : AGCBIT;
    \OT1207/\   : AGCBIT;
    \ISSWAR\    : AGCBIT;
    \OT1207\    : AGCBIT;
    \RYWD16\    : AGCBIT;
    \S4BTAK\    : AGCBIT;
    \RYWD14\    : AGCBIT;
    \DISDAC\    : AGCBIT;
    \RYWD13\    : AGCBIT;
    \STARON\    : AGCBIT;
    \RYWD12\    : AGCBIT;
    \TVCNAB\    : AGCBIT;
    \RLYB11\    : AGCBIT;
    \RC-Z-R\    : AGCBIT;
    \RLYB10\    : AGCBIT;
    \RC-Z+R\    : AGCBIT;
    \RLYB09\    : AGCBIT;
    \RC+Z-R\    : AGCBIT;
    \RLYB08\    : AGCBIT;
    \RC+Z+R\    : AGCBIT;
    \RLYB07\    : AGCBIT;
    \RC-Y-R\    : AGCBIT;
    \RLYB06\    : AGCBIT;
    \RC-Y+R\    : AGCBIT;
    \RLYB05\    : AGCBIT;
    \RC+Y-R\    : AGCBIT;
    \RLYB04\    : AGCBIT;
    \RC+Y+R\    : AGCBIT;
    \RLYB03\    : AGCBIT;
    \RC-X-Y\    : AGCBIT;
    \RLYB02\    : AGCBIT;
    \RC-X+Y\    : AGCBIT;
    \RLYB01\    : AGCBIT;
    \RC-X-P\    : AGCBIT;
    \ELSNCN\    : AGCBIT;
    \THRST+\    : AGCBIT;
    \LRRANG\    : AGCBIT;
    \SHFTDP\    : AGCBIT;
    \THRST-\    : AGCBIT;
    \LRZVEL\    : AGCBIT;
    \SHFTDM\    : AGCBIT;
    \EMS+\      : AGCBIT;
    \LRYVEL\    : AGCBIT;
    \TRNDP\     : AGCBIT;
    \EMS-\      : AGCBIT;
    \LRXVEL\    : AGCBIT;
    \TRNDM\     : AGCBIT;
    \ALT1\      : AGCBIT;
    \RRRANG\    : AGCBIT;
    \GYRSET\    : AGCBIT;
    \ALT0\      : AGCBIT;
    \RRRARA\    : AGCBIT;
    \GYRRST\    : AGCBIT;
    \ALRT1\     : AGCBIT;
    \RRSYNC\    : AGCBIT;
    \OTLNK0\    : AGCBIT;
    \ALRT0\     : AGCBIT;
    \LRSYNC\    : AGCBIT;
    \OTLNK1\    : AGCBIT;
    \DKDATB\    : AGCBIT;
    \DKDATA\    : AGCBIT;
    \GYZM\      : AGCBIT;
    \GYYM\      : AGCBIT;
    \GYXM\      : AGCBIT;
    \GYZP\      : AGCBIT;
    \GYYP\      : AGCBIT;
    \GYXP\      : AGCBIT;
  end record; -- t_OUTPUTS

end AGCIO;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library UNISIM;
use UNISIM.VComponents.all;

use work.AGCPACK.all;
use work.AGCIO.all;

entity AGC_LOGIC is
  port(
    SYSCLOCK  : in  AGCBIT;
    SYSRESET  : in  AGCBIT;
    SYSERROR  : out AGCBIT;
    \CLOCK\   : in  AGCBIT;
    ECADR     : out AGCBITARRAY( 11 downto 1 );
    FCADR     : out AGCBITARRAY( 16 downto 1 );
    SAXX      : in  AGCBITARRAY( 15 downto 0 );
    GEMXX     : out AGCBITARRAY( 15 downto 0 );
    EWRITE    : out AGCBIT;
    EREAD     : out AGCBIT;
    ESTART    : out AGCBIT;
    FREAD     : out AGCBIT;
    INPUTS    : in  t_INPUTS;
    OUTPUTS   : out t_OUTPUTS;
    VGADEBUG  : out t_debug
  );
end AGC_LOGIC;

architecture Rtl of AGC_LOGIC is

  -- ************************************
  -- ***                              ***
  -- ***  INPUT signal declarations.  ***
  -- ***                              ***
  -- ************************************

  signal \SAP\      : AGCBIT;
  signal \SA01\     : AGCBIT;
  signal \SA02\     : AGCBIT;
  signal \SA03\     : AGCBIT;
  signal \SA04\     : AGCBIT;
  signal \SA05\     : AGCBIT;
  signal \SA06\     : AGCBIT;
  signal \SA07\     : AGCBIT;
  signal \SA08\     : AGCBIT;
  signal \SA09\     : AGCBIT;
  signal \SA10\     : AGCBIT;
  signal \SA11\     : AGCBIT;
  signal \SA12\     : AGCBIT;
  signal \SA13\     : AGCBIT;
  signal \SA14\     : AGCBIT;
  signal \SA16\     : AGCBIT;

  signal \NHVFAL\    : AGCBIT;
  signal \MAINRS\    : AGCBIT;
  signal \SBYBUT\    : AGCBIT;
  signal \IN3212\    : AGCBIT;
  signal \CAURST\    : AGCBIT;
  signal \IN3213\    : AGCBIT;
  signal \NKEY1\     : AGCBIT;
  signal \IN3214\    : AGCBIT;
  signal \NKEY2\     : AGCBIT;
  signal \MKEY1\     : AGCBIT;
  signal \NKEY3\     : AGCBIT;
  signal \MKEY2\     : AGCBIT;
  signal \NKEY4\     : AGCBIT;
  signal \MKEY3\     : AGCBIT;
  signal \NKEY5\     : AGCBIT;
  signal \MKEY4\     : AGCBIT;
  signal \NAVRST\    : AGCBIT;
  signal \MKEY5\     : AGCBIT;
  signal \IN3216\    : AGCBIT;
  signal \GATEX/\    : AGCBIT;
  signal \GATEY/\    : AGCBIT;
  signal \GATEZ/\    : AGCBIT;
  signal \SIGNX\     : AGCBIT;
  signal \SIGNY\     : AGCBIT;
  signal \SIGNZ\     : AGCBIT;
  signal \BMGXP\     : AGCBIT;
  signal \CDUXM\     : AGCBIT;
  signal \DKSTRT\    : AGCBIT;
  signal \BMGXM\     : AGCBIT;
  signal \CDUYP\     : AGCBIT;
  signal \DKEND\     : AGCBIT;
  signal \BMGYP\     : AGCBIT;
  signal \CDUYM\     : AGCBIT;
  signal \DKBSNC\    : AGCBIT;
  signal \BMGYM\     : AGCBIT;
  signal \CDUZP\     : AGCBIT;
  signal \UPL0\      : AGCBIT;
  signal \BMGZP\     : AGCBIT;
  signal \CDUZM\     : AGCBIT;
  signal \UPL1\      : AGCBIT;
  signal \BMGZM\     : AGCBIT;
  signal \PIPAX+\    : AGCBIT;
  signal \RRIN0\     : AGCBIT;
  signal \SHAFTP\    : AGCBIT;
  signal \PIPAX-\    : AGCBIT;
  signal \RRIN1\     : AGCBIT;
  signal \SHAFTM\    : AGCBIT;
  signal \PIPAY+\    : AGCBIT;
  signal \LRIN0\     : AGCBIT;
  signal \TRNP\      : AGCBIT;
  signal \PIPAY-\    : AGCBIT;
  signal \LRIN1\     : AGCBIT;
  signal \TRNM\      : AGCBIT;
  signal \PIPAZ+\    : AGCBIT;
  signal \XLNK0\     : AGCBIT;
  signal \CDUXP\     : AGCBIT;
  signal \PIPAZ-\    : AGCBIT;
  signal \XLNK1\     : AGCBIT;
  signal \ULLTHR\    : AGCBIT;
  signal \MNIM+Y\    : AGCBIT;
  signal \RRPONA\    : AGCBIT;
  signal \LFTOFF\    : AGCBIT;
  signal \MNIM-Y\    : AGCBIT;
  signal \RRRLSC\    : AGCBIT;
  signal \GUIREL\    : AGCBIT;
  signal \MNIM+R\    : AGCBIT;
  signal \MANR+P\    : AGCBIT;
  signal \TRAN+X\    : AGCBIT;
  signal \MNIM-R\    : AGCBIT;
  signal \MANR-P\    : AGCBIT;
  signal \TRAN-X\    : AGCBIT;
  signal \TRST9\     : AGCBIT;
  signal \MANR+Y\    : AGCBIT;
  signal \TRAN+Y\    : AGCBIT;
  signal \TRST10\    : AGCBIT;
  signal \MANR-Y\    : AGCBIT;
  signal \TRAN-Y\    : AGCBIT;
  signal \HOLFUN\    : AGCBIT;
  signal \MANR+R\    : AGCBIT;
  signal \TRAN+Z\    : AGCBIT;
  signal \FREFUN\    : AGCBIT;
  signal \MANR-R\    : AGCBIT;
  signal \TRAN-Z\    : AGCBIT;
  signal \S4BSAB\    : AGCBIT;
  signal \ISSTOR\    : AGCBIT;
  signal \OPCDFL\    : AGCBIT;
  signal \SMSEPR\    : AGCBIT;
  signal \OPCDEL\    : AGCBIT;
  signal \MRKRST\    : AGCBIT;
  signal \IN3008\    : AGCBIT;
  signal \CDUFAL\    : AGCBIT;
  signal \ZEROP\     : AGCBIT;
  signal \BLKUPL/\   : AGCBIT;
  signal \TEMPIN\    : AGCBIT;
  signal \MARK\      : AGCBIT;
  signal \SPSRDY\    : AGCBIT;
  signal \IMUFAL\    : AGCBIT;
  signal \OPMSW3\    : AGCBIT;
  signal \GCAPCL\    : AGCBIT;
  signal \LEMATT\    : AGCBIT;
  signal \MRKREJ\    : AGCBIT;
  signal \ROLGOF\    : AGCBIT;
  signal \IMUOPR\    : AGCBIT;
  signal \STRPRS\    : AGCBIT;
  signal \PCHGOF\    : AGCBIT;
  signal \IMUCAG\    : AGCBIT;
  signal \MNIM+P\    : AGCBIT;
  signal \LVDAGD\    : AGCBIT;
  signal \IN3301\    : AGCBIT;
  signal \MNIM-P\    : AGCBIT;
  signal \LRRLSC\    : AGCBIT;
  signal \CTLSAT\    : AGCBIT;
  signal \2FSFAL\    : AGCBIT;
  signal \FLTOUT\    : AGCBIT;
  signal \OPMSW2\    : AGCBIT;
  signal \SCAFAL\    : AGCBIT;
  signal \STRT2\     : AGCBIT;
  signal \VFAIL\     : AGCBIT;

  -- ***********************************
  -- ***                             ***
  -- ***  Gate signal declarations.  ***
  -- ***                             ***
  -- ***********************************

  signal  \38101\    : AGCBIT; signal  \CHAT05\   : AGCBIT;
  signal  \38102\    : AGCBIT; signal  \F10A\     : AGCBIT;
  signal  \38103\    : AGCBIT;
  signal \$38103\    : AGCBIT;
  signal  \38104\    : AGCBIT;
  signal \$38104\    : AGCBIT;
  signal  \38105\    : AGCBIT;
  signal \$38105\    : AGCBIT;
  signal  \38106\    : AGCBIT; signal  \FS10\     : AGCBIT;
  signal  \38107\    : AGCBIT; signal  \F10B\     : AGCBIT;
  signal  \38111\    : AGCBIT; signal  \CHAT06\   : AGCBIT;
  signal  \38112\    : AGCBIT; signal  \F11A\     : AGCBIT;
  signal  \38113\    : AGCBIT;
  signal \$38113\    : AGCBIT;
  signal  \38114\    : AGCBIT;
  signal \$38114\    : AGCBIT;
  signal  \38115\    : AGCBIT;
  signal \$38115\    : AGCBIT;
  signal  \38116\    : AGCBIT; signal  \FS11\     : AGCBIT;
  signal  \38117\    : AGCBIT; signal  \F11B\     : AGCBIT;
  signal  \38121\    : AGCBIT; signal  \CHAT07\   : AGCBIT;
  signal  \38122\    : AGCBIT; signal  \F12A\     : AGCBIT;
  signal  \38123\    : AGCBIT;
  signal \$38123\    : AGCBIT;
  signal  \38124\    : AGCBIT;
  signal \$38124\    : AGCBIT;
  signal  \38125\    : AGCBIT;
  signal \$38125\    : AGCBIT;
  signal  \38126\    : AGCBIT; signal  \FS12\     : AGCBIT;
  signal  \38127\    : AGCBIT; signal  \F12B\     : AGCBIT;
  signal  \38131\    : AGCBIT; signal  \CHAT08\   : AGCBIT;
  signal  \38132\    : AGCBIT; signal  \F13A\     : AGCBIT;
  signal  \38133\    : AGCBIT;
  signal \$38133\    : AGCBIT;
  signal  \38134\    : AGCBIT;
  signal \$38134\    : AGCBIT;
  signal  \38135\    : AGCBIT;
  signal \$38135\    : AGCBIT;
  signal  \38136\    : AGCBIT; signal  \FS13\     : AGCBIT;
  signal  \38137\    : AGCBIT; signal  \F13B\     : AGCBIT;
  signal  \38141\    : AGCBIT; signal  \CHAT09\   : AGCBIT;
  signal  \38142\    : AGCBIT; signal  \F14A\     : AGCBIT;
  signal  \38143\    : AGCBIT;
  signal \$38143\    : AGCBIT;
  signal  \38144\    : AGCBIT;
  signal \$38144\    : AGCBIT;
  signal  \38145\    : AGCBIT;
  signal \$38145\    : AGCBIT;
  signal  \38146\    : AGCBIT; signal  \FS14\     : AGCBIT;
  signal  \38147\    : AGCBIT; signal  \F14B\     : AGCBIT;
  signal  \38151\    : AGCBIT; signal  \CHAT10\   : AGCBIT;
  signal  \38152\    : AGCBIT; signal  \F15A\     : AGCBIT;
  signal  \38153\    : AGCBIT;
  signal \$38153\    : AGCBIT;
  signal  \38154\    : AGCBIT;
  signal \$38154\    : AGCBIT;
  signal  \38155\    : AGCBIT;
  signal \$38155\    : AGCBIT;
  signal  \38156\    : AGCBIT; signal  \FS15\     : AGCBIT;
  signal  \38157\    : AGCBIT; signal  \F15B\     : AGCBIT;
  signal  \38161\    : AGCBIT; signal  \CHAT11\   : AGCBIT;
  signal  \38162\    : AGCBIT; signal  \F16A\     : AGCBIT;
  signal  \38163\    : AGCBIT;
  signal \$38163\    : AGCBIT;
  signal  \38164\    : AGCBIT;
  signal \$38164\    : AGCBIT;
  signal  \38165\    : AGCBIT;
  signal \$38165\    : AGCBIT;
  signal  \38166\    : AGCBIT; signal  \FS16\     : AGCBIT;
  signal  \38167\    : AGCBIT; signal  \F16B\     : AGCBIT;
  signal  \38171\    : AGCBIT; signal  \CHAT12\   : AGCBIT;
  signal  \38172\    : AGCBIT; signal  \F17A\     : AGCBIT;
  signal  \38173\    : AGCBIT;
  signal \$38173\    : AGCBIT;
  signal  \38174\    : AGCBIT;
  signal \$38174\    : AGCBIT;
  signal  \38175\    : AGCBIT;
  signal \$38175\    : AGCBIT;
  signal  \38176\    : AGCBIT; signal  \FS17\     : AGCBIT;
  signal  \38177\    : AGCBIT; signal  \F17B\     : AGCBIT;
  signal  \38190\    : AGCBIT; signal  \FS06/\    : AGCBIT;
  signal  \38191\    : AGCBIT; signal  \FS07/\    : AGCBIT;
  signal  \38201\    : AGCBIT; signal  \FS02A\    : AGCBIT;
  signal  \38202\    : AGCBIT; signal  \F02A\     : AGCBIT;
  signal  \38203\    : AGCBIT;
  signal \$38203\    : AGCBIT;
  signal  \38204\    : AGCBIT;
  signal \$38204\    : AGCBIT;
  signal  \38205\    : AGCBIT;
  signal \$38205\    : AGCBIT;
  signal  \38206\    : AGCBIT; signal  \FS02\     : AGCBIT;
  signal  \38207\    : AGCBIT; signal  \F02B\     : AGCBIT;
  signal  \38211\    : AGCBIT; signal  \FS03A\    : AGCBIT;
  signal  \38212\    : AGCBIT; signal  \F03A\     : AGCBIT;
  signal  \38213\    : AGCBIT;
  signal \$38213\    : AGCBIT;
  signal  \38214\    : AGCBIT;
  signal \$38214\    : AGCBIT;
  signal  \38215\    : AGCBIT;
  signal \$38215\    : AGCBIT;
  signal  \38216\    : AGCBIT; signal  \FS03\     : AGCBIT;
  signal  \38217\    : AGCBIT; signal  \F03B\     : AGCBIT;
  signal  \38221\    : AGCBIT; signal  \FS04A\    : AGCBIT;
  signal  \38222\    : AGCBIT; signal  \F04A\     : AGCBIT;
  signal  \38223\    : AGCBIT;
  signal \$38223\    : AGCBIT;
  signal  \38224\    : AGCBIT;
  signal \$38224\    : AGCBIT;
  signal  \38225\    : AGCBIT;
  signal \$38225\    : AGCBIT;
  signal  \38226\    : AGCBIT; signal  \FS04\     : AGCBIT;
  signal  \38227\    : AGCBIT; signal  \F04B\     : AGCBIT;
  signal  \38231\    : AGCBIT; signal  \FS05A\    : AGCBIT;
  signal  \38232\    : AGCBIT; signal  \F05A\     : AGCBIT;
  signal  \38233\    : AGCBIT;
  signal \$38233\    : AGCBIT;
  signal  \38234\    : AGCBIT;
  signal \$38234\    : AGCBIT;
  signal  \38235\    : AGCBIT;
  signal \$38235\    : AGCBIT;
  signal  \38236\    : AGCBIT; signal  \FS05\     : AGCBIT;
  signal  \38237\    : AGCBIT; signal  \F05B\     : AGCBIT;
  signal  \38241\    : AGCBIT; signal  \CHAT01\   : AGCBIT;
  signal  \38242\    : AGCBIT; signal  \F06A\     : AGCBIT;
  signal  \38243\    : AGCBIT;
  signal \$38243\    : AGCBIT;
  signal  \38244\    : AGCBIT;
  signal \$38244\    : AGCBIT;
  signal  \38245\    : AGCBIT;
  signal \$38245\    : AGCBIT;
  signal  \38246\    : AGCBIT; signal  \FS06\     : AGCBIT;
  signal  \38247\    : AGCBIT; signal  \F06B\     : AGCBIT;
  signal  \38251\    : AGCBIT; signal  \CHAT02\   : AGCBIT;
  signal  \38252\    : AGCBIT; signal  \F07A\     : AGCBIT;
  signal  \38253\    : AGCBIT;
  signal \$38253\    : AGCBIT;
  signal  \38254\    : AGCBIT;
  signal \$38254\    : AGCBIT;
  signal  \38255\    : AGCBIT;
  signal \$38255\    : AGCBIT;
  signal  \38256\    : AGCBIT; signal  \FS07\     : AGCBIT;
  signal  \38257\    : AGCBIT; signal  \F07B\     : AGCBIT;
  signal  \38261\    : AGCBIT; signal  \CHAT03\   : AGCBIT;
  signal  \38262\    : AGCBIT; signal  \F08A\     : AGCBIT;
  signal  \38263\    : AGCBIT;
  signal \$38263\    : AGCBIT;
  signal  \38264\    : AGCBIT;
  signal \$38264\    : AGCBIT;
  signal  \38265\    : AGCBIT;
  signal \$38265\    : AGCBIT;
  signal  \38266\    : AGCBIT; signal  \FS08\     : AGCBIT;
  signal  \38267\    : AGCBIT; signal  \F08B\     : AGCBIT;
  signal  \38271\    : AGCBIT; signal  \CHAT04\   : AGCBIT;
  signal  \38272\    : AGCBIT; signal  \F09A\     : AGCBIT;
  signal  \38273\    : AGCBIT;
  signal \$38273\    : AGCBIT;
  signal  \38274\    : AGCBIT;
  signal \$38274\    : AGCBIT;
  signal  \38275\    : AGCBIT;
  signal \$38275\    : AGCBIT;
  signal  \38276\    : AGCBIT; signal  \FS09\     : AGCBIT;
  signal  \38277\    : AGCBIT; signal  \F09B\     : AGCBIT;
  signal  \38290\    : AGCBIT; signal  \FS08/\    : AGCBIT;
  signal  \38291\    : AGCBIT; signal  \FS07A\    : AGCBIT;
  signal  \38301\    : AGCBIT; signal  \CHAT13\   : AGCBIT;
  signal  \38302\    : AGCBIT; signal  \F18A\     : AGCBIT;
  signal  \38303\    : AGCBIT;
  signal \$38303\    : AGCBIT;
  signal  \38304\    : AGCBIT;
  signal \$38304\    : AGCBIT;
  signal  \38305\    : AGCBIT;
  signal \$38305\    : AGCBIT;
  signal  \38306\    : AGCBIT; signal  \FS18\     : AGCBIT;
  signal  \38307\    : AGCBIT; signal  \F18B\     : AGCBIT;
  signal  \38311\    : AGCBIT; signal  \CHAT14\   : AGCBIT;
  signal  \38312\    : AGCBIT; signal  \F19A\     : AGCBIT;
  signal  \38313\    : AGCBIT;
  signal \$38313\    : AGCBIT;
  signal  \38314\    : AGCBIT;
  signal \$38314\    : AGCBIT;
  signal  \38315\    : AGCBIT;
  signal \$38315\    : AGCBIT;
  signal  \38316\    : AGCBIT; signal  \FS19\     : AGCBIT;
  signal  \38317\    : AGCBIT; signal  \F19B\     : AGCBIT;
  signal  \38321\    : AGCBIT; signal  \CHBT01\   : AGCBIT;
  signal  \38322\    : AGCBIT; signal  \F20A\     : AGCBIT;
  signal  \38323\    : AGCBIT;
  signal \$38323\    : AGCBIT;
  signal  \38324\    : AGCBIT;
  signal \$38324\    : AGCBIT;
  signal  \38325\    : AGCBIT;
  signal \$38325\    : AGCBIT;
  signal  \38326\    : AGCBIT; signal  \FS20\     : AGCBIT;
  signal  \38327\    : AGCBIT; signal  \F20B\     : AGCBIT;
  signal  \38331\    : AGCBIT; signal  \CHBT02\   : AGCBIT;
  signal  \38332\    : AGCBIT; signal  \F21A\     : AGCBIT;
  signal  \38333\    : AGCBIT;
  signal \$38333\    : AGCBIT;
  signal  \38334\    : AGCBIT;
  signal \$38334\    : AGCBIT;
  signal  \38335\    : AGCBIT;
  signal \$38335\    : AGCBIT;
  signal  \38336\    : AGCBIT; signal  \FS21\     : AGCBIT;
  signal  \38337\    : AGCBIT; signal  \F21B\     : AGCBIT;
  signal  \38341\    : AGCBIT; signal  \CHBT03\   : AGCBIT;
  signal  \38342\    : AGCBIT; signal  \F22A\     : AGCBIT;
  signal  \38343\    : AGCBIT;
  signal \$38343\    : AGCBIT;
  signal  \38344\    : AGCBIT;
  signal \$38344\    : AGCBIT;
  signal  \38345\    : AGCBIT;
  signal \$38345\    : AGCBIT;
  signal  \38346\    : AGCBIT; signal  \FS22\     : AGCBIT;
  signal  \38347\    : AGCBIT; signal  \F22B\     : AGCBIT;
  signal  \38351\    : AGCBIT; signal  \CHBT04\   : AGCBIT;
  signal  \38352\    : AGCBIT; signal  \F23A\     : AGCBIT;
  signal  \38353\    : AGCBIT;
  signal \$38353\    : AGCBIT;
  signal  \38354\    : AGCBIT;
  signal \$38354\    : AGCBIT;
  signal  \38355\    : AGCBIT;
  signal \$38355\    : AGCBIT;
  signal  \38356\    : AGCBIT; signal  \FS23\     : AGCBIT;
  signal  \38357\    : AGCBIT; signal  \F23B\     : AGCBIT;
  signal  \38361\    : AGCBIT; signal  \CHBT05\   : AGCBIT;
  signal  \38362\    : AGCBIT; signal  \F24A\     : AGCBIT;
  signal  \38363\    : AGCBIT;
  signal \$38363\    : AGCBIT;
  signal  \38364\    : AGCBIT;
  signal \$38364\    : AGCBIT;
  signal  \38365\    : AGCBIT;
  signal \$38365\    : AGCBIT;
  signal  \38366\    : AGCBIT; signal  \FS24\     : AGCBIT;
  signal  \38367\    : AGCBIT; signal  \F24B\     : AGCBIT;
  signal  \38371\    : AGCBIT; signal  \CHBT06\   : AGCBIT;
  signal  \38372\    : AGCBIT; signal  \F25A\     : AGCBIT;
  signal  \38373\    : AGCBIT;
  signal \$38373\    : AGCBIT;
  signal  \38374\    : AGCBIT;
  signal \$38374\    : AGCBIT;
  signal  \38375\    : AGCBIT;
  signal \$38375\    : AGCBIT;
  signal  \38376\    : AGCBIT; signal  \FS25\     : AGCBIT;
  signal  \38377\    : AGCBIT; signal  \F25B\     : AGCBIT;
  signal  \38390\    : AGCBIT; signal  \F18AX\    : AGCBIT;
  signal  \38391\    : AGCBIT; signal  \F07A/\    : AGCBIT;
  signal  \38401\    : AGCBIT; signal  \CHBT07\   : AGCBIT;
  signal  \38402\    : AGCBIT; signal  \F26A\     : AGCBIT;
  signal  \38403\    : AGCBIT;
  signal \$38403\    : AGCBIT;
  signal  \38404\    : AGCBIT;
  signal \$38404\    : AGCBIT;
  signal  \38405\    : AGCBIT;
  signal \$38405\    : AGCBIT;
  signal  \38406\    : AGCBIT; signal  \FS26\     : AGCBIT;
  signal  \38407\    : AGCBIT; signal  \F26B\     : AGCBIT;
  signal  \38411\    : AGCBIT; signal  \CHBT08\   : AGCBIT;
  signal  \38412\    : AGCBIT; signal  \F27A\     : AGCBIT;
  signal  \38413\    : AGCBIT;
  signal \$38413\    : AGCBIT;
  signal  \38414\    : AGCBIT;
  signal \$38414\    : AGCBIT;
  signal  \38415\    : AGCBIT;
  signal \$38415\    : AGCBIT;
  signal  \38416\    : AGCBIT; signal  \FS27\     : AGCBIT;
  signal  \38417\    : AGCBIT; signal  \F27B\     : AGCBIT;
  signal  \38421\    : AGCBIT; signal  \CHBT09\   : AGCBIT;
  signal  \38422\    : AGCBIT; signal  \F28A\     : AGCBIT;
  signal  \38423\    : AGCBIT;
  signal \$38423\    : AGCBIT;
  signal  \38424\    : AGCBIT;
  signal \$38424\    : AGCBIT;
  signal  \38425\    : AGCBIT;
  signal \$38425\    : AGCBIT;
  signal  \38426\    : AGCBIT; signal  \FS28\     : AGCBIT;
  signal  \38427\    : AGCBIT; signal  \F28B\     : AGCBIT;
  signal  \38431\    : AGCBIT; signal  \CHBT10\   : AGCBIT;
  signal  \38432\    : AGCBIT; signal  \F29A\     : AGCBIT;
  signal  \38433\    : AGCBIT;
  signal \$38433\    : AGCBIT;
  signal  \38434\    : AGCBIT;
  signal \$38434\    : AGCBIT;
  signal  \38435\    : AGCBIT;
  signal \$38435\    : AGCBIT;
  signal  \38436\    : AGCBIT; signal  \FS29\     : AGCBIT;
  signal  \38437\    : AGCBIT; signal  \F29B\     : AGCBIT;
  signal  \38441\    : AGCBIT; signal  \CHBT11\   : AGCBIT;
  signal  \38442\    : AGCBIT; signal  \F30A\     : AGCBIT;
  signal  \38443\    : AGCBIT;
  signal \$38443\    : AGCBIT;
  signal  \38444\    : AGCBIT;
  signal \$38444\    : AGCBIT;
  signal  \38445\    : AGCBIT;
  signal \$38445\    : AGCBIT;
  signal  \38446\    : AGCBIT; signal  \FS30\     : AGCBIT;
  signal  \38447\    : AGCBIT; signal  \F30B\     : AGCBIT;
  signal  \38451\    : AGCBIT; signal  \CHBT12\   : AGCBIT;
  signal  \38452\    : AGCBIT; signal  \F31A\     : AGCBIT;
  signal  \38453\    : AGCBIT;
  signal \$38453\    : AGCBIT;
  signal  \38454\    : AGCBIT;
  signal \$38454\    : AGCBIT;
  signal  \38455\    : AGCBIT;
  signal \$38455\    : AGCBIT;
  signal  \38456\    : AGCBIT; signal  \FS31\     : AGCBIT;
  signal  \38457\    : AGCBIT; signal  \F31B\     : AGCBIT;
  signal  \38461\    : AGCBIT; signal  \CHBT13\   : AGCBIT;
  signal  \38462\    : AGCBIT; signal  \F32A\     : AGCBIT;
  signal  \38463\    : AGCBIT;
  signal \$38463\    : AGCBIT;
  signal  \38464\    : AGCBIT;
  signal \$38464\    : AGCBIT;
  signal  \38465\    : AGCBIT;
  signal \$38465\    : AGCBIT;
  signal  \38466\    : AGCBIT; signal  \FS32\     : AGCBIT;
  signal  \38467\    : AGCBIT; signal  \F32B\     : AGCBIT;
  signal  \38471\    : AGCBIT; signal  \CHBT14\   : AGCBIT;
  signal  \38472\    : AGCBIT; signal  \F33A\     : AGCBIT;
  signal  \38473\    : AGCBIT;
  signal \$38473\    : AGCBIT;
  signal  \38474\    : AGCBIT;
  signal \$38474\    : AGCBIT;
  signal  \38475\    : AGCBIT;
  signal \$38475\    : AGCBIT;
  signal  \38476\    : AGCBIT; signal  \FS33\     : AGCBIT;
  signal  \38477\    : AGCBIT; signal  \F33B\     : AGCBIT;
  signal  \38490\    : AGCBIT; signal  \F18A/\    : AGCBIT;
  signal  \38491\    : AGCBIT; signal  \F03B/\    : AGCBIT;
  signal  \37101\    : AGCBIT;
  signal  \37102\    : AGCBIT;
  signal \$37102\    : AGCBIT;
  signal  \37103\    : AGCBIT;
  signal \$37103\    : AGCBIT;
  signal  \37104\    : AGCBIT; signal  \PHS2\     : AGCBIT;
  signal  \37105\    : AGCBIT;
  signal \$37105\    : AGCBIT;
  signal  \37106\    : AGCBIT;
  signal  \37107\    : AGCBIT;
  signal  \37108\    : AGCBIT; signal  \PHS4\     : AGCBIT;
  signal  \37109\    : AGCBIT; signal  \PHS4/\    : AGCBIT;
  signal  \37111\    : AGCBIT;
  signal  \37112\    : AGCBIT;
  signal \$37112\    : AGCBIT;
  signal  \37113\    : AGCBIT;
  signal \$37113\    : AGCBIT;
  signal  \37114\    : AGCBIT;
  signal  \37115\    : AGCBIT; signal  \RINGA/\   : AGCBIT;
  signal  \37117\    : AGCBIT;
  signal \$37117\    : AGCBIT;
  signal  \37118\    : AGCBIT;
  signal  \37119\    : AGCBIT; signal  \RINGB/\   : AGCBIT;
  signal  \37121\    : AGCBIT;
  signal  \37122\    : AGCBIT; signal  \ODDSET/\  : AGCBIT;
  signal  \37125\    : AGCBIT; signal  \EVNSET\   : AGCBIT;
  signal  \37126\    : AGCBIT; signal  \EVNSET/\  : AGCBIT;
  signal  \37129\    : AGCBIT; signal  \RT\       : AGCBIT;
  signal  \37130\    : AGCBIT; signal  \WT\       : AGCBIT;
  signal  \37131\    : AGCBIT; signal  \WT/\      : AGCBIT;
  signal  \37135\    : AGCBIT; signal  \TT/\      : AGCBIT;
  signal \&37136\    : AGCBIT;
  signal  \37137\    : AGCBIT; signal  \CLK\      : AGCBIT;
  signal \&37138\    : AGCBIT;
  signal  \37139\    : AGCBIT;
  signal  \37140\    : AGCBIT; signal  \CT\       : AGCBIT;
  signal  \37142\    : AGCBIT; signal  \CT/\      : AGCBIT;
  signal  \37148\    : AGCBIT;
  signal  \37149\    : AGCBIT;
  signal \$37149\    : AGCBIT;
  signal  \37150\    : AGCBIT;
  signal  \37151\    : AGCBIT; signal  \OVFSTB/\  : AGCBIT;
  signal  \37152\    : AGCBIT;
  signal \$37152\    : AGCBIT;
  signal  \37153\    : AGCBIT;
  signal \$37153\    : AGCBIT;
  signal  \37154\    : AGCBIT;
  signal \$37154\    : AGCBIT;
  signal  \37155\    : AGCBIT; signal  \PHS2/\    : AGCBIT;
  signal  \37201\    : AGCBIT;
  signal  \37202\    : AGCBIT;
  signal  \37203\    : AGCBIT; signal  \P01\      : AGCBIT;
  signal \$37203\    : AGCBIT;
  signal  \37204\    : AGCBIT; signal  \P01/\     : AGCBIT;
  signal  \37205\    : AGCBIT;
  signal  \37206\    : AGCBIT;
  signal  \37207\    : AGCBIT; signal  \P02\      : AGCBIT;
  signal \$37207\    : AGCBIT;
  signal  \37208\    : AGCBIT; signal  \P02/\     : AGCBIT;
  signal  \37209\    : AGCBIT;
  signal  \37210\    : AGCBIT;
  signal  \37211\    : AGCBIT; signal  \P03\      : AGCBIT;
  signal \$37211\    : AGCBIT;
  signal  \37212\    : AGCBIT; signal  \P03/\     : AGCBIT;
  signal  \37213\    : AGCBIT;
  signal  \37214\    : AGCBIT;
  signal  \37215\    : AGCBIT; signal  \P04\      : AGCBIT;
  signal \$37215\    : AGCBIT;
  signal  \37216\    : AGCBIT; signal  \P04/\     : AGCBIT;
  signal  \37217\    : AGCBIT;
  signal  \37218\    : AGCBIT;
  signal  \37219\    : AGCBIT; signal  \P05\      : AGCBIT;
  signal \$37219\    : AGCBIT;
  signal  \37220\    : AGCBIT; signal  \P05/\     : AGCBIT;
  signal  \37221\    : AGCBIT; signal  \F01D\     : AGCBIT;
  signal  \37222\    : AGCBIT; signal  \F01B\     : AGCBIT;
  signal \$37222\    : AGCBIT;
  signal  \37223\    : AGCBIT; signal  \F01A\     : AGCBIT;
  signal \$37223\    : AGCBIT;
  signal  \37224\    : AGCBIT; signal  \F01C\     : AGCBIT;
  signal  \37225\    : AGCBIT; signal  \FS01/\    : AGCBIT;
  signal \$37225\    : AGCBIT;
  signal  \37226\    : AGCBIT; signal  \FS01\     : AGCBIT;
  signal \&37227\    : AGCBIT;
  signal  \37228\    : AGCBIT; signal  \GOSET/\   : AGCBIT;
  signal \$37228\    : AGCBIT;
  signal  \37229\    : AGCBIT;
  signal  \37230\    : AGCBIT;
  signal  \37231\    : AGCBIT;
  signal  \37232\    : AGCBIT;
  signal  \37233\    : AGCBIT;
  signal \$37233\    : AGCBIT;
  signal  \37234\    : AGCBIT; signal  \STOPA\    : AGCBIT;
  signal  \37235\    : AGCBIT;
  signal  \37236\    : AGCBIT;
  signal  \37237\    : AGCBIT;
  signal  \37238\    : AGCBIT;
  signal \$37238\    : AGCBIT;
  signal  \37239\    : AGCBIT;
  signal  \37240\    : AGCBIT; signal  \GOJAM/\   : AGCBIT;
  signal \&37241\    : AGCBIT;
  signal  \37242\    : AGCBIT; signal  \STOP/\    : AGCBIT;
  signal  \37243\    : AGCBIT; signal  \STOP\     : AGCBIT;
  signal \&37244\    : AGCBIT;
  signal  \37245\    : AGCBIT; signal  \GOJAM\    : AGCBIT;
  signal \&37251\    : AGCBIT;
  signal  \37255\    : AGCBIT; signal  \SB0\      : AGCBIT;
  signal  \37256\    : AGCBIT; signal  \SB1\      : AGCBIT;
  signal  \37257\    : AGCBIT; signal  \SB2\      : AGCBIT;
  signal  \37258\    : AGCBIT; signal  \SB4\      : AGCBIT;
  signal  \37259\    : AGCBIT; signal  \EDSET\    : AGCBIT;
  signal  \37301\    : AGCBIT; signal  \T12\      : AGCBIT;
  signal  \37302\    : AGCBIT; signal  \T12DC/\   : AGCBIT;
  signal  \37303\    : AGCBIT;
  signal \$37303\    : AGCBIT;
  signal  \37304\    : AGCBIT;
  signal  \37305\    : AGCBIT; signal  \T01DC/\   : AGCBIT;
  signal \$37305\    : AGCBIT;
  signal  \37306\    : AGCBIT;
  signal  \37307\    : AGCBIT; signal  \T01\      : AGCBIT;
  signal  \37308\    : AGCBIT;
  signal  \37309\    : AGCBIT; signal  \T02DC/\   : AGCBIT;
  signal \$37309\    : AGCBIT;
  signal  \37310\    : AGCBIT;
  signal  \37311\    : AGCBIT; signal  \T02\      : AGCBIT;
  signal  \37312\    : AGCBIT;
  signal  \37313\    : AGCBIT; signal  \T03DC/\   : AGCBIT;
  signal \$37313\    : AGCBIT;
  signal  \37314\    : AGCBIT;
  signal  \37315\    : AGCBIT; signal  \T03\      : AGCBIT;
  signal  \37316\    : AGCBIT;
  signal  \37317\    : AGCBIT;
  signal \$37317\    : AGCBIT;
  signal  \37318\    : AGCBIT;
  signal  \37319\    : AGCBIT; signal  \T04\      : AGCBIT;
  signal  \37320\    : AGCBIT;
  signal  \37321\    : AGCBIT;
  signal \$37321\    : AGCBIT;
  signal  \37322\    : AGCBIT;
  signal  \37323\    : AGCBIT; signal  \T05\      : AGCBIT;
  signal  \37325\    : AGCBIT;
  signal  \37326\    : AGCBIT; signal  \T06DC/\   : AGCBIT;
  signal \$37326\    : AGCBIT;
  signal  \37327\    : AGCBIT;
  signal  \37328\    : AGCBIT; signal  \T06\      : AGCBIT;
  signal  \37329\    : AGCBIT;
  signal  \37330\    : AGCBIT; signal  \T07DC/\   : AGCBIT;
  signal \$37330\    : AGCBIT;
  signal  \37331\    : AGCBIT;
  signal  \37332\    : AGCBIT; signal  \T07\      : AGCBIT;
  signal  \37333\    : AGCBIT;
  signal  \37334\    : AGCBIT; signal  \T08DC/\   : AGCBIT;
  signal \$37334\    : AGCBIT;
  signal  \37335\    : AGCBIT;
  signal  \37336\    : AGCBIT; signal  \T08\      : AGCBIT;
  signal  \37337\    : AGCBIT;
  signal  \37338\    : AGCBIT; signal  \T09DC/\   : AGCBIT;
  signal \$37338\    : AGCBIT;
  signal  \37339\    : AGCBIT;
  signal  \37340\    : AGCBIT; signal  \T09\      : AGCBIT;
  signal  \37341\    : AGCBIT;
  signal  \37342\    : AGCBIT; signal  \T10DC/\   : AGCBIT;
  signal \$37342\    : AGCBIT;
  signal  \37343\    : AGCBIT;
  signal  \37344\    : AGCBIT; signal  \T10\      : AGCBIT;
  signal  \37345\    : AGCBIT;
  signal \$37345\    : AGCBIT;
  signal  \37346\    : AGCBIT;
  signal \$37346\    : AGCBIT;
  signal  \37347\    : AGCBIT;
  signal \$37347\    : AGCBIT;
  signal  \37348\    : AGCBIT;
  signal  \37349\    : AGCBIT; signal  \T11\      : AGCBIT;
  signal  \37350\    : AGCBIT; signal  \RT/\      : AGCBIT;
  signal  \37353\    : AGCBIT; signal  \OVF\      : AGCBIT;
  signal  \37354\    : AGCBIT; signal  \UNF\      : AGCBIT;
  signal  \37355\    : AGCBIT; signal  \T12SET\   : AGCBIT;
  signal \&37356\    : AGCBIT;
  signal \&37357\    : AGCBIT;
  signal \&37358\    : AGCBIT;
  signal \&37360\    : AGCBIT;
  signal  \37401\    : AGCBIT; signal  \T01/\     : AGCBIT;
  signal \&37404\    : AGCBIT;
  signal  \37405\    : AGCBIT; signal  \T02/\     : AGCBIT;
  signal \&37407\    : AGCBIT;
  signal  \37408\    : AGCBIT; signal  \T03/\     : AGCBIT;
  signal \&37411\    : AGCBIT;
  signal  \37412\    : AGCBIT; signal  \T04/\     : AGCBIT;
  signal \&37415\    : AGCBIT;
  signal  \37416\    : AGCBIT; signal  \T05/\     : AGCBIT;
  signal \&37422\    : AGCBIT;
  signal  \37423\    : AGCBIT; signal  \T06/\     : AGCBIT;
  signal \&37427\    : AGCBIT;
  signal  \37428\    : AGCBIT; signal  \T07/\     : AGCBIT;
  signal \&37432\    : AGCBIT;
  signal  \37433\    : AGCBIT; signal  \T08/\     : AGCBIT;
  signal \&37437\    : AGCBIT;
  signal  \37438\    : AGCBIT; signal  \T09/\     : AGCBIT;
  signal \&37442\    : AGCBIT;
  signal  \37443\    : AGCBIT; signal  \T10/\     : AGCBIT;
  signal \&37447\    : AGCBIT;
  signal  \37448\    : AGCBIT; signal  \T11/\     : AGCBIT;
  signal \&37450\    : AGCBIT;
  signal  \37451\    : AGCBIT; signal  \T12/\     : AGCBIT;
  signal \&37454\    : AGCBIT;
  signal  \37455\    : AGCBIT; signal  \OVF/\     : AGCBIT;
  signal  \37456\    : AGCBIT; signal  \UNF/\     : AGCBIT;
  signal  \30001\    : AGCBIT;
  signal \$30001\    : AGCBIT;
  signal  \30002\    : AGCBIT;
  signal  \30003\    : AGCBIT;
  signal  \30004\    : AGCBIT; signal  \NISQL/\   : AGCBIT;
  signal  \30005\    : AGCBIT;
  signal  \30006\    : AGCBIT;
  signal  \30007\    : AGCBIT; signal  \CSQG\     : AGCBIT;
  signal  \30009\    : AGCBIT; signal  \RBSQ\     : AGCBIT;
  signal  \30010\    : AGCBIT;
  signal  \30011\    : AGCBIT; signal  \WSQG/\    : AGCBIT;
  signal  \30013\    : AGCBIT;
  signal  \30014\    : AGCBIT;
  signal  \30015\    : AGCBIT;
  signal  \30016\    : AGCBIT;
  signal \$30016\    : AGCBIT;
  signal  \30017\    : AGCBIT; signal  \SQR16\    : AGCBIT;
  signal  \30018\    : AGCBIT;
  signal \$30018\    : AGCBIT;
  signal  \30019\    : AGCBIT; signal  \SQR14\    : AGCBIT;
  signal  \30020\    : AGCBIT;
  signal \$30020\    : AGCBIT;
  signal  \30021\    : AGCBIT; signal  \SQR13\    : AGCBIT;
  signal \&30022\    : AGCBIT;
  signal  \30023\    : AGCBIT;
  signal  \30024\    : AGCBIT;
  signal \&30025\    : AGCBIT;
  signal \&30028\    : AGCBIT;
  signal  \30031\    : AGCBIT;
  signal  \30032\    : AGCBIT;
  signal  \30034\    : AGCBIT;
  signal  \30036\    : AGCBIT;
  signal  \30037\    : AGCBIT;
  signal  \30038\    : AGCBIT;
  signal  \30039\    : AGCBIT; signal  \SQ5\      : AGCBIT;
  signal  \30040\    : AGCBIT;
  signal  \30041\    : AGCBIT;
  signal  \30042\    : AGCBIT;
  signal  \30043\    : AGCBIT;
  signal  \30044\    : AGCBIT;
  signal  \30045\    : AGCBIT; signal  \SQ0/\     : AGCBIT;
  signal  \30048\    : AGCBIT; signal  \SQ1/\     : AGCBIT;
  signal  \30049\    : AGCBIT; signal  \SQ2/\     : AGCBIT;
  signal  \30053\    : AGCBIT; signal  \SQ3/\     : AGCBIT;
  signal  \30054\    : AGCBIT; signal  \SQ4/\     : AGCBIT;
  signal  \30055\    : AGCBIT; signal  \SQ6/\     : AGCBIT;
  signal  \30056\    : AGCBIT; signal  \SQ7/\     : AGCBIT;
  signal  \30057\    : AGCBIT; signal  \CON1\     : AGCBIT;
  signal  \30058\    : AGCBIT; signal  \CON2\     : AGCBIT;
  signal \&30059\    : AGCBIT;
  signal  \30061\    : AGCBIT; signal  \INKBT1\   : AGCBIT;
  signal  \30101\    : AGCBIT;
  signal  \30103\    : AGCBIT;
  signal \$30103\    : AGCBIT;
  signal  \30104\    : AGCBIT; signal  \INHINT\   : AGCBIT;
  signal  \30105\    : AGCBIT; signal  \IIP/\     : AGCBIT;
  signal \$30105\    : AGCBIT;
  signal  \30106\    : AGCBIT; signal  \IIP\      : AGCBIT;
  signal  \30107\    : AGCBIT; signal  \STRTFC\   : AGCBIT;
  signal  \30108\    : AGCBIT;
  signal  \30109\    : AGCBIT;
  signal \$30109\    : AGCBIT;
  signal  \30110\    : AGCBIT; signal  \FUTEXT\   : AGCBIT;
  signal \&30111\    : AGCBIT;
  signal \&30112\    : AGCBIT;
  signal  \30113\    : AGCBIT;
  signal  \30114\    : AGCBIT;
  signal  \30115\    : AGCBIT;
  signal \&30116\    : AGCBIT;
  signal  \30117\    : AGCBIT; signal  \RPTSET\   : AGCBIT;
  signal \&30118\    : AGCBIT;
  signal  \30119\    : AGCBIT;
  signal \$30119\    : AGCBIT;
  signal  \30120\    : AGCBIT;
  signal  \30121\    : AGCBIT;
  signal \$30121\    : AGCBIT;
  signal  \30122\    : AGCBIT;
  signal \&30123\    : AGCBIT;
  signal  \30124\    : AGCBIT; signal  \SQEXT/\   : AGCBIT;
  signal  \30127\    : AGCBIT; signal  \RPTFRC\   : AGCBIT;
  signal  \30129\    : AGCBIT;
  signal  \30130\    : AGCBIT;
  signal  \30131\    : AGCBIT;
  signal  \30132\    : AGCBIT;
  signal \$30132\    : AGCBIT;
  signal  \30133\    : AGCBIT; signal  \SQR12\    : AGCBIT;
  signal  \30134\    : AGCBIT;
  signal \$30134\    : AGCBIT;
  signal  \30135\    : AGCBIT; signal  \SQR11\    : AGCBIT;
  signal  \30136\    : AGCBIT;
  signal \$30136\    : AGCBIT;
  signal  \30137\    : AGCBIT;
  signal \&30138\    : AGCBIT;
  signal \&30139\    : AGCBIT;
  signal \&30140\    : AGCBIT;
  signal  \30141\    : AGCBIT; signal  \QC0\      : AGCBIT;
  signal  \30142\    : AGCBIT;
  signal  \30143\    : AGCBIT;
  signal  \30144\    : AGCBIT;
  signal  \30145\    : AGCBIT; signal  \QC0/\     : AGCBIT;
  signal  \30148\    : AGCBIT; signal  \QC1/\     : AGCBIT;
  signal  \30151\    : AGCBIT; signal  \QC2/\     : AGCBIT;
  signal  \30152\    : AGCBIT; signal  \QC3/\     : AGCBIT;
  signal  \30154\    : AGCBIT; signal  \SQR10\    : AGCBIT;
  signal  \30156\    : AGCBIT; signal  \SQR10/\   : AGCBIT;
  signal  \30157\    : AGCBIT; signal  \SQR12/\   : AGCBIT;
  signal  \30160\    : AGCBIT; signal  \SQEXT\    : AGCBIT;
  signal  \30301\    : AGCBIT;
  signal  \30302\    : AGCBIT;
  signal  \30303\    : AGCBIT; signal  \SQ5QC0/\  : AGCBIT;
  signal  \30304\    : AGCBIT;
  signal  \30305\    : AGCBIT; signal  \IC1\      : AGCBIT;
  signal  \30306\    : AGCBIT; signal  \IC2\      : AGCBIT;
  signal  \30309\    : AGCBIT; signal  \IC2/\     : AGCBIT;
  signal  \30310\    : AGCBIT; signal  \SQ5/\     : AGCBIT;
  signal  \30313\    : AGCBIT; signal  \IC11\     : AGCBIT;
  signal  \30314\    : AGCBIT;
  signal  \30315\    : AGCBIT;
  signal  \30316\    : AGCBIT; signal  \EXST1/\   : AGCBIT;
  signal  \30317\    : AGCBIT; signal  \IC6\      : AGCBIT;
  signal  \30318\    : AGCBIT; signal  \IC7\      : AGCBIT;
  signal  \30319\    : AGCBIT; signal  \TC0\      : AGCBIT;
  signal  \30320\    : AGCBIT; signal  \TCF0\     : AGCBIT;
  signal  \30321\    : AGCBIT; signal  \NEXST0\   : AGCBIT;
  signal  \30322\    : AGCBIT; signal  \TC0/\     : AGCBIT;
  signal  \30323\    : AGCBIT; signal  \IC3/\     : AGCBIT;
  signal  \30324\    : AGCBIT; signal  \NEXST0/\  : AGCBIT;
  signal  \30326\    : AGCBIT; signal  \IC3\      : AGCBIT;
  signal  \30327\    : AGCBIT; signal  \DCS0\     : AGCBIT;
  signal  \30328\    : AGCBIT; signal  \DCA0\     : AGCBIT;
  signal  \30329\    : AGCBIT; signal  \IC4/\     : AGCBIT;
  signal  \30330\    : AGCBIT; signal  \IC4\      : AGCBIT;
  signal  \30331\    : AGCBIT; signal  \IC13/\    : AGCBIT;
  signal \&30332\    : AGCBIT;
  signal  \30333\    : AGCBIT; signal  \IC13\     : AGCBIT;
  signal  \30335\    : AGCBIT;
  signal  \30336\    : AGCBIT;
  signal  \30337\    : AGCBIT;
  signal  \30338\    : AGCBIT; signal  \IC5\      : AGCBIT;
  signal  \30339\    : AGCBIT; signal  \IC5/\     : AGCBIT;
  signal  \30340\    : AGCBIT; signal  \IC9/\     : AGCBIT;
  signal  \30341\    : AGCBIT; signal  \LXCH0\    : AGCBIT;
  signal  \30342\    : AGCBIT; signal  \QXCH0\    : AGCBIT;
  signal  \30343\    : AGCBIT; signal  \QXCH0/\   : AGCBIT;
  signal \&30344\    : AGCBIT;
  signal  \30345\    : AGCBIT; signal  \IC9\      : AGCBIT;
  signal  \30346\    : AGCBIT; signal  \IC8/\     : AGCBIT;
  signal  \30347\    : AGCBIT;
  signal  \30348\    : AGCBIT; signal  \TS0\      : AGCBIT;
  signal  \30349\    : AGCBIT; signal  \EXST0/\   : AGCBIT;
  signal  \30350\    : AGCBIT; signal  \TS0/\     : AGCBIT;
  signal  \30352\    : AGCBIT; signal  \DXCH0\    : AGCBIT;
  signal  \30354\    : AGCBIT; signal  \DAS0\     : AGCBIT;
  signal  \30356\    : AGCBIT; signal  \IC10/\    : AGCBIT;
  signal  \30357\    : AGCBIT; signal  \IC10\     : AGCBIT;
  signal  \30360\    : AGCBIT;
  signal  \30401\    : AGCBIT; signal  \DAS0/\    : AGCBIT;
  signal  \30403\    : AGCBIT; signal  \BZF0\     : AGCBIT;
  signal  \30404\    : AGCBIT; signal  \BZF0/\    : AGCBIT;
  signal  \30405\    : AGCBIT; signal  \BMF0\     : AGCBIT;
  signal  \30406\    : AGCBIT; signal  \BMF0/\    : AGCBIT;
  signal  \30407\    : AGCBIT;
  signal  \30408\    : AGCBIT;
  signal  \30409\    : AGCBIT; signal  \IC16/\    : AGCBIT;
  signal  \30410\    : AGCBIT; signal  \IC15/\    : AGCBIT;
  signal  \30411\    : AGCBIT; signal  \IC16\     : AGCBIT;
  signal  \30412\    : AGCBIT; signal  \IC17\     : AGCBIT;
  signal  \30413\    : AGCBIT; signal  \IC15\     : AGCBIT;
  signal  \30415\    : AGCBIT; signal  \CCS0\     : AGCBIT;
  signal  \30416\    : AGCBIT; signal  \CCS0/\    : AGCBIT;
  signal  \30417\    : AGCBIT;
  signal \&30418\    : AGCBIT;
  signal  \30419\    : AGCBIT; signal  \DAS1/\    : AGCBIT;
  signal  \30421\    : AGCBIT; signal  \DAS1\     : AGCBIT;
  signal  \30422\    : AGCBIT; signal  \IC12/\    : AGCBIT;
  signal  \30423\    : AGCBIT; signal  \IC12\     : AGCBIT;
  signal  \30424\    : AGCBIT; signal  \ADS0\     : AGCBIT;
  signal  \30425\    : AGCBIT; signal  \INCR0\    : AGCBIT;
  signal  \30426\    : AGCBIT; signal  \MSU0\     : AGCBIT;
  signal  \30427\    : AGCBIT; signal  \MSU0/\    : AGCBIT;
  signal  \30428\    : AGCBIT; signal  \AUG0\     : AGCBIT;
  signal  \30429\    : AGCBIT; signal  \AUG0/\    : AGCBIT;
  signal  \30430\    : AGCBIT; signal  \DIM0\     : AGCBIT;
  signal  \30431\    : AGCBIT; signal  \DIM0/\    : AGCBIT;
  signal  \30432\    : AGCBIT; signal  \MP3\      : AGCBIT;
  signal  \30433\    : AGCBIT; signal  \MP3/\     : AGCBIT;
  signal  \30435\    : AGCBIT; signal  \MP1\      : AGCBIT;
  signal  \30436\    : AGCBIT; signal  \MP1/\     : AGCBIT;
  signal  \30437\    : AGCBIT; signal  \MP0\      : AGCBIT;
  signal \&30438\    : AGCBIT;
  signal  \30439\    : AGCBIT; signal  \MP0/\     : AGCBIT;
  signal  \30441\    : AGCBIT; signal  \TCSAJ3\   : AGCBIT;
  signal  \30442\    : AGCBIT; signal  \TCSAJ3/\  : AGCBIT;
  signal  \30443\    : AGCBIT; signal  \RSM3\     : AGCBIT;
  signal  \30444\    : AGCBIT; signal  \RSM3/\    : AGCBIT;
  signal  \30445\    : AGCBIT; signal  \SU0\      : AGCBIT;
  signal  \30446\    : AGCBIT; signal  \MASK0\    : AGCBIT;
  signal  \30447\    : AGCBIT; signal  \MASK0/\   : AGCBIT;
  signal  \30448\    : AGCBIT; signal  \AD0\      : AGCBIT;
  signal  \30449\    : AGCBIT; signal  \NDX0\     : AGCBIT;
  signal  \30450\    : AGCBIT; signal  \NDX0/\    : AGCBIT;
  signal  \30451\    : AGCBIT; signal  \NDXX1\    : AGCBIT;
  signal  \30452\    : AGCBIT; signal  \NDXX1/\   : AGCBIT;
  signal  \30453\    : AGCBIT; signal  \GOJ1\     : AGCBIT;
  signal  \30454\    : AGCBIT; signal  \GOJ1/\    : AGCBIT;
  signal  \30455\    : AGCBIT;
  signal  \30456\    : AGCBIT; signal  \IC14\     : AGCBIT;
  signal  \36101\    : AGCBIT; signal  \DIVSTG\   : AGCBIT;
  signal  \36102\    : AGCBIT; signal  \T12USE/\  : AGCBIT;
  signal \$36102\    : AGCBIT;
  signal  \36103\    : AGCBIT;
  signal  \36104\    : AGCBIT;
  signal  \36105\    : AGCBIT;
  signal  \36106\    : AGCBIT; signal  \ST0/\     : AGCBIT;
  signal  \36108\    : AGCBIT; signal  \MP3A\     : AGCBIT;
  signal  \36109\    : AGCBIT;
  signal \$36109\    : AGCBIT;
  signal  \36110\    : AGCBIT;
  signal \&36112\    : AGCBIT;
  signal  \36113\    : AGCBIT;
  signal \$36113\    : AGCBIT;
  signal  \36114\    : AGCBIT;
  signal  \36115\    : AGCBIT;
  signal \$36115\    : AGCBIT;
  signal \&36116\    : AGCBIT;
  signal  \36117\    : AGCBIT; signal  \ST1/\     : AGCBIT;
  signal  \36118\    : AGCBIT;
  signal \$36118\    : AGCBIT;
  signal  \36119\    : AGCBIT;
  signal  \36120\    : AGCBIT; signal  \STG1\     : AGCBIT;
  signal \$36120\    : AGCBIT;
  signal  \36121\    : AGCBIT; signal  \ST1D\     : AGCBIT;
  signal  \36124\    : AGCBIT;
  signal \&36125\    : AGCBIT;
  signal  \36126\    : AGCBIT; signal  \ST1376/\  : AGCBIT;
  signal  \36127\    : AGCBIT; signal  \DV1376\   : AGCBIT;
  signal  \36128\    : AGCBIT; signal  \DV1376/\  : AGCBIT;
  signal \&36129\    : AGCBIT;
  signal  \36130\    : AGCBIT;
  signal \$36130\    : AGCBIT;
  signal  \36131\    : AGCBIT;
  signal  \36132\    : AGCBIT;
  signal \$36132\    : AGCBIT;
  signal \&36134\    : AGCBIT;
  signal  \36135\    : AGCBIT;
  signal \$36135\    : AGCBIT;
  signal  \36136\    : AGCBIT;
  signal  \36137\    : AGCBIT; signal  \STG2\     : AGCBIT;
  signal \$36137\    : AGCBIT;
  signal  \36138\    : AGCBIT; signal  \STD2\     : AGCBIT;
  signal  \36139\    : AGCBIT;
  signal  \36140\    : AGCBIT;
  signal  \36141\    : AGCBIT; signal  \ST3/\     : AGCBIT;
  signal  \36142\    : AGCBIT;
  signal \&36143\    : AGCBIT;
  signal  \36144\    : AGCBIT;
  signal  \36145\    : AGCBIT; signal  \ST4/\     : AGCBIT;
  signal  \36146\    : AGCBIT;
  signal \$36146\    : AGCBIT;
  signal  \36147\    : AGCBIT;
  signal  \36148\    : AGCBIT;
  signal \$36148\    : AGCBIT;
  signal  \36149\    : AGCBIT;
  signal \$36149\    : AGCBIT;
  signal  \36150\    : AGCBIT;
  signal  \36151\    : AGCBIT; signal  \STG3\     : AGCBIT;
  signal  \36152\    : AGCBIT;
  signal  \36153\    : AGCBIT; signal  \ST376\    : AGCBIT;
  signal  \36154\    : AGCBIT; signal  \ST376/\   : AGCBIT;
  signal  \36155\    : AGCBIT;
  signal  \36156\    : AGCBIT;
  signal  \36157\    : AGCBIT; signal  \DV3764\   : AGCBIT;
  signal \&36158\    : AGCBIT;
  signal \&36159\    : AGCBIT;
  signal \&36161\    : AGCBIT;
  signal  \36201\    : AGCBIT;
  signal  \36202\    : AGCBIT; signal  \DIV/\     : AGCBIT;
  signal  \36204\    : AGCBIT; signal  \DV0\      : AGCBIT;
  signal  \36205\    : AGCBIT; signal  \DV0/\     : AGCBIT;
  signal  \36206\    : AGCBIT; signal  \DV376\    : AGCBIT;
  signal  \36207\    : AGCBIT; signal  \DV376/\   : AGCBIT;
  signal  \36208\    : AGCBIT; signal  \DV4\      : AGCBIT;
  signal  \36209\    : AGCBIT; signal  \DV1\      : AGCBIT;
  signal  \36210\    : AGCBIT; signal  \DV1/\     : AGCBIT;
  signal  \36213\    : AGCBIT;
  signal  \36214\    : AGCBIT; signal  \SGUM\     : AGCBIT;
  signal \&36215\    : AGCBIT;
  signal  \36216\    : AGCBIT;
  signal  \36217\    : AGCBIT;
  signal  \36218\    : AGCBIT;
  signal \&36219\    : AGCBIT;
  signal  \36220\    : AGCBIT; signal  \BR1\      : AGCBIT;
  signal  \36221\    : AGCBIT;
  signal  \36222\    : AGCBIT;
  signal \$36222\    : AGCBIT;
  signal  \36224\    : AGCBIT;
  signal \&36225\    : AGCBIT;
  signal  \36226\    : AGCBIT; signal  \BR1/\     : AGCBIT;
  signal  \36227\    : AGCBIT;
  signal  \36228\    : AGCBIT;
  signal \$36228\    : AGCBIT;
  signal  \36230\    : AGCBIT;
  signal  \36231\    : AGCBIT;
  signal \&36232\    : AGCBIT;
  signal  \36233\    : AGCBIT;
  signal  \36236\    : AGCBIT;
  signal \&36237\    : AGCBIT;
  signal  \36238\    : AGCBIT; signal  \BR2\      : AGCBIT;
  signal  \36239\    : AGCBIT;
  signal  \36240\    : AGCBIT;
  signal  \36241\    : AGCBIT;
  signal \$36241\    : AGCBIT;
  signal  \36243\    : AGCBIT;
  signal  \36244\    : AGCBIT;
  signal \&36245\    : AGCBIT;
  signal  \36246\    : AGCBIT; signal  \BR2/\     : AGCBIT;
  signal \&36247\    : AGCBIT;
  signal  \36249\    : AGCBIT;
  signal \$36249\    : AGCBIT;
  signal \&36251\    : AGCBIT;
  signal  \36252\    : AGCBIT;
  signal \&36253\    : AGCBIT;
  signal \&36254\    : AGCBIT;
  signal \&36255\    : AGCBIT;
  signal \&36260\    : AGCBIT;
  signal \&36262\    : AGCBIT;
  signal  \36263\    : AGCBIT; signal  \TRSM/\    : AGCBIT;
  signal  \36264\    : AGCBIT; signal  \DVST/\    : AGCBIT;
  signal  \36301\    : AGCBIT; signal  \DV4/\     : AGCBIT;
  signal  \36303\    : AGCBIT;
  signal  \36304\    : AGCBIT;
  signal  \36305\    : AGCBIT; signal  \READ0\    : AGCBIT;
  signal  \36306\    : AGCBIT; signal  \READ0/\   : AGCBIT;
  signal  \36308\    : AGCBIT; signal  \WRITE0\   : AGCBIT;
  signal  \36309\    : AGCBIT; signal  \WRITE0/\  : AGCBIT;
  signal  \36310\    : AGCBIT; signal  \RAND0\    : AGCBIT;
  signal  \36312\    : AGCBIT; signal  \WAND0\    : AGCBIT;
  signal  \36313\    : AGCBIT; signal  \INOUT/\   : AGCBIT;
  signal  \36314\    : AGCBIT; signal  \INOUT\    : AGCBIT;
  signal  \36315\    : AGCBIT; signal  \ROR0\     : AGCBIT;
  signal  \36316\    : AGCBIT; signal  \WOR0\     : AGCBIT;
  signal  \36317\    : AGCBIT; signal  \WOR0/\    : AGCBIT;
  signal  \36318\    : AGCBIT; signal  \RXOR0\    : AGCBIT;
  signal  \36319\    : AGCBIT; signal  \RXOR0/\   : AGCBIT;
  signal  \36320\    : AGCBIT; signal  \RUPT0\    : AGCBIT;
  signal  \36321\    : AGCBIT; signal  \RUPT0/\   : AGCBIT;
  signal  \36322\    : AGCBIT; signal  \8PP4\     : AGCBIT;
  signal  \36323\    : AGCBIT; signal  \RUPT1\    : AGCBIT;
  signal  \36324\    : AGCBIT; signal  \RUPT1/\   : AGCBIT;
  signal \&36325\    : AGCBIT;
  signal  \36326\    : AGCBIT;
  signal  \36327\    : AGCBIT; signal  \PRINC\    : AGCBIT;
  signal  \36328\    : AGCBIT;
  signal  \36329\    : AGCBIT;
  signal  \36331\    : AGCBIT; signal  \RRPA\     : AGCBIT;
  signal  \36332\    : AGCBIT; signal  \3XP7\     : AGCBIT;
  signal  \36333\    : AGCBIT;
  signal  \36334\    : AGCBIT;
  signal \&36335\    : AGCBIT;
  signal  \36336\    : AGCBIT; signal  \9XP1\     : AGCBIT;
  signal  \36337\    : AGCBIT;
  signal  \36338\    : AGCBIT;
  signal \&36339\    : AGCBIT;
  signal  \36340\    : AGCBIT;
  signal  \36341\    : AGCBIT; signal  \5XP28\    : AGCBIT;
  signal  \36342\    : AGCBIT;
  signal  \36343\    : AGCBIT;
  signal  \36344\    : AGCBIT; signal  \5XP11\    : AGCBIT;
  signal \&36345\    : AGCBIT;
  signal \&36346\    : AGCBIT;
  signal \&36347\    : AGCBIT;
  signal  \36348\    : AGCBIT;
  signal  \36349\    : AGCBIT;
  signal  \36350\    : AGCBIT; signal  \WCH/\     : AGCBIT;
  signal  \36351\    : AGCBIT;
  signal  \36352\    : AGCBIT; signal  \2XP3\     : AGCBIT;
  signal  \36353\    : AGCBIT;
  signal  \36354\    : AGCBIT;
  signal \&36355\    : AGCBIT;
  signal  \36360\    : AGCBIT;
  signal  \36401\    : AGCBIT;
  signal  \36402\    : AGCBIT; signal  \R15\      : AGCBIT;
  signal  \36403\    : AGCBIT; signal  \RB2\      : AGCBIT;
  signal  \36404\    : AGCBIT; signal  \1XP10\    : AGCBIT;
  signal  \36405\    : AGCBIT; signal  \2PP1\     : AGCBIT;
  signal  \36406\    : AGCBIT;
  signal  \36407\    : AGCBIT;
  signal  \36408\    : AGCBIT; signal  \2XP5\     : AGCBIT;
  signal \&36409\    : AGCBIT;
  signal  \36410\    : AGCBIT; signal  \RSC/\     : AGCBIT;
  signal \&36411\    : AGCBIT;
  signal \&36412\    : AGCBIT;
  signal  \36413\    : AGCBIT;
  signal  \36414\    : AGCBIT;
  signal \&36415\    : AGCBIT;
  signal  \36416\    : AGCBIT; signal  \3XP2\     : AGCBIT;
  signal  \36417\    : AGCBIT; signal  \BR1B2\    : AGCBIT;
  signal  \36418\    : AGCBIT; signal  \BR1B2/\   : AGCBIT;
  signal  \36419\    : AGCBIT; signal  \BR12B\    : AGCBIT;
  signal  \36420\    : AGCBIT; signal  \BR12B/\   : AGCBIT;
  signal  \36421\    : AGCBIT; signal  \BRDIF/\   : AGCBIT;
  signal  \36422\    : AGCBIT; signal  \BR1B2B\   : AGCBIT;
  signal  \36423\    : AGCBIT; signal  \BR1B2B/\  : AGCBIT;
  signal  \36424\    : AGCBIT;
  signal  \36425\    : AGCBIT;
  signal \&36426\    : AGCBIT;
  signal  \36427\    : AGCBIT;
  signal \&36428\    : AGCBIT;
  signal  \36429\    : AGCBIT; signal  \4XP5\     : AGCBIT;
  signal \&36430\    : AGCBIT;
  signal  \36431\    : AGCBIT;
  signal  \36432\    : AGCBIT; signal  \8XP5\     : AGCBIT;
  signal  \36433\    : AGCBIT; signal  \4XP11\    : AGCBIT;
  signal  \36434\    : AGCBIT; signal  \8XP6\     : AGCBIT;
  signal  \36435\    : AGCBIT;
  signal  \36436\    : AGCBIT;
  signal  \36437\    : AGCBIT;
  signal  \36438\    : AGCBIT;
  signal  \36439\    : AGCBIT;
  signal \&36440\    : AGCBIT;
  signal \&36441\    : AGCBIT;
  signal \&36442\    : AGCBIT;
  signal  \36443\    : AGCBIT; signal  \B15X\     : AGCBIT;
  signal  \36444\    : AGCBIT;
  signal  \36445\    : AGCBIT; signal  \5XP4\     : AGCBIT;
  signal  \36446\    : AGCBIT;
  signal  \36447\    : AGCBIT; signal  \6XP5\     : AGCBIT;
  signal  \36448\    : AGCBIT; signal  \KRPT\     : AGCBIT;
  signal  \36449\    : AGCBIT; signal  \TL15\     : AGCBIT;
  signal  \36450\    : AGCBIT; signal  \MP0T10\   : AGCBIT;
  signal  \36451\    : AGCBIT;
  signal \&36452\    : AGCBIT;
  signal \&36453\    : AGCBIT;
  signal \&36454\    : AGCBIT;
  signal  \36455\    : AGCBIT; signal  \TSGN2\    : AGCBIT;
  signal  \36456\    : AGCBIT;
  signal  \36457\    : AGCBIT; signal  \7XP19\    : AGCBIT;
  signal \&36459\    : AGCBIT;
  signal \&36460\    : AGCBIT;
  signal  \39101\    : AGCBIT;
  signal  \39102\    : AGCBIT;
  signal  \39103\    : AGCBIT;
  signal \&39104\    : AGCBIT;
  signal  \39105\    : AGCBIT;
  signal  \39106\    : AGCBIT;
  signal \&39107\    : AGCBIT;
  signal  \39108\    : AGCBIT;
  signal  \39109\    : AGCBIT;
  signal \&39110\    : AGCBIT;
  signal  \39111\    : AGCBIT;
  signal  \39112\    : AGCBIT;
  signal  \39113\    : AGCBIT; signal  \NISQ/\    : AGCBIT;
  signal  \39115\    : AGCBIT; signal  \DVST\     : AGCBIT;
  signal  \39116\    : AGCBIT;
  signal  \39117\    : AGCBIT; signal  \2XP7\     : AGCBIT;
  signal  \39120\    : AGCBIT;
  signal  \39121\    : AGCBIT;
  signal  \39122\    : AGCBIT; signal  \3XP6\     : AGCBIT;
  signal \&39123\    : AGCBIT;
  signal  \39124\    : AGCBIT;
  signal  \39125\    : AGCBIT;
  signal  \39126\    : AGCBIT; signal  \TPZG/\    : AGCBIT;
  signal  \39127\    : AGCBIT;
  signal \&39128\    : AGCBIT;
  signal  \39129\    : AGCBIT;
  signal \&39130\    : AGCBIT;
  signal  \39131\    : AGCBIT;
  signal  \39132\    : AGCBIT; signal  \PARTC\    : AGCBIT;
  signal  \39133\    : AGCBIT;
  signal  \39134\    : AGCBIT;
  signal \&39135\    : AGCBIT;
  signal  \39136\    : AGCBIT; signal  \5XP12\    : AGCBIT;
  signal  \39137\    : AGCBIT; signal  \TSGN/\    : AGCBIT;
  signal  \39138\    : AGCBIT;
  signal \&39139\    : AGCBIT;
  signal  \39140\    : AGCBIT;
  signal \&39141\    : AGCBIT;
  signal  \39143\    : AGCBIT;
  signal \&39144\    : AGCBIT;
  signal  \39145\    : AGCBIT;
  signal \&39146\    : AGCBIT;
  signal  \39147\    : AGCBIT; signal  \7XP9\     : AGCBIT;
  signal \&39148\    : AGCBIT;
  signal  \39149\    : AGCBIT;
  signal  \39150\    : AGCBIT; signal  \7XP4\     : AGCBIT;
  signal  \39151\    : AGCBIT; signal  \PTWOX\    : AGCBIT;
  signal  \39152\    : AGCBIT;
  signal \&39153\    : AGCBIT;
  signal \&39154\    : AGCBIT;
  signal \&39155\    : AGCBIT;
  signal \&39156\    : AGCBIT;
  signal  \39201\    : AGCBIT;
  signal \&39202\    : AGCBIT;
  signal  \39203\    : AGCBIT;
  signal \&39204\    : AGCBIT;
  signal  \39205\    : AGCBIT; signal  \TSUDO/\   : AGCBIT;
  signal \&39206\    : AGCBIT;
  signal  \39207\    : AGCBIT; signal  \RAD\      : AGCBIT;
  signal \&39208\    : AGCBIT;
  signal  \39209\    : AGCBIT;
  signal  \39210\    : AGCBIT; signal  \8XP15\    : AGCBIT;
  signal  \39211\    : AGCBIT;
  signal  \39212\    : AGCBIT; signal  \8XP3\     : AGCBIT;
  signal  \39213\    : AGCBIT;
  signal  \39214\    : AGCBIT;
  signal \&39215\    : AGCBIT;
  signal  \39216\    : AGCBIT;
  signal  \39217\    : AGCBIT;
  signal  \39219\    : AGCBIT; signal  \RSTRT\    : AGCBIT;
  signal  \39220\    : AGCBIT; signal  \8XP12\    : AGCBIT;
  signal  \39221\    : AGCBIT;
  signal  \39222\    : AGCBIT;
  signal  \39223\    : AGCBIT;
  signal  \39224\    : AGCBIT; signal  \9XP5\     : AGCBIT;
  signal  \39225\    : AGCBIT;
  signal \&39226\    : AGCBIT;
  signal  \39227\    : AGCBIT;
  signal \&39228\    : AGCBIT;
  signal  \39229\    : AGCBIT; signal  \10XP6\    : AGCBIT;
  signal  \39230\    : AGCBIT;
  signal  \39231\    : AGCBIT; signal  \10XP1\    : AGCBIT;
  signal  \39232\    : AGCBIT;
  signal  \39233\    : AGCBIT;
  signal \&39234\    : AGCBIT;
  signal  \39235\    : AGCBIT;
  signal  \39236\    : AGCBIT; signal  \10XP7\    : AGCBIT;
  signal  \39237\    : AGCBIT;
  signal  \39238\    : AGCBIT; signal  \10XP8\    : AGCBIT;
  signal  \39239\    : AGCBIT;
  signal  \39240\    : AGCBIT; signal  \11XP2\    : AGCBIT;
  signal  \39241\    : AGCBIT;
  signal \&39242\    : AGCBIT;
  signal  \39243\    : AGCBIT;
  signal \&39244\    : AGCBIT;
  signal  \39245\    : AGCBIT;
  signal  \39248\    : AGCBIT;
  signal  \39249\    : AGCBIT; signal  \GNHNC\    : AGCBIT;
  signal \$39249\    : AGCBIT;
  signal  \39250\    : AGCBIT;
  signal \&39251\    : AGCBIT;
  signal \&39252\    : AGCBIT;
  signal \&39253\    : AGCBIT;
  signal  \39254\    : AGCBIT;
  signal  \39255\    : AGCBIT; signal  \PINC/\    : AGCBIT;
  signal \$39255\    : AGCBIT;
  signal  \39256\    : AGCBIT; signal  \PINC\     : AGCBIT;
  signal \&39261\    : AGCBIT;
  signal  \39301\    : AGCBIT;
  signal \&39302\    : AGCBIT;
  signal \&39303\    : AGCBIT;
  signal  \39304\    : AGCBIT; signal  \RL10BB\   : AGCBIT;
  signal \&39305\    : AGCBIT;
  signal  \39306\    : AGCBIT; signal  \R6\       : AGCBIT;
  signal  \39307\    : AGCBIT;
  signal  \39308\    : AGCBIT; signal  \2XP8\     : AGCBIT;
  signal  \39309\    : AGCBIT; signal  \RSCT\     : AGCBIT;
  signal  \39310\    : AGCBIT;
  signal \&39311\    : AGCBIT;
  signal  \39312\    : AGCBIT;
  signal  \39313\    : AGCBIT;
  signal  \39314\    : AGCBIT; signal  \RQ\       : AGCBIT;
  signal \&39315\    : AGCBIT;
  signal \&39316\    : AGCBIT;
  signal  \39318\    : AGCBIT;
  signal  \39319\    : AGCBIT;
  signal  \39320\    : AGCBIT;
  signal  \39321\    : AGCBIT; signal  \RL/\      : AGCBIT;
  signal  \39322\    : AGCBIT; signal  \RA/\      : AGCBIT;
  signal  \39323\    : AGCBIT; signal  \TRSM\     : AGCBIT;
  signal  \39324\    : AGCBIT;
  signal \&39325\    : AGCBIT;
  signal \&39326\    : AGCBIT;
  signal  \39327\    : AGCBIT;
  signal \&39328\    : AGCBIT;
  signal  \39329\    : AGCBIT;
  signal  \39330\    : AGCBIT;
  signal  \39331\    : AGCBIT; signal  \WY12/\    : AGCBIT;
  signal  \39332\    : AGCBIT; signal  \5XP9\     : AGCBIT;
  signal  \39333\    : AGCBIT; signal  \WY/\      : AGCBIT;
  signal \&39334\    : AGCBIT;
  signal  \39335\    : AGCBIT;
  signal \&39336\    : AGCBIT;
  signal  \39337\    : AGCBIT; signal  \5XP13\    : AGCBIT;
  signal \&39338\    : AGCBIT;
  signal  \39339\    : AGCBIT; signal  \5XP15\    : AGCBIT;
  signal  \39340\    : AGCBIT; signal  \5XP21\    : AGCBIT;
  signal  \39341\    : AGCBIT;
  signal  \39342\    : AGCBIT;
  signal  \39343\    : AGCBIT;
  signal  \39344\    : AGCBIT;
  signal \&39345\    : AGCBIT;
  signal  \39346\    : AGCBIT; signal  \SCAD\     : AGCBIT;
  signal  \39347\    : AGCBIT; signal  \SCAD/\    : AGCBIT;
  signal  \39348\    : AGCBIT;
  signal \&39349\    : AGCBIT;
  signal  \39350\    : AGCBIT; signal  \NDR100/\  : AGCBIT;
  signal  \39352\    : AGCBIT; signal  \OCTAD2\   : AGCBIT;
  signal  \39353\    : AGCBIT; signal  \OCTAD3\   : AGCBIT;
  signal  \39354\    : AGCBIT; signal  \OCTAD4\   : AGCBIT;
  signal  \39355\    : AGCBIT; signal  \OCTAD5\   : AGCBIT;
  signal  \39356\    : AGCBIT; signal  \OCTAD6\   : AGCBIT;
  signal  \39401\    : AGCBIT;
  signal  \39402\    : AGCBIT; signal  \DV1B1B\   : AGCBIT;
  signal  \39403\    : AGCBIT;
  signal  \39404\    : AGCBIT;
  signal  \39405\    : AGCBIT;
  signal  \39406\    : AGCBIT;
  signal  \39407\    : AGCBIT; signal  \5XP19\    : AGCBIT;
  signal  \39408\    : AGCBIT;
  signal  \39409\    : AGCBIT;
  signal \&39410\    : AGCBIT;
  signal  \39411\    : AGCBIT;
  signal  \39412\    : AGCBIT;
  signal \&39413\    : AGCBIT;
  signal \&39414\    : AGCBIT;
  signal  \39415\    : AGCBIT;
  signal  \39416\    : AGCBIT;
  signal \&39417\    : AGCBIT;
  signal \&39418\    : AGCBIT;
  signal  \39419\    : AGCBIT; signal  \6XP8\     : AGCBIT;
  signal  \39420\    : AGCBIT; signal  \6XP7\     : AGCBIT;
  signal  \39421\    : AGCBIT; signal  \6XP2\     : AGCBIT;
  signal \&39422\    : AGCBIT;
  signal \&39423\    : AGCBIT;
  signal \&39424\    : AGCBIT;
  signal  \39425\    : AGCBIT;
  signal  \39426\    : AGCBIT; signal  \U2BBK\    : AGCBIT;
  signal  \39427\    : AGCBIT;
  signal  \39428\    : AGCBIT;
  signal \&39429\    : AGCBIT;
  signal \&39430\    : AGCBIT;
  signal  \39431\    : AGCBIT; signal  \RSTSTG\   : AGCBIT;
  signal  \39432\    : AGCBIT;
  signal \&39433\    : AGCBIT;
  signal \&39434\    : AGCBIT;
  signal \&39435\    : AGCBIT;
  signal  \39436\    : AGCBIT;
  signal \&39437\    : AGCBIT;
  signal \&39438\    : AGCBIT;
  signal  \39439\    : AGCBIT;
  signal  \39440\    : AGCBIT; signal  \TMZ/\     : AGCBIT;
  signal  \39441\    : AGCBIT;
  signal  \39442\    : AGCBIT; signal  \10XP10\   : AGCBIT;
  signal \&39443\    : AGCBIT;
  signal \&39444\    : AGCBIT;
  signal  \39445\    : AGCBIT;
  signal  \39446\    : AGCBIT; signal  \DV4B1B\   : AGCBIT;
  signal  \39447\    : AGCBIT;
  signal  \39448\    : AGCBIT;
  signal  \39449\    : AGCBIT;
  signal  \39450\    : AGCBIT; signal  \11XP6\    : AGCBIT;
  signal  \39451\    : AGCBIT;
  signal  \39452\    : AGCBIT;
  signal  \40101\    : AGCBIT;
  signal  \40102\    : AGCBIT;
  signal  \40103\    : AGCBIT;
  signal  \40104\    : AGCBIT;
  signal  \40105\    : AGCBIT;
  signal  \40106\    : AGCBIT; signal  \DVXP1\    : AGCBIT;
  signal  \40107\    : AGCBIT; signal  \A2X/\     : AGCBIT;
  signal  \40108\    : AGCBIT; signal  \L2GD/\    : AGCBIT;
  signal  \40109\    : AGCBIT; signal  \RB/\      : AGCBIT;
  signal  \40110\    : AGCBIT; signal  \WYD/\     : AGCBIT;
  signal  \40111\    : AGCBIT;
  signal \&40112\    : AGCBIT;
  signal  \40113\    : AGCBIT;
  signal  \40114\    : AGCBIT;
  signal  \40115\    : AGCBIT;
  signal  \40116\    : AGCBIT;
  signal  \40117\    : AGCBIT; signal  \ZIP\      : AGCBIT;
  signal  \40118\    : AGCBIT;
  signal \&40119\    : AGCBIT;
  signal  \40120\    : AGCBIT;
  signal  \40121\    : AGCBIT;
  signal  \40122\    : AGCBIT;
  signal  \40123\    : AGCBIT;
  signal  \40124\    : AGCBIT;
  signal  \40125\    : AGCBIT;
  signal  \40126\    : AGCBIT;
  signal  \40127\    : AGCBIT;
  signal  \40128\    : AGCBIT;
  signal  \40129\    : AGCBIT;
  signal  \40130\    : AGCBIT; signal  \ZIPCI\    : AGCBIT;
  signal  \40131\    : AGCBIT; signal  \RC/\      : AGCBIT;
  signal  \40132\    : AGCBIT; signal  \RCH/\     : AGCBIT;
  signal  \40133\    : AGCBIT;
  signal  \40134\    : AGCBIT;
  signal  \40135\    : AGCBIT;
  signal  \40136\    : AGCBIT;
  signal  \40137\    : AGCBIT;
  signal  \40138\    : AGCBIT;
  signal  \40139\    : AGCBIT; signal  \TSGU/\    : AGCBIT;
  signal  \40140\    : AGCBIT; signal  \WL/\      : AGCBIT;
  signal \&40141\    : AGCBIT;
  signal  \40142\    : AGCBIT;
  signal  \40143\    : AGCBIT;
  signal  \40144\    : AGCBIT;
  signal  \40145\    : AGCBIT;
  signal  \40146\    : AGCBIT; signal  \RG/\      : AGCBIT;
  signal  \40147\    : AGCBIT;
  signal \&40148\    : AGCBIT;
  signal  \40149\    : AGCBIT;
  signal  \40150\    : AGCBIT;
  signal  \40151\    : AGCBIT;
  signal  \40152\    : AGCBIT; signal  \ZAP/\     : AGCBIT;
  signal \&40153\    : AGCBIT;
  signal  \40154\    : AGCBIT; signal  \ZAP\      : AGCBIT;
  signal  \40155\    : AGCBIT; signal  \WB/\      : AGCBIT;
  signal  \40156\    : AGCBIT; signal  \RU/\      : AGCBIT;
  signal \&40157\    : AGCBIT;
  signal  \40158\    : AGCBIT; signal  \WZ/\      : AGCBIT;
  signal  \40160\    : AGCBIT; signal  \MCRO/\    : AGCBIT;
  signal  \40201\    : AGCBIT; signal  \RB1F\     : AGCBIT;
  signal  \40202\    : AGCBIT; signal  \CLXC\     : AGCBIT;
  signal \&40203\    : AGCBIT;
  signal \&40204\    : AGCBIT;
  signal  \40206\    : AGCBIT; signal  \WQ/\      : AGCBIT;
  signal  \40207\    : AGCBIT; signal  \TOV/\     : AGCBIT;
  signal  \40208\    : AGCBIT; signal  \WSC/\     : AGCBIT;
  signal  \40209\    : AGCBIT; signal  \WG/\      : AGCBIT;
  signal  \40210\    : AGCBIT; signal  \MONEX\    : AGCBIT;
  signal  \40213\    : AGCBIT;
  signal  \40214\    : AGCBIT; signal  \TWOX\     : AGCBIT;
  signal  \40215\    : AGCBIT;
  signal  \40216\    : AGCBIT; signal  \BXVX\     : AGCBIT;
  signal  \40217\    : AGCBIT;
  signal  \40220\    : AGCBIT; signal  \PIFL/\    : AGCBIT;
  signal \$40220\    : AGCBIT;
  signal  \40221\    : AGCBIT;
  signal  \40222\    : AGCBIT;
  signal \&40224\    : AGCBIT;
  signal \&40225\    : AGCBIT;
  signal \&40226\    : AGCBIT;
  signal \&40227\    : AGCBIT;
  signal \&40228\    : AGCBIT;
  signal \&40229\    : AGCBIT;
  signal \&40230\    : AGCBIT;
  signal \&40231\    : AGCBIT;
  signal \&40232\    : AGCBIT;
  signal \&40233\    : AGCBIT;
  signal \&40234\    : AGCBIT;
  signal \&40235\    : AGCBIT;
  signal \&40236\    : AGCBIT;
  signal \&40237\    : AGCBIT;
  signal \&40238\    : AGCBIT;
  signal \&40239\    : AGCBIT;
  signal  \40240\    : AGCBIT;
  signal  \40241\    : AGCBIT; signal  \CGMC\     : AGCBIT;
  signal  \40242\    : AGCBIT;
  signal \$40242\    : AGCBIT;
  signal  \40243\    : AGCBIT;
  signal  \40244\    : AGCBIT;
  signal \$40244\    : AGCBIT;
  signal  \40245\    : AGCBIT;
  signal \$40245\    : AGCBIT;
  signal  \40246\    : AGCBIT;
  signal \$40246\    : AGCBIT;
  signal  \40247\    : AGCBIT;
  signal  \40248\    : AGCBIT;
  signal \&40249\    : AGCBIT;
  signal  \40250\    : AGCBIT;
  signal  \40251\    : AGCBIT; signal  \TIMR\     : AGCBIT;
  signal  \40253\    : AGCBIT;
  signal \$40253\    : AGCBIT;
  signal  \40254\    : AGCBIT;
  signal \$40254\    : AGCBIT;
  signal  \40255\    : AGCBIT;
  signal \$40255\    : AGCBIT;
  signal  \40256\    : AGCBIT;
  signal \$40256\    : AGCBIT;
  signal  \40257\    : AGCBIT;
  signal \$40257\    : AGCBIT;
  signal  \40258\    : AGCBIT;
  signal \$40258\    : AGCBIT;
  signal  \40302\    : AGCBIT;
  signal  \40303\    : AGCBIT;
  signal  \40304\    : AGCBIT;
  signal  \40305\    : AGCBIT; signal  \6XP10\    : AGCBIT;
  signal \&40306\    : AGCBIT;
  signal  \40307\    : AGCBIT;
  signal  \40309\    : AGCBIT;
  signal  \40310\    : AGCBIT;
  signal  \40311\    : AGCBIT; signal  \MONEX/\   : AGCBIT;
  signal  \40312\    : AGCBIT;
  signal  \40313\    : AGCBIT;
  signal  \40314\    : AGCBIT;
  signal \&40315\    : AGCBIT;
  signal  \40317\    : AGCBIT;
  signal  \40318\    : AGCBIT;
  signal  \40320\    : AGCBIT; signal  \POUT\     : AGCBIT;
  signal  \40321\    : AGCBIT; signal  \MOUT\     : AGCBIT;
  signal  \40322\    : AGCBIT; signal  \ZOUT\     : AGCBIT;
  signal  \40323\    : AGCBIT;
  signal  \40324\    : AGCBIT;
  signal  \40325\    : AGCBIT;
  signal  \40326\    : AGCBIT;
  signal  \40327\    : AGCBIT; signal  \7XP7\     : AGCBIT;
  signal \&40328\    : AGCBIT;
  signal  \40329\    : AGCBIT;
  signal  \40330\    : AGCBIT;
  signal  \40331\    : AGCBIT; signal  \7XP14\    : AGCBIT;
  signal  \40333\    : AGCBIT;
  signal  \40334\    : AGCBIT;
  signal  \40335\    : AGCBIT;
  signal  \40336\    : AGCBIT;
  signal  \40337\    : AGCBIT;
  signal  \40338\    : AGCBIT;
  signal \&40339\    : AGCBIT;
  signal  \40340\    : AGCBIT;
  signal  \40341\    : AGCBIT; signal  \WOVR\     : AGCBIT;
  signal \&40342\    : AGCBIT;
  signal \&40343\    : AGCBIT;
  signal \&40344\    : AGCBIT;
  signal  \40345\    : AGCBIT;
  signal  \40346\    : AGCBIT;
  signal \&40347\    : AGCBIT;
  signal \&40348\    : AGCBIT;
  signal  \40349\    : AGCBIT; signal  \8XP4\     : AGCBIT;
  signal  \40350\    : AGCBIT; signal  \8XP10\    : AGCBIT;
  signal \&40351\    : AGCBIT;
  signal  \40352\    : AGCBIT;
  signal  \40353\    : AGCBIT;
  signal  \40354\    : AGCBIT;
  signal  \40355\    : AGCBIT;
  signal \&40356\    : AGCBIT;
  signal  \40357\    : AGCBIT; signal  \RD_BANK\  : AGCBIT;
  signal \&40358\    : AGCBIT;
  signal  \40401\    : AGCBIT;
  signal  \40402\    : AGCBIT; signal  \EXT\      : AGCBIT;
  signal  \40403\    : AGCBIT; signal  \10XP9\    : AGCBIT;
  signal  \40405\    : AGCBIT;
  signal \&40406\    : AGCBIT;
  signal  \40407\    : AGCBIT;
  signal  \40408\    : AGCBIT;
  signal  \40409\    : AGCBIT;
  signal  \40410\    : AGCBIT;
  signal  \40411\    : AGCBIT;
  signal \&40412\    : AGCBIT;
  signal  \40413\    : AGCBIT;
  signal  \40414\    : AGCBIT; signal  \WA/\      : AGCBIT;
  signal \&40415\    : AGCBIT;
  signal \&40416\    : AGCBIT;
  signal \&40417\    : AGCBIT;
  signal \&40418\    : AGCBIT;
  signal  \40419\    : AGCBIT; signal  \RUS/\     : AGCBIT;
  signal  \40420\    : AGCBIT; signal  \RZ/\      : AGCBIT;
  signal \&40421\    : AGCBIT;
  signal  \40422\    : AGCBIT;
  signal  \40423\    : AGCBIT; signal  \ST1\      : AGCBIT;
  signal  \40424\    : AGCBIT; signal  \ST2/\     : AGCBIT;
  signal  \40425\    : AGCBIT; signal  \ST2\      : AGCBIT;
  signal  \40426\    : AGCBIT;
  signal \$40426\    : AGCBIT;
  signal  \40427\    : AGCBIT; signal  \NEAC\     : AGCBIT;
  signal \&40428\    : AGCBIT;
  signal  \40430\    : AGCBIT; signal  \WS/\      : AGCBIT;
  signal  \40431\    : AGCBIT; signal  \CI/\      : AGCBIT;
  signal  \40432\    : AGCBIT;
  signal \&40433\    : AGCBIT;
  signal  \40434\    : AGCBIT; signal  \PONEX\    : AGCBIT;
  signal  \40435\    : AGCBIT; signal  \R1C/\     : AGCBIT;
  signal  \40436\    : AGCBIT; signal  \RB1/\     : AGCBIT;
  signal  \40438\    : AGCBIT;
  signal  \40439\    : AGCBIT;
  signal \$40439\    : AGCBIT;
  signal  \40440\    : AGCBIT; signal  \PSEUDO\   : AGCBIT;
  signal \&40441\    : AGCBIT;
  signal  \33101\    : AGCBIT; signal  \WALSG/\   : AGCBIT;
  signal  \33102\    : AGCBIT; signal  \WALSG\    : AGCBIT;
  signal  \33105\    : AGCBIT;
  signal  \33106\    : AGCBIT;
  signal  \33107\    : AGCBIT;
  signal  \33108\    : AGCBIT;
  signal  \33109\    : AGCBIT; signal  \WYLOG/\   : AGCBIT;
  signal  \33111\    : AGCBIT;
  signal  \33112\    : AGCBIT; signal  \WYHIG/\   : AGCBIT;
  signal  \33113\    : AGCBIT;
  signal \&33114\    : AGCBIT;
  signal \&33115\    : AGCBIT;
  signal  \33116\    : AGCBIT; signal  \CUG\      : AGCBIT;
  signal  \33122\    : AGCBIT;
  signal \&33123\    : AGCBIT;
  signal  \33124\    : AGCBIT;
  signal  \33125\    : AGCBIT;
  signal  \33126\    : AGCBIT; signal  \WYDG/\    : AGCBIT;
  signal  \33129\    : AGCBIT; signal  \WYDLOG/\  : AGCBIT;
  signal  \33130\    : AGCBIT;
  signal  \33131\    : AGCBIT; signal  \WBG/\     : AGCBIT;
  signal \&33135\    : AGCBIT;
  signal  \33136\    : AGCBIT; signal  \CBG\      : AGCBIT;
  signal \&33138\    : AGCBIT;
  signal \&33139\    : AGCBIT;
  signal  \33140\    : AGCBIT; signal  \WGNORM\   : AGCBIT;
  signal  \33141\    : AGCBIT; signal  \WG1G/\    : AGCBIT;
  signal  \33144\    : AGCBIT;
  signal  \33145\    : AGCBIT; signal  \WG2G/\    : AGCBIT;
  signal  \33146\    : AGCBIT; signal  \WG4G/\    : AGCBIT;
  signal  \33149\    : AGCBIT;
  signal  \33150\    : AGCBIT; signal  \WG5G/\    : AGCBIT;
  signal  \33151\    : AGCBIT;
  signal  \33152\    : AGCBIT; signal  \WG3G/\    : AGCBIT;
  signal  \33155\    : AGCBIT;
  signal  \33156\    : AGCBIT; signal  \WEDOPG/\  : AGCBIT;
  signal  \33160\    : AGCBIT; signal  \PIPSAM\   : AGCBIT;
  signal  \33201\    : AGCBIT;
  signal  \33202\    : AGCBIT; signal  \WZG/\     : AGCBIT;
  signal  \33204\    : AGCBIT;
  signal \&33207\    : AGCBIT;
  signal  \33208\    : AGCBIT; signal  \CZG\      : AGCBIT;
  signal  \33211\    : AGCBIT;
  signal  \33212\    : AGCBIT;
  signal  \33213\    : AGCBIT;
  signal  \33214\    : AGCBIT; signal  \WLG/\     : AGCBIT;
  signal  \33217\    : AGCBIT;
  signal \&33218\    : AGCBIT;
  signal  \33219\    : AGCBIT;
  signal \&33220\    : AGCBIT;
  signal  \33221\    : AGCBIT; signal  \CLG2G\    : AGCBIT;
  signal  \33222\    : AGCBIT;
  signal \&33223\    : AGCBIT;
  signal  \33224\    : AGCBIT; signal  \CLG1G\    : AGCBIT;
  signal  \33227\    : AGCBIT;
  signal  \33228\    : AGCBIT;
  signal  \33229\    : AGCBIT; signal  \WAG/\     : AGCBIT;
  signal  \33232\    : AGCBIT;
  signal  \33233\    : AGCBIT;
  signal  \33234\    : AGCBIT; signal  \CAG\      : AGCBIT;
  signal  \33237\    : AGCBIT;
  signal  \33238\    : AGCBIT; signal  \WSG/\     : AGCBIT;
  signal \&33241\    : AGCBIT;
  signal  \33242\    : AGCBIT; signal  \CSG\      : AGCBIT;
  signal  \33244\    : AGCBIT;
  signal  \33245\    : AGCBIT;
  signal  \33246\    : AGCBIT;
  signal  \33247\    : AGCBIT; signal  \WQG/\     : AGCBIT;
  signal \&33251\    : AGCBIT;
  signal  \33252\    : AGCBIT; signal  \CQG\      : AGCBIT;
  signal \&33255\    : AGCBIT;
  signal  \33257\    : AGCBIT; signal  \P04A\     : AGCBIT;
  signal  \33301\    : AGCBIT;
  signal  \33302\    : AGCBIT; signal  \WEBG/\    : AGCBIT;
  signal \&33303\    : AGCBIT;
  signal  \33305\    : AGCBIT;
  signal  \33306\    : AGCBIT; signal  \CEBG\     : AGCBIT;
  signal  \33307\    : AGCBIT;
  signal  \33308\    : AGCBIT; signal  \WFBG/\    : AGCBIT;
  signal  \33310\    : AGCBIT; signal  \CFBG\     : AGCBIT;
  signal \&33311\    : AGCBIT;
  signal  \33312\    : AGCBIT;
  signal  \33313\    : AGCBIT; signal  \WBBEG/\   : AGCBIT;
  signal \&33315\    : AGCBIT;
  signal  \33316\    : AGCBIT; signal  \RGG1\     : AGCBIT;
  signal  \33317\    : AGCBIT; signal  \RGG/\     : AGCBIT;
  signal \&33320\    : AGCBIT;
  signal  \33321\    : AGCBIT;
  signal  \33322\    : AGCBIT;
  signal  \33323\    : AGCBIT; signal  \RAG/\     : AGCBIT;
  signal \&33326\    : AGCBIT;
  signal  \33327\    : AGCBIT;
  signal  \33328\    : AGCBIT; signal  \REBG/\    : AGCBIT;
  signal  \33329\    : AGCBIT; signal  \RLG2\     : AGCBIT;
  signal  \33330\    : AGCBIT; signal  \RLG/\     : AGCBIT;
  signal  \33331\    : AGCBIT; signal  \RLG1\     : AGCBIT;
  signal  \33333\    : AGCBIT; signal  \RLG3\     : AGCBIT;
  signal \&33335\    : AGCBIT;
  signal  \33336\    : AGCBIT;
  signal  \33337\    : AGCBIT;
  signal  \33338\    : AGCBIT; signal  \RZG/\     : AGCBIT;
  signal  \33341\    : AGCBIT;
  signal  \33342\    : AGCBIT; signal  \RULOG/\   : AGCBIT;
  signal  \33345\    : AGCBIT;
  signal  \33346\    : AGCBIT;
  signal \&33347\    : AGCBIT;
  signal  \33348\    : AGCBIT; signal  \RUG/\     : AGCBIT;
  signal  \33349\    : AGCBIT; signal  \RUSG/\    : AGCBIT;
  signal  \33350\    : AGCBIT;
  signal  \33351\    : AGCBIT; signal  \RBHG/\    : AGCBIT;
  signal  \33352\    : AGCBIT;
  signal  \33353\    : AGCBIT; signal  \RBLG/\    : AGCBIT;
  signal  \33355\    : AGCBIT;
  signal  \33356\    : AGCBIT; signal  \CI01/\    : AGCBIT;
  signal \$33356\    : AGCBIT;
  signal  \33359\    : AGCBIT;
  signal  \33401\    : AGCBIT;
  signal  \33402\    : AGCBIT; signal  \RCG/\     : AGCBIT;
  signal  \33405\    : AGCBIT;
  signal  \33406\    : AGCBIT; signal  \RQG/\     : AGCBIT;
  signal  \33407\    : AGCBIT;
  signal  \33409\    : AGCBIT;
  signal  \33411\    : AGCBIT;
  signal  \33412\    : AGCBIT; signal  \RFBG/\    : AGCBIT;
  signal  \33413\    : AGCBIT;
  signal  \33414\    : AGCBIT; signal  \RBBEG/\   : AGCBIT;
  signal  \33415\    : AGCBIT; signal  \G2LSG\    : AGCBIT;
  signal  \33416\    : AGCBIT; signal  \G2LSG/\   : AGCBIT;
  signal  \33419\    : AGCBIT;
  signal  \33420\    : AGCBIT; signal  \L2GDG/\   : AGCBIT;
  signal  \33423\    : AGCBIT;
  signal  \33424\    : AGCBIT; signal  \A2XG/\    : AGCBIT;
  signal  \33427\    : AGCBIT;
  signal  \33428\    : AGCBIT;
  signal  \33429\    : AGCBIT;
  signal  \33430\    : AGCBIT; signal  \CGG\      : AGCBIT;
  signal  \33433\    : AGCBIT; signal  \YT0\      : AGCBIT;
  signal  \33434\    : AGCBIT; signal  \YT0/\     : AGCBIT;
  signal \&33435\    : AGCBIT;
  signal  \33436\    : AGCBIT; signal  \YT1\      : AGCBIT;
  signal  \33437\    : AGCBIT; signal  \YT1/\     : AGCBIT;
  signal \&33438\    : AGCBIT;
  signal  \33439\    : AGCBIT; signal  \YT2\      : AGCBIT;
  signal  \33440\    : AGCBIT; signal  \YT2/\     : AGCBIT;
  signal \&33441\    : AGCBIT;
  signal  \33442\    : AGCBIT; signal  \YT3\      : AGCBIT;
  signal  \33443\    : AGCBIT; signal  \YT3/\     : AGCBIT;
  signal \&33444\    : AGCBIT;
  signal  \33445\    : AGCBIT; signal  \YT4\      : AGCBIT;
  signal  \33446\    : AGCBIT; signal  \YT4/\     : AGCBIT;
  signal \&33447\    : AGCBIT;
  signal  \33448\    : AGCBIT; signal  \YT5\      : AGCBIT;
  signal  \33449\    : AGCBIT; signal  \YT5/\     : AGCBIT;
  signal \&33450\    : AGCBIT;
  signal  \33451\    : AGCBIT; signal  \YT6\      : AGCBIT;
  signal  \33452\    : AGCBIT; signal  \YT6/\     : AGCBIT;
  signal \&33453\    : AGCBIT;
  signal  \33454\    : AGCBIT; signal  \YT7\      : AGCBIT;
  signal  \33455\    : AGCBIT; signal  \YT7/\     : AGCBIT;
  signal \&33456\    : AGCBIT;
  signal  \33457\    : AGCBIT; signal  \CINORM\   : AGCBIT;
  signal  \33458\    : AGCBIT;
  signal \$33458\    : AGCBIT;
  signal  \33459\    : AGCBIT; signal  \CIFF\     : AGCBIT;
  signal  \33460\    : AGCBIT; signal  \RBBK\     : AGCBIT;
  signal  \51101\    : AGCBIT; signal  \CO04\     : AGCBIT;
  signal  \51102\    : AGCBIT;
  signal  \51103\    : AGCBIT;
  signal \$51103\    : AGCBIT;
  signal  \51104\    : AGCBIT;
  signal  \51105\    : AGCBIT;
  signal  \51106\    : AGCBIT;
  signal  \51107\    : AGCBIT;
  signal \$51107\    : AGCBIT;
  signal  \51108\    : AGCBIT;
  signal  \51109\    : AGCBIT;
  signal  \51110\    : AGCBIT; signal  \XUY01/\   : AGCBIT;
  signal  \51111\    : AGCBIT;
  signal  \51112\    : AGCBIT; signal  \SUMA01/\  : AGCBIT;
  signal  \51113\    : AGCBIT;
  signal  \51114\    : AGCBIT; signal  \CI02/\    : AGCBIT;
  signal  \51115\    : AGCBIT; signal  \SUMB01/\  : AGCBIT;
  signal  \51117\    : AGCBIT;
  signal  \51118\    : AGCBIT;
  signal  \51119\    : AGCBIT;
  signal  \51120\    : AGCBIT; signal  \A01/\     : AGCBIT;
  signal \$51120\    : AGCBIT;
  signal  \51121\    : AGCBIT;
  signal  \51122\    : AGCBIT;
  signal \&51123\    : AGCBIT;
  signal  \51124\    : AGCBIT;
  signal  \51125\    : AGCBIT;
  signal  \51126\    : AGCBIT; signal  \L01/\     : AGCBIT;
  signal \$51126\    : AGCBIT;
  signal  \51127\    : AGCBIT;
  signal  \51128\    : AGCBIT;
  signal  \51129\    : AGCBIT;
  signal  \51130\    : AGCBIT;
  signal \$51130\    : AGCBIT;
  signal  \51131\    : AGCBIT;
  signal  \51132\    : AGCBIT;
  signal \&51133\    : AGCBIT;
  signal  \51134\    : AGCBIT;
  signal  \51135\    : AGCBIT; signal  \Z01/\     : AGCBIT;
  signal \$51135\    : AGCBIT;
  signal  \51136\    : AGCBIT;
  signal  \51137\    : AGCBIT;
  signal  \51138\    : AGCBIT;
  signal  \51139\    : AGCBIT;
  signal \$51139\    : AGCBIT;
  signal  \51140\    : AGCBIT;
  signal  \51141\    : AGCBIT;
  signal  \51142\    : AGCBIT;
  signal  \51143\    : AGCBIT;
  signal  \51144\    : AGCBIT;
  signal  \51145\    : AGCBIT;
  signal  \51146\    : AGCBIT;
  signal \&51147\    : AGCBIT;
  signal  \51148\    : AGCBIT; signal  \G01/\     : AGCBIT;
  signal \$51148\    : AGCBIT;
  signal  \51149\    : AGCBIT; signal  \G01\      : AGCBIT;
  signal \&51150\    : AGCBIT;
  signal  \51151\    : AGCBIT;
  signal  \51152\    : AGCBIT; signal  \WL01\     : AGCBIT;
  signal \&51153\    : AGCBIT;
  signal  \51154\    : AGCBIT; signal  \WL01/\    : AGCBIT;
  signal  \51157\    : AGCBIT; signal  \RL01/\    : AGCBIT;
  signal \&51158\    : AGCBIT;
  signal  \51161\    : AGCBIT; signal  \CLEARA\   : AGCBIT;
  signal \&51162\    : AGCBIT;
  signal \&51163\    : AGCBIT;
  signal \&51201\    : AGCBIT;
  signal  \51202\    : AGCBIT;
  signal  \51203\    : AGCBIT;
  signal \$51203\    : AGCBIT;
  signal  \51204\    : AGCBIT;
  signal  \51205\    : AGCBIT;
  signal  \51206\    : AGCBIT;
  signal  \51207\    : AGCBIT;
  signal \$51207\    : AGCBIT;
  signal  \51208\    : AGCBIT;
  signal  \51209\    : AGCBIT;
  signal  \51210\    : AGCBIT; signal  \XUY02/\   : AGCBIT;
  signal  \51211\    : AGCBIT;
  signal  \51212\    : AGCBIT; signal  \SUMA02/\  : AGCBIT;
  signal  \51213\    : AGCBIT;
  signal  \51214\    : AGCBIT; signal  \CI03/\    : AGCBIT;
  signal  \51215\    : AGCBIT; signal  \SUMB02/\  : AGCBIT;
  signal  \51217\    : AGCBIT;
  signal  \51218\    : AGCBIT;
  signal  \51219\    : AGCBIT;
  signal  \51220\    : AGCBIT; signal  \A02/\     : AGCBIT;
  signal \$51220\    : AGCBIT;
  signal  \51221\    : AGCBIT;
  signal  \51222\    : AGCBIT;
  signal \&51223\    : AGCBIT;
  signal  \51224\    : AGCBIT;
  signal  \51225\    : AGCBIT;
  signal  \51226\    : AGCBIT; signal  \L02/\     : AGCBIT;
  signal \$51226\    : AGCBIT;
  signal  \51227\    : AGCBIT;
  signal  \51228\    : AGCBIT;
  signal  \51229\    : AGCBIT;
  signal  \51230\    : AGCBIT;
  signal \$51230\    : AGCBIT;
  signal  \51231\    : AGCBIT;
  signal  \51232\    : AGCBIT;
  signal \&51233\    : AGCBIT;
  signal  \51234\    : AGCBIT;
  signal  \51235\    : AGCBIT; signal  \Z02/\     : AGCBIT;
  signal \$51235\    : AGCBIT;
  signal  \51236\    : AGCBIT;
  signal  \51237\    : AGCBIT;
  signal  \51238\    : AGCBIT;
  signal  \51239\    : AGCBIT;
  signal \$51239\    : AGCBIT;
  signal  \51240\    : AGCBIT;
  signal  \51241\    : AGCBIT;
  signal  \51242\    : AGCBIT;
  signal  \51243\    : AGCBIT;
  signal  \51244\    : AGCBIT;
  signal  \51245\    : AGCBIT;
  signal  \51246\    : AGCBIT;
  signal \&51247\    : AGCBIT;
  signal  \51248\    : AGCBIT; signal  \G02/\     : AGCBIT;
  signal \$51248\    : AGCBIT;
  signal  \51249\    : AGCBIT; signal  \G02\      : AGCBIT;
  signal \&51250\    : AGCBIT;
  signal  \51251\    : AGCBIT;
  signal  \51252\    : AGCBIT; signal  \WL02\     : AGCBIT;
  signal \&51253\    : AGCBIT;
  signal  \51254\    : AGCBIT; signal  \WL02/\    : AGCBIT;
  signal  \51257\    : AGCBIT; signal  \RL02/\    : AGCBIT;
  signal \&51258\    : AGCBIT;
  signal  \51261\    : AGCBIT; signal  \S08A/\    : AGCBIT;
  signal  \51262\    : AGCBIT; signal  \S08A\     : AGCBIT;
  signal \&51263\    : AGCBIT;
  signal \&51301\    : AGCBIT;
  signal  \51302\    : AGCBIT;
  signal  \51303\    : AGCBIT;
  signal \$51303\    : AGCBIT;
  signal  \51304\    : AGCBIT;
  signal  \51305\    : AGCBIT;
  signal  \51306\    : AGCBIT;
  signal  \51307\    : AGCBIT;
  signal \$51307\    : AGCBIT;
  signal  \51308\    : AGCBIT;
  signal  \51309\    : AGCBIT;
  signal  \51310\    : AGCBIT; signal  \XUY04/\   : AGCBIT;
  signal  \51311\    : AGCBIT;
  signal  \51312\    : AGCBIT; signal  \SUMA04/\  : AGCBIT;
  signal  \51313\    : AGCBIT;
  signal  \51314\    : AGCBIT; signal  \CI05/\    : AGCBIT;
  signal  \51315\    : AGCBIT; signal  \SUMB04/\  : AGCBIT;
  signal  \51317\    : AGCBIT;
  signal  \51318\    : AGCBIT;
  signal  \51319\    : AGCBIT;
  signal  \51320\    : AGCBIT; signal  \A04/\     : AGCBIT;
  signal \$51320\    : AGCBIT;
  signal  \51321\    : AGCBIT;
  signal  \51322\    : AGCBIT;
  signal \&51323\    : AGCBIT;
  signal  \51324\    : AGCBIT;
  signal  \51325\    : AGCBIT;
  signal  \51326\    : AGCBIT; signal  \L04/\     : AGCBIT;
  signal \$51326\    : AGCBIT;
  signal  \51327\    : AGCBIT;
  signal  \51328\    : AGCBIT;
  signal  \51329\    : AGCBIT;
  signal  \51330\    : AGCBIT;
  signal \$51330\    : AGCBIT;
  signal  \51331\    : AGCBIT;
  signal  \51332\    : AGCBIT;
  signal \&51333\    : AGCBIT;
  signal  \51334\    : AGCBIT;
  signal  \51335\    : AGCBIT; signal  \Z04/\     : AGCBIT;
  signal \$51335\    : AGCBIT;
  signal  \51336\    : AGCBIT;
  signal  \51337\    : AGCBIT;
  signal  \51338\    : AGCBIT;
  signal  \51339\    : AGCBIT;
  signal \$51339\    : AGCBIT;
  signal  \51340\    : AGCBIT;
  signal  \51341\    : AGCBIT;
  signal  \51342\    : AGCBIT;
  signal  \51343\    : AGCBIT;
  signal  \51344\    : AGCBIT;
  signal  \51345\    : AGCBIT;
  signal  \51346\    : AGCBIT;
  signal \&51347\    : AGCBIT;
  signal  \51348\    : AGCBIT; signal  \G04/\     : AGCBIT;
  signal \$51348\    : AGCBIT;
  signal  \51349\    : AGCBIT; signal  \G04\      : AGCBIT;
  signal \&51350\    : AGCBIT;
  signal  \51351\    : AGCBIT;
  signal  \51352\    : AGCBIT; signal  \WL04\     : AGCBIT;
  signal \&51353\    : AGCBIT;
  signal  \51354\    : AGCBIT; signal  \WL04/\    : AGCBIT;
  signal  \51357\    : AGCBIT; signal  \RL04/\    : AGCBIT;
  signal \&51358\    : AGCBIT;
  signal  \51361\    : AGCBIT; signal  \CLEARC\   : AGCBIT;
  signal  \51362\    : AGCBIT; signal  \CLEARD\   : AGCBIT;
  signal \&51363\    : AGCBIT;
  signal  \51401\    : AGCBIT; signal  \CO06\     : AGCBIT;
  signal  \51402\    : AGCBIT;
  signal  \51403\    : AGCBIT;
  signal \$51403\    : AGCBIT;
  signal  \51404\    : AGCBIT;
  signal  \51405\    : AGCBIT;
  signal  \51406\    : AGCBIT;
  signal  \51407\    : AGCBIT;
  signal \$51407\    : AGCBIT;
  signal  \51408\    : AGCBIT;
  signal  \51409\    : AGCBIT;
  signal  \51410\    : AGCBIT; signal  \XUY03/\   : AGCBIT;
  signal  \51411\    : AGCBIT;
  signal  \51412\    : AGCBIT; signal  \SUMA03/\  : AGCBIT;
  signal  \51413\    : AGCBIT;
  signal  \51414\    : AGCBIT; signal  \CI04/\    : AGCBIT;
  signal  \51415\    : AGCBIT; signal  \SUMB03/\  : AGCBIT;
  signal  \51417\    : AGCBIT;
  signal  \51418\    : AGCBIT;
  signal  \51419\    : AGCBIT;
  signal  \51420\    : AGCBIT; signal  \A03/\     : AGCBIT;
  signal \$51420\    : AGCBIT;
  signal  \51421\    : AGCBIT;
  signal  \51422\    : AGCBIT;
  signal \&51423\    : AGCBIT;
  signal  \51424\    : AGCBIT;
  signal  \51425\    : AGCBIT;
  signal  \51426\    : AGCBIT; signal  \L03/\     : AGCBIT;
  signal \$51426\    : AGCBIT;
  signal  \51427\    : AGCBIT;
  signal  \51428\    : AGCBIT;
  signal  \51429\    : AGCBIT;
  signal  \51430\    : AGCBIT;
  signal \$51430\    : AGCBIT;
  signal  \51431\    : AGCBIT;
  signal  \51432\    : AGCBIT;
  signal \&51433\    : AGCBIT;
  signal  \51434\    : AGCBIT;
  signal  \51435\    : AGCBIT; signal  \Z03/\     : AGCBIT;
  signal \$51435\    : AGCBIT;
  signal  \51436\    : AGCBIT;
  signal  \51437\    : AGCBIT;
  signal  \51438\    : AGCBIT;
  signal  \51439\    : AGCBIT;
  signal \$51439\    : AGCBIT;
  signal  \51440\    : AGCBIT;
  signal  \51441\    : AGCBIT;
  signal  \51442\    : AGCBIT;
  signal  \51443\    : AGCBIT;
  signal  \51444\    : AGCBIT;
  signal  \51445\    : AGCBIT;
  signal  \51446\    : AGCBIT;
  signal \&51447\    : AGCBIT;
  signal  \51448\    : AGCBIT; signal  \G03/\     : AGCBIT;
  signal \$51448\    : AGCBIT;
  signal  \51449\    : AGCBIT; signal  \G03\      : AGCBIT;
  signal \&51450\    : AGCBIT;
  signal  \51451\    : AGCBIT;
  signal  \51452\    : AGCBIT; signal  \WL03\     : AGCBIT;
  signal \&51453\    : AGCBIT;
  signal  \51454\    : AGCBIT; signal  \WL03/\    : AGCBIT;
  signal  \51457\    : AGCBIT; signal  \RL03/\    : AGCBIT;
  signal \&51458\    : AGCBIT;
  signal  \51461\    : AGCBIT; signal  \CLEARB\   : AGCBIT;
  signal \&51462\    : AGCBIT;
  signal \&51463\    : AGCBIT;
  signal  \52101\    : AGCBIT; signal  \CO08\     : AGCBIT;
  signal  \52102\    : AGCBIT;
  signal  \52103\    : AGCBIT;
  signal \$52103\    : AGCBIT;
  signal  \52104\    : AGCBIT;
  signal  \52105\    : AGCBIT;
  signal  \52106\    : AGCBIT;
  signal  \52107\    : AGCBIT;
  signal \$52107\    : AGCBIT;
  signal  \52108\    : AGCBIT;
  signal  \52109\    : AGCBIT;
  signal  \52110\    : AGCBIT; signal  \XUY05/\   : AGCBIT;
  signal  \52111\    : AGCBIT;
  signal  \52112\    : AGCBIT; signal  \SUMA05/\  : AGCBIT;
  signal  \52113\    : AGCBIT;
  signal  \52114\    : AGCBIT; signal  \CI06/\    : AGCBIT;
  signal  \52115\    : AGCBIT; signal  \SUMB05/\  : AGCBIT;
  signal  \52117\    : AGCBIT;
  signal  \52118\    : AGCBIT;
  signal  \52119\    : AGCBIT;
  signal  \52120\    : AGCBIT; signal  \A05/\     : AGCBIT;
  signal \$52120\    : AGCBIT;
  signal  \52121\    : AGCBIT;
  signal  \52122\    : AGCBIT;
  signal \&52123\    : AGCBIT;
  signal  \52124\    : AGCBIT;
  signal  \52125\    : AGCBIT;
  signal  \52126\    : AGCBIT; signal  \L05/\     : AGCBIT;
  signal \$52126\    : AGCBIT;
  signal  \52127\    : AGCBIT;
  signal  \52128\    : AGCBIT;
  signal  \52129\    : AGCBIT;
  signal  \52130\    : AGCBIT;
  signal \$52130\    : AGCBIT;
  signal  \52131\    : AGCBIT;
  signal  \52132\    : AGCBIT;
  signal \&52133\    : AGCBIT;
  signal  \52134\    : AGCBIT;
  signal  \52135\    : AGCBIT; signal  \Z05/\     : AGCBIT;
  signal \$52135\    : AGCBIT;
  signal  \52136\    : AGCBIT;
  signal  \52137\    : AGCBIT;
  signal  \52138\    : AGCBIT;
  signal  \52139\    : AGCBIT;
  signal \$52139\    : AGCBIT;
  signal  \52140\    : AGCBIT;
  signal  \52141\    : AGCBIT;
  signal  \52142\    : AGCBIT;
  signal  \52143\    : AGCBIT;
  signal  \52144\    : AGCBIT;
  signal  \52145\    : AGCBIT;
  signal  \52146\    : AGCBIT;
  signal \&52147\    : AGCBIT;
  signal  \52148\    : AGCBIT; signal  \G05/\     : AGCBIT;
  signal \$52148\    : AGCBIT;
  signal  \52149\    : AGCBIT; signal  \G05\      : AGCBIT;
  signal \&52150\    : AGCBIT;
  signal  \52151\    : AGCBIT;
  signal  \52152\    : AGCBIT; signal  \WL05\     : AGCBIT;
  signal \&52153\    : AGCBIT;
  signal  \52154\    : AGCBIT; signal  \WL05/\    : AGCBIT;
  signal  \52157\    : AGCBIT; signal  \RL05/\    : AGCBIT;
  signal \&52158\    : AGCBIT;
  signal \&52162\    : AGCBIT;
  signal \&52163\    : AGCBIT;
  signal \&52201\    : AGCBIT;
  signal  \52202\    : AGCBIT;
  signal  \52203\    : AGCBIT;
  signal \$52203\    : AGCBIT;
  signal  \52204\    : AGCBIT;
  signal  \52205\    : AGCBIT;
  signal  \52206\    : AGCBIT;
  signal  \52207\    : AGCBIT;
  signal \$52207\    : AGCBIT;
  signal  \52208\    : AGCBIT;
  signal  \52209\    : AGCBIT;
  signal  \52210\    : AGCBIT; signal  \XUY06/\   : AGCBIT;
  signal  \52211\    : AGCBIT;
  signal  \52212\    : AGCBIT; signal  \SUMA06/\  : AGCBIT;
  signal  \52213\    : AGCBIT;
  signal  \52214\    : AGCBIT; signal  \CI07/\    : AGCBIT;
  signal  \52215\    : AGCBIT; signal  \SUMB06/\  : AGCBIT;
  signal  \52217\    : AGCBIT;
  signal  \52218\    : AGCBIT;
  signal  \52219\    : AGCBIT;
  signal  \52220\    : AGCBIT; signal  \A06/\     : AGCBIT;
  signal \$52220\    : AGCBIT;
  signal  \52221\    : AGCBIT;
  signal  \52222\    : AGCBIT;
  signal \&52223\    : AGCBIT;
  signal  \52224\    : AGCBIT;
  signal  \52225\    : AGCBIT;
  signal  \52226\    : AGCBIT; signal  \L06/\     : AGCBIT;
  signal \$52226\    : AGCBIT;
  signal  \52227\    : AGCBIT;
  signal  \52228\    : AGCBIT;
  signal  \52229\    : AGCBIT;
  signal  \52230\    : AGCBIT;
  signal \$52230\    : AGCBIT;
  signal  \52231\    : AGCBIT;
  signal  \52232\    : AGCBIT;
  signal \&52233\    : AGCBIT;
  signal  \52234\    : AGCBIT;
  signal  \52235\    : AGCBIT; signal  \Z06/\     : AGCBIT;
  signal \$52235\    : AGCBIT;
  signal  \52236\    : AGCBIT;
  signal  \52237\    : AGCBIT;
  signal  \52238\    : AGCBIT;
  signal  \52239\    : AGCBIT;
  signal \$52239\    : AGCBIT;
  signal  \52240\    : AGCBIT;
  signal  \52241\    : AGCBIT;
  signal  \52242\    : AGCBIT;
  signal  \52243\    : AGCBIT;
  signal  \52244\    : AGCBIT;
  signal  \52245\    : AGCBIT;
  signal  \52246\    : AGCBIT;
  signal \&52247\    : AGCBIT;
  signal  \52248\    : AGCBIT; signal  \G06/\     : AGCBIT;
  signal \$52248\    : AGCBIT;
  signal  \52249\    : AGCBIT; signal  \G06\      : AGCBIT;
  signal \&52250\    : AGCBIT;
  signal  \52251\    : AGCBIT;
  signal  \52252\    : AGCBIT; signal  \WL06\     : AGCBIT;
  signal \&52253\    : AGCBIT;
  signal  \52254\    : AGCBIT; signal  \WL06/\    : AGCBIT;
  signal  \52257\    : AGCBIT; signal  \RL06/\    : AGCBIT;
  signal \&52258\    : AGCBIT;
  signal  \52261\    : AGCBIT; signal  \PIPSAM/\  : AGCBIT;
  signal \&52301\    : AGCBIT;
  signal  \52302\    : AGCBIT;
  signal  \52303\    : AGCBIT;
  signal \$52303\    : AGCBIT;
  signal  \52304\    : AGCBIT;
  signal  \52305\    : AGCBIT;
  signal  \52306\    : AGCBIT;
  signal  \52307\    : AGCBIT;
  signal \$52307\    : AGCBIT;
  signal  \52308\    : AGCBIT;
  signal  \52309\    : AGCBIT;
  signal  \52310\    : AGCBIT; signal  \XUY08/\   : AGCBIT;
  signal  \52311\    : AGCBIT;
  signal  \52312\    : AGCBIT; signal  \SUMA08/\  : AGCBIT;
  signal  \52313\    : AGCBIT;
  signal  \52314\    : AGCBIT; signal  \CI09/\    : AGCBIT;
  signal  \52315\    : AGCBIT; signal  \SUMB08/\  : AGCBIT;
  signal  \52317\    : AGCBIT;
  signal  \52318\    : AGCBIT;
  signal  \52319\    : AGCBIT;
  signal  \52320\    : AGCBIT; signal  \A08/\     : AGCBIT;
  signal \$52320\    : AGCBIT;
  signal  \52321\    : AGCBIT;
  signal  \52322\    : AGCBIT;
  signal \&52323\    : AGCBIT;
  signal  \52324\    : AGCBIT;
  signal  \52325\    : AGCBIT;
  signal  \52326\    : AGCBIT; signal  \L08/\     : AGCBIT;
  signal \$52326\    : AGCBIT;
  signal  \52327\    : AGCBIT;
  signal  \52328\    : AGCBIT;
  signal  \52329\    : AGCBIT;
  signal  \52330\    : AGCBIT;
  signal \$52330\    : AGCBIT;
  signal  \52331\    : AGCBIT;
  signal  \52332\    : AGCBIT;
  signal \&52333\    : AGCBIT;
  signal  \52334\    : AGCBIT;
  signal  \52335\    : AGCBIT; signal  \Z08/\     : AGCBIT;
  signal \$52335\    : AGCBIT;
  signal  \52336\    : AGCBIT;
  signal  \52337\    : AGCBIT;
  signal  \52338\    : AGCBIT;
  signal  \52339\    : AGCBIT;
  signal \$52339\    : AGCBIT;
  signal  \52340\    : AGCBIT;
  signal  \52341\    : AGCBIT;
  signal  \52342\    : AGCBIT;
  signal  \52343\    : AGCBIT;
  signal  \52344\    : AGCBIT;
  signal  \52345\    : AGCBIT;
  signal  \52346\    : AGCBIT;
  signal \&52347\    : AGCBIT;
  signal  \52348\    : AGCBIT; signal  \G08/\     : AGCBIT;
  signal \$52348\    : AGCBIT;
  signal  \52349\    : AGCBIT; signal  \G08\      : AGCBIT;
  signal \&52350\    : AGCBIT;
  signal  \52351\    : AGCBIT;
  signal  \52352\    : AGCBIT; signal  \WL08\     : AGCBIT;
  signal \&52353\    : AGCBIT;
  signal  \52354\    : AGCBIT; signal  \WL08/\    : AGCBIT;
  signal  \52357\    : AGCBIT; signal  \RL08/\    : AGCBIT;
  signal \&52358\    : AGCBIT;
  signal  \52361\    : AGCBIT; signal  \PIPGX-\   : AGCBIT;
  signal  \52362\    : AGCBIT; signal  \PIPGY+\   : AGCBIT;
  signal \&52363\    : AGCBIT;
  signal  \52401\    : AGCBIT; signal  \CO10\     : AGCBIT;
  signal  \52402\    : AGCBIT;
  signal  \52403\    : AGCBIT;
  signal \$52403\    : AGCBIT;
  signal  \52404\    : AGCBIT;
  signal  \52405\    : AGCBIT;
  signal  \52406\    : AGCBIT;
  signal  \52407\    : AGCBIT;
  signal \$52407\    : AGCBIT;
  signal  \52408\    : AGCBIT;
  signal  \52409\    : AGCBIT;
  signal  \52410\    : AGCBIT; signal  \XUY07/\   : AGCBIT;
  signal  \52411\    : AGCBIT;
  signal  \52412\    : AGCBIT; signal  \SUMA07/\  : AGCBIT;
  signal  \52413\    : AGCBIT;
  signal  \52414\    : AGCBIT; signal  \CI08/\    : AGCBIT;
  signal  \52415\    : AGCBIT; signal  \SUMB07/\  : AGCBIT;
  signal  \52417\    : AGCBIT;
  signal  \52418\    : AGCBIT;
  signal  \52419\    : AGCBIT;
  signal  \52420\    : AGCBIT; signal  \A07/\     : AGCBIT;
  signal \$52420\    : AGCBIT;
  signal  \52421\    : AGCBIT;
  signal  \52422\    : AGCBIT;
  signal \&52423\    : AGCBIT;
  signal  \52424\    : AGCBIT;
  signal  \52425\    : AGCBIT;
  signal  \52426\    : AGCBIT; signal  \L07/\     : AGCBIT;
  signal \$52426\    : AGCBIT;
  signal  \52427\    : AGCBIT;
  signal  \52428\    : AGCBIT;
  signal  \52429\    : AGCBIT;
  signal  \52430\    : AGCBIT;
  signal \$52430\    : AGCBIT;
  signal  \52431\    : AGCBIT;
  signal  \52432\    : AGCBIT;
  signal \&52433\    : AGCBIT;
  signal  \52434\    : AGCBIT;
  signal  \52435\    : AGCBIT; signal  \Z07/\     : AGCBIT;
  signal \$52435\    : AGCBIT;
  signal  \52436\    : AGCBIT;
  signal  \52437\    : AGCBIT;
  signal  \52438\    : AGCBIT;
  signal  \52439\    : AGCBIT;
  signal \$52439\    : AGCBIT;
  signal  \52440\    : AGCBIT;
  signal  \52441\    : AGCBIT;
  signal  \52442\    : AGCBIT;
  signal  \52443\    : AGCBIT;
  signal  \52444\    : AGCBIT;
  signal  \52445\    : AGCBIT;
  signal  \52446\    : AGCBIT;
  signal \&52447\    : AGCBIT;
  signal  \52448\    : AGCBIT; signal  \G07/\     : AGCBIT;
  signal \$52448\    : AGCBIT;
  signal  \52449\    : AGCBIT; signal  \G07\      : AGCBIT;
  signal \&52450\    : AGCBIT;
  signal  \52451\    : AGCBIT;
  signal  \52452\    : AGCBIT; signal  \WL07\     : AGCBIT;
  signal \&52453\    : AGCBIT;
  signal  \52454\    : AGCBIT; signal  \WL07/\    : AGCBIT;
  signal  \52457\    : AGCBIT; signal  \RL07/\    : AGCBIT;
  signal \&52458\    : AGCBIT;
  signal  \52461\    : AGCBIT; signal  \PIPGX+\   : AGCBIT;
  signal \&52462\    : AGCBIT;
  signal \&52463\    : AGCBIT;
  signal  \53101\    : AGCBIT; signal  \CO12\     : AGCBIT;
  signal  \53102\    : AGCBIT;
  signal  \53103\    : AGCBIT;
  signal \$53103\    : AGCBIT;
  signal  \53104\    : AGCBIT;
  signal  \53105\    : AGCBIT;
  signal  \53106\    : AGCBIT;
  signal  \53107\    : AGCBIT;
  signal \$53107\    : AGCBIT;
  signal  \53108\    : AGCBIT;
  signal  \53109\    : AGCBIT;
  signal  \53110\    : AGCBIT; signal  \XUY09/\   : AGCBIT;
  signal  \53111\    : AGCBIT;
  signal  \53112\    : AGCBIT; signal  \SUMA09/\  : AGCBIT;
  signal  \53113\    : AGCBIT;
  signal  \53114\    : AGCBIT; signal  \CI10/\    : AGCBIT;
  signal  \53115\    : AGCBIT; signal  \SUMB09/\  : AGCBIT;
  signal  \53117\    : AGCBIT;
  signal  \53118\    : AGCBIT;
  signal  \53119\    : AGCBIT;
  signal  \53120\    : AGCBIT; signal  \A09/\     : AGCBIT;
  signal \$53120\    : AGCBIT;
  signal  \53121\    : AGCBIT;
  signal  \53122\    : AGCBIT;
  signal \&53123\    : AGCBIT;
  signal  \53124\    : AGCBIT;
  signal  \53125\    : AGCBIT;
  signal  \53126\    : AGCBIT; signal  \L09/\     : AGCBIT;
  signal \$53126\    : AGCBIT;
  signal  \53127\    : AGCBIT;
  signal  \53128\    : AGCBIT;
  signal  \53129\    : AGCBIT;
  signal  \53130\    : AGCBIT;
  signal \$53130\    : AGCBIT;
  signal  \53131\    : AGCBIT;
  signal  \53132\    : AGCBIT;
  signal \&53133\    : AGCBIT;
  signal  \53134\    : AGCBIT;
  signal  \53135\    : AGCBIT; signal  \Z09/\     : AGCBIT;
  signal \$53135\    : AGCBIT;
  signal  \53136\    : AGCBIT;
  signal  \53137\    : AGCBIT;
  signal  \53138\    : AGCBIT;
  signal  \53139\    : AGCBIT;
  signal \$53139\    : AGCBIT;
  signal  \53140\    : AGCBIT;
  signal  \53141\    : AGCBIT;
  signal  \53142\    : AGCBIT;
  signal  \53143\    : AGCBIT;
  signal  \53144\    : AGCBIT;
  signal  \53145\    : AGCBIT;
  signal  \53146\    : AGCBIT;
  signal \&53147\    : AGCBIT;
  signal  \53148\    : AGCBIT; signal  \G09/\     : AGCBIT;
  signal \$53148\    : AGCBIT;
  signal  \53149\    : AGCBIT; signal  \G09\      : AGCBIT;
  signal \&53150\    : AGCBIT;
  signal  \53151\    : AGCBIT;
  signal  \53152\    : AGCBIT; signal  \WL09\     : AGCBIT;
  signal \&53153\    : AGCBIT;
  signal  \53154\    : AGCBIT; signal  \WL09/\    : AGCBIT;
  signal  \53157\    : AGCBIT; signal  \RL09/\    : AGCBIT;
  signal \&53158\    : AGCBIT;
  signal  \53161\    : AGCBIT; signal  \PIPGY-\   : AGCBIT;
  signal \&53201\    : AGCBIT;
  signal  \53202\    : AGCBIT;
  signal  \53203\    : AGCBIT;
  signal \$53203\    : AGCBIT;
  signal  \53204\    : AGCBIT;
  signal  \53205\    : AGCBIT;
  signal  \53206\    : AGCBIT;
  signal  \53207\    : AGCBIT;
  signal \$53207\    : AGCBIT;
  signal  \53208\    : AGCBIT;
  signal  \53209\    : AGCBIT;
  signal  \53210\    : AGCBIT; signal  \XUY10/\   : AGCBIT;
  signal  \53211\    : AGCBIT;
  signal  \53212\    : AGCBIT; signal  \SUMA10/\  : AGCBIT;
  signal  \53213\    : AGCBIT;
  signal  \53214\    : AGCBIT; signal  \CI11/\    : AGCBIT;
  signal  \53215\    : AGCBIT; signal  \SUMB10/\  : AGCBIT;
  signal  \53217\    : AGCBIT;
  signal  \53218\    : AGCBIT;
  signal  \53219\    : AGCBIT;
  signal  \53220\    : AGCBIT; signal  \A10/\     : AGCBIT;
  signal \$53220\    : AGCBIT;
  signal  \53221\    : AGCBIT;
  signal  \53222\    : AGCBIT;
  signal \&53223\    : AGCBIT;
  signal  \53224\    : AGCBIT;
  signal  \53225\    : AGCBIT;
  signal  \53226\    : AGCBIT; signal  \L10/\     : AGCBIT;
  signal \$53226\    : AGCBIT;
  signal  \53227\    : AGCBIT;
  signal  \53228\    : AGCBIT;
  signal  \53229\    : AGCBIT;
  signal  \53230\    : AGCBIT;
  signal \$53230\    : AGCBIT;
  signal  \53231\    : AGCBIT;
  signal  \53232\    : AGCBIT;
  signal \&53233\    : AGCBIT;
  signal  \53234\    : AGCBIT;
  signal  \53235\    : AGCBIT; signal  \Z10/\     : AGCBIT;
  signal \$53235\    : AGCBIT;
  signal  \53236\    : AGCBIT;
  signal  \53237\    : AGCBIT;
  signal  \53238\    : AGCBIT;
  signal  \53239\    : AGCBIT;
  signal \$53239\    : AGCBIT;
  signal  \53240\    : AGCBIT;
  signal  \53241\    : AGCBIT;
  signal  \53242\    : AGCBIT;
  signal  \53243\    : AGCBIT;
  signal  \53244\    : AGCBIT;
  signal  \53245\    : AGCBIT;
  signal  \53246\    : AGCBIT;
  signal \&53247\    : AGCBIT;
  signal  \53248\    : AGCBIT; signal  \G10/\     : AGCBIT;
  signal \$53248\    : AGCBIT;
  signal  \53249\    : AGCBIT; signal  \G10\      : AGCBIT;
  signal \&53250\    : AGCBIT;
  signal  \53251\    : AGCBIT;
  signal  \53252\    : AGCBIT; signal  \WL10\     : AGCBIT;
  signal \&53253\    : AGCBIT;
  signal  \53254\    : AGCBIT; signal  \WL10/\    : AGCBIT;
  signal  \53257\    : AGCBIT; signal  \RL10/\    : AGCBIT;
  signal \&53258\    : AGCBIT;
  signal  \53261\    : AGCBIT; signal  \PIPGZ+\   : AGCBIT;
  signal  \53262\    : AGCBIT; signal  \PIPGZ-\   : AGCBIT;
  signal \&53301\    : AGCBIT;
  signal  \53302\    : AGCBIT;
  signal  \53303\    : AGCBIT;
  signal \$53303\    : AGCBIT;
  signal  \53304\    : AGCBIT;
  signal  \53305\    : AGCBIT;
  signal  \53306\    : AGCBIT;
  signal  \53307\    : AGCBIT;
  signal \$53307\    : AGCBIT;
  signal  \53308\    : AGCBIT;
  signal  \53309\    : AGCBIT;
  signal  \53310\    : AGCBIT; signal  \XUY12/\   : AGCBIT;
  signal  \53311\    : AGCBIT;
  signal  \53312\    : AGCBIT; signal  \SUMA12/\  : AGCBIT;
  signal  \53313\    : AGCBIT;
  signal  \53314\    : AGCBIT; signal  \CI13/\    : AGCBIT;
  signal  \53315\    : AGCBIT; signal  \SUMB12/\  : AGCBIT;
  signal  \53317\    : AGCBIT;
  signal  \53318\    : AGCBIT;
  signal  \53319\    : AGCBIT;
  signal  \53320\    : AGCBIT; signal  \A12/\     : AGCBIT;
  signal \$53320\    : AGCBIT;
  signal  \53321\    : AGCBIT;
  signal  \53322\    : AGCBIT;
  signal \&53323\    : AGCBIT;
  signal  \53324\    : AGCBIT;
  signal  \53325\    : AGCBIT;
  signal  \53326\    : AGCBIT; signal  \L12/\     : AGCBIT;
  signal \$53326\    : AGCBIT;
  signal  \53327\    : AGCBIT;
  signal  \53328\    : AGCBIT;
  signal  \53329\    : AGCBIT;
  signal  \53330\    : AGCBIT;
  signal \$53330\    : AGCBIT;
  signal  \53331\    : AGCBIT;
  signal  \53332\    : AGCBIT;
  signal \&53333\    : AGCBIT;
  signal  \53334\    : AGCBIT;
  signal  \53335\    : AGCBIT; signal  \Z12/\     : AGCBIT;
  signal \$53335\    : AGCBIT;
  signal  \53336\    : AGCBIT;
  signal  \53337\    : AGCBIT;
  signal  \53338\    : AGCBIT;
  signal  \53339\    : AGCBIT;
  signal \$53339\    : AGCBIT;
  signal  \53340\    : AGCBIT;
  signal  \53341\    : AGCBIT;
  signal  \53342\    : AGCBIT;
  signal  \53343\    : AGCBIT;
  signal  \53344\    : AGCBIT;
  signal  \53345\    : AGCBIT;
  signal  \53346\    : AGCBIT;
  signal \&53347\    : AGCBIT;
  signal  \53348\    : AGCBIT; signal  \G12/\     : AGCBIT;
  signal \$53348\    : AGCBIT;
  signal  \53349\    : AGCBIT; signal  \G12\      : AGCBIT;
  signal \&53350\    : AGCBIT;
  signal  \53351\    : AGCBIT;
  signal  \53352\    : AGCBIT; signal  \WL12\     : AGCBIT;
  signal \&53353\    : AGCBIT;
  signal  \53354\    : AGCBIT; signal  \WL12/\    : AGCBIT;
  signal  \53357\    : AGCBIT; signal  \RL12/\    : AGCBIT;
  signal \&53358\    : AGCBIT;
  signal  \53361\    : AGCBIT; signal  \PIPAX-/\  : AGCBIT;
  signal  \53362\    : AGCBIT; signal  \PIPAY+/\  : AGCBIT;
  signal \&53363\    : AGCBIT;
  signal  \53401\    : AGCBIT; signal  \CO14\     : AGCBIT;
  signal  \53402\    : AGCBIT;
  signal  \53403\    : AGCBIT;
  signal \$53403\    : AGCBIT;
  signal  \53404\    : AGCBIT;
  signal  \53405\    : AGCBIT;
  signal  \53406\    : AGCBIT;
  signal  \53407\    : AGCBIT;
  signal \$53407\    : AGCBIT;
  signal  \53408\    : AGCBIT;
  signal  \53409\    : AGCBIT;
  signal  \53410\    : AGCBIT; signal  \XUY11/\   : AGCBIT;
  signal  \53411\    : AGCBIT;
  signal  \53412\    : AGCBIT; signal  \SUMA11/\  : AGCBIT;
  signal  \53413\    : AGCBIT;
  signal  \53414\    : AGCBIT; signal  \CI12/\    : AGCBIT;
  signal  \53415\    : AGCBIT; signal  \SUMB11/\  : AGCBIT;
  signal  \53417\    : AGCBIT;
  signal  \53418\    : AGCBIT;
  signal  \53419\    : AGCBIT;
  signal  \53420\    : AGCBIT; signal  \A11/\     : AGCBIT;
  signal \$53420\    : AGCBIT;
  signal  \53421\    : AGCBIT;
  signal  \53422\    : AGCBIT;
  signal \&53423\    : AGCBIT;
  signal  \53424\    : AGCBIT;
  signal  \53425\    : AGCBIT;
  signal  \53426\    : AGCBIT; signal  \L11/\     : AGCBIT;
  signal \$53426\    : AGCBIT;
  signal  \53427\    : AGCBIT;
  signal  \53428\    : AGCBIT;
  signal  \53429\    : AGCBIT;
  signal  \53430\    : AGCBIT;
  signal \$53430\    : AGCBIT;
  signal  \53431\    : AGCBIT;
  signal  \53432\    : AGCBIT;
  signal \&53433\    : AGCBIT;
  signal  \53434\    : AGCBIT;
  signal  \53435\    : AGCBIT; signal  \Z11/\     : AGCBIT;
  signal \$53435\    : AGCBIT;
  signal  \53436\    : AGCBIT;
  signal  \53437\    : AGCBIT;
  signal  \53438\    : AGCBIT;
  signal  \53439\    : AGCBIT;
  signal \$53439\    : AGCBIT;
  signal  \53440\    : AGCBIT;
  signal  \53441\    : AGCBIT;
  signal  \53442\    : AGCBIT;
  signal  \53443\    : AGCBIT;
  signal  \53444\    : AGCBIT;
  signal  \53445\    : AGCBIT;
  signal  \53446\    : AGCBIT;
  signal \&53447\    : AGCBIT;
  signal  \53448\    : AGCBIT; signal  \G11/\     : AGCBIT;
  signal \$53448\    : AGCBIT;
  signal  \53449\    : AGCBIT; signal  \G11\      : AGCBIT;
  signal \&53450\    : AGCBIT;
  signal  \53451\    : AGCBIT;
  signal  \53452\    : AGCBIT; signal  \WL11\     : AGCBIT;
  signal \&53453\    : AGCBIT;
  signal  \53454\    : AGCBIT; signal  \WL11/\    : AGCBIT;
  signal  \53457\    : AGCBIT; signal  \RL11/\    : AGCBIT;
  signal \&53458\    : AGCBIT;
  signal  \53461\    : AGCBIT; signal  \PIPAX+/\  : AGCBIT;
  signal \&53462\    : AGCBIT;
  signal \&53463\    : AGCBIT;
  signal  \54101\    : AGCBIT; signal  \CO16\     : AGCBIT;
  signal  \54102\    : AGCBIT;
  signal  \54103\    : AGCBIT;
  signal \$54103\    : AGCBIT;
  signal  \54104\    : AGCBIT;
  signal  \54105\    : AGCBIT;
  signal  \54106\    : AGCBIT;
  signal  \54107\    : AGCBIT;
  signal \$54107\    : AGCBIT;
  signal  \54108\    : AGCBIT;
  signal  \54109\    : AGCBIT;
  signal  \54110\    : AGCBIT; signal  \XUY13/\   : AGCBIT;
  signal  \54111\    : AGCBIT;
  signal  \54112\    : AGCBIT; signal  \SUMA13/\  : AGCBIT;
  signal  \54113\    : AGCBIT;
  signal  \54114\    : AGCBIT; signal  \CI14/\    : AGCBIT;
  signal  \54115\    : AGCBIT; signal  \SUMB13/\  : AGCBIT;
  signal  \54117\    : AGCBIT;
  signal  \54118\    : AGCBIT;
  signal  \54119\    : AGCBIT;
  signal  \54120\    : AGCBIT; signal  \A13/\     : AGCBIT;
  signal \$54120\    : AGCBIT;
  signal  \54121\    : AGCBIT;
  signal  \54122\    : AGCBIT;
  signal \&54123\    : AGCBIT;
  signal  \54124\    : AGCBIT;
  signal  \54125\    : AGCBIT;
  signal  \54126\    : AGCBIT; signal  \L13/\     : AGCBIT;
  signal \$54126\    : AGCBIT;
  signal  \54127\    : AGCBIT;
  signal  \54128\    : AGCBIT;
  signal  \54129\    : AGCBIT;
  signal  \54130\    : AGCBIT;
  signal \$54130\    : AGCBIT;
  signal  \54131\    : AGCBIT;
  signal  \54132\    : AGCBIT;
  signal \&54133\    : AGCBIT;
  signal  \54134\    : AGCBIT;
  signal  \54135\    : AGCBIT; signal  \Z13/\     : AGCBIT;
  signal \$54135\    : AGCBIT;
  signal  \54136\    : AGCBIT;
  signal  \54137\    : AGCBIT;
  signal  \54138\    : AGCBIT;
  signal  \54139\    : AGCBIT;
  signal \$54139\    : AGCBIT;
  signal  \54140\    : AGCBIT;
  signal  \54141\    : AGCBIT;
  signal  \54142\    : AGCBIT;
  signal  \54143\    : AGCBIT;
  signal  \54144\    : AGCBIT;
  signal  \54145\    : AGCBIT;
  signal  \54146\    : AGCBIT;
  signal \&54147\    : AGCBIT;
  signal  \54148\    : AGCBIT; signal  \G13/\     : AGCBIT;
  signal \$54148\    : AGCBIT;
  signal  \54149\    : AGCBIT; signal  \G13\      : AGCBIT;
  signal \&54150\    : AGCBIT;
  signal  \54151\    : AGCBIT;
  signal  \54152\    : AGCBIT; signal  \WL13\     : AGCBIT;
  signal \&54153\    : AGCBIT;
  signal  \54154\    : AGCBIT; signal  \WL13/\    : AGCBIT;
  signal  \54157\    : AGCBIT; signal  \RL13/\    : AGCBIT;
  signal \&54158\    : AGCBIT;
  signal  \54161\    : AGCBIT; signal  \WHOMP/\   : AGCBIT;
  signal \$54161\    : AGCBIT;
  signal \&54162\    : AGCBIT;
  signal \&54163\    : AGCBIT;
  signal \&54201\    : AGCBIT;
  signal  \54202\    : AGCBIT;
  signal  \54203\    : AGCBIT;
  signal \$54203\    : AGCBIT;
  signal  \54204\    : AGCBIT;
  signal  \54205\    : AGCBIT;
  signal  \54206\    : AGCBIT;
  signal  \54207\    : AGCBIT;
  signal \$54207\    : AGCBIT;
  signal  \54208\    : AGCBIT;
  signal  \54209\    : AGCBIT;
  signal  \54210\    : AGCBIT; signal  \XUY14/\   : AGCBIT;
  signal  \54211\    : AGCBIT;
  signal  \54212\    : AGCBIT; signal  \SUMA14/\  : AGCBIT;
  signal  \54213\    : AGCBIT;
  signal  \54214\    : AGCBIT; signal  \CI15/\    : AGCBIT;
  signal  \54215\    : AGCBIT; signal  \SUMB14/\  : AGCBIT;
  signal  \54217\    : AGCBIT;
  signal  \54218\    : AGCBIT;
  signal  \54219\    : AGCBIT;
  signal  \54220\    : AGCBIT; signal  \A14/\     : AGCBIT;
  signal \$54220\    : AGCBIT;
  signal  \54221\    : AGCBIT;
  signal  \54222\    : AGCBIT;
  signal \&54223\    : AGCBIT;
  signal  \54224\    : AGCBIT;
  signal  \54225\    : AGCBIT;
  signal  \54226\    : AGCBIT; signal  \L14/\     : AGCBIT;
  signal \$54226\    : AGCBIT;
  signal  \54227\    : AGCBIT;
  signal  \54228\    : AGCBIT;
  signal  \54229\    : AGCBIT;
  signal  \54230\    : AGCBIT;
  signal \$54230\    : AGCBIT;
  signal  \54231\    : AGCBIT;
  signal  \54232\    : AGCBIT;
  signal \&54233\    : AGCBIT;
  signal  \54234\    : AGCBIT;
  signal  \54235\    : AGCBIT; signal  \Z14/\     : AGCBIT;
  signal \$54235\    : AGCBIT;
  signal  \54236\    : AGCBIT;
  signal  \54237\    : AGCBIT;
  signal  \54238\    : AGCBIT;
  signal  \54239\    : AGCBIT;
  signal \$54239\    : AGCBIT;
  signal  \54240\    : AGCBIT;
  signal  \54241\    : AGCBIT;
  signal  \54242\    : AGCBIT;
  signal  \54243\    : AGCBIT;
  signal  \54244\    : AGCBIT;
  signal  \54245\    : AGCBIT;
  signal  \54246\    : AGCBIT;
  signal \&54247\    : AGCBIT;
  signal  \54248\    : AGCBIT; signal  \G14/\     : AGCBIT;
  signal \$54248\    : AGCBIT;
  signal  \54249\    : AGCBIT; signal  \G14\      : AGCBIT;
  signal \&54250\    : AGCBIT;
  signal  \54251\    : AGCBIT;
  signal  \54252\    : AGCBIT; signal  \WL14\     : AGCBIT;
  signal \&54253\    : AGCBIT;
  signal  \54254\    : AGCBIT; signal  \WL14/\    : AGCBIT;
  signal  \54257\    : AGCBIT; signal  \RL14/\    : AGCBIT;
  signal \&54258\    : AGCBIT;
  signal  \54261\    : AGCBIT; signal  \GTRST/\   : AGCBIT;
  signal  \54262\    : AGCBIT; signal  \WHOMP\    : AGCBIT;
  signal \$54262\    : AGCBIT;
  signal \&54263\    : AGCBIT;
  signal \&54301\    : AGCBIT;
  signal  \54302\    : AGCBIT;
  signal  \54303\    : AGCBIT;
  signal \$54303\    : AGCBIT;
  signal  \54304\    : AGCBIT;
  signal  \54305\    : AGCBIT;
  signal  \54306\    : AGCBIT;
  signal  \54307\    : AGCBIT;
  signal \$54307\    : AGCBIT;
  signal  \54308\    : AGCBIT;
  signal  \54309\    : AGCBIT;
  signal  \54310\    : AGCBIT; signal  \XUY16/\   : AGCBIT;
  signal  \54311\    : AGCBIT;
  signal  \54312\    : AGCBIT; signal  \SUMA16/\  : AGCBIT;
  signal  \54313\    : AGCBIT;
  signal  \54314\    : AGCBIT; signal  \EAC/\     : AGCBIT;
  signal  \54315\    : AGCBIT; signal  \SUMB16/\  : AGCBIT;
  signal  \54317\    : AGCBIT;
  signal  \54318\    : AGCBIT;
  signal  \54319\    : AGCBIT;
  signal  \54320\    : AGCBIT; signal  \A16/\     : AGCBIT;
  signal \$54320\    : AGCBIT;
  signal  \54321\    : AGCBIT;
  signal  \54322\    : AGCBIT;
  signal \&54323\    : AGCBIT;
  signal  \54324\    : AGCBIT;
  signal  \54325\    : AGCBIT;
  signal  \54326\    : AGCBIT; signal  \L16/\     : AGCBIT;
  signal \$54326\    : AGCBIT;
  signal  \54327\    : AGCBIT;
  signal  \54328\    : AGCBIT; signal  \RL16\     : AGCBIT;
  signal  \54329\    : AGCBIT;
  signal  \54330\    : AGCBIT;
  signal \$54330\    : AGCBIT;
  signal  \54331\    : AGCBIT;
  signal  \54332\    : AGCBIT;
  signal \&54333\    : AGCBIT;
  signal  \54334\    : AGCBIT;
  signal  \54335\    : AGCBIT; signal  \Z16/\     : AGCBIT;
  signal \$54335\    : AGCBIT;
  signal  \54336\    : AGCBIT;
  signal  \54337\    : AGCBIT;
  signal  \54338\    : AGCBIT;
  signal  \54339\    : AGCBIT;
  signal \$54339\    : AGCBIT;
  signal  \54340\    : AGCBIT;
  signal  \54341\    : AGCBIT;
  signal  \54342\    : AGCBIT;
  signal  \54343\    : AGCBIT;
  signal  \54344\    : AGCBIT;
  signal  \54345\    : AGCBIT;
  signal  \54346\    : AGCBIT;
  signal \&54347\    : AGCBIT;
  signal  \54348\    : AGCBIT; signal  \G16/\     : AGCBIT;
  signal \$54348\    : AGCBIT;
  signal  \54349\    : AGCBIT; signal  \G16\      : AGCBIT;
  signal \&54350\    : AGCBIT;
  signal  \54351\    : AGCBIT;
  signal  \54352\    : AGCBIT; signal  \WL16\     : AGCBIT;
  signal \&54353\    : AGCBIT;
  signal  \54354\    : AGCBIT; signal  \WL16/\    : AGCBIT;
  signal  \54357\    : AGCBIT; signal  \RL16/\    : AGCBIT;
  signal \&54358\    : AGCBIT;
  signal  \54361\    : AGCBIT; signal  \PIPAZ+/\  : AGCBIT;
  signal  \54362\    : AGCBIT; signal  \PIPAZ-/\  : AGCBIT;
  signal \&54363\    : AGCBIT;
  signal  \54401\    : AGCBIT; signal  \CO02\     : AGCBIT;
  signal  \54402\    : AGCBIT;
  signal  \54403\    : AGCBIT;
  signal \$54403\    : AGCBIT;
  signal  \54404\    : AGCBIT;
  signal  \54405\    : AGCBIT;
  signal  \54406\    : AGCBIT;
  signal  \54407\    : AGCBIT;
  signal \$54407\    : AGCBIT;
  signal  \54408\    : AGCBIT;
  signal  \54409\    : AGCBIT;
  signal  \54410\    : AGCBIT; signal  \XUY15/\   : AGCBIT;
  signal  \54411\    : AGCBIT;
  signal  \54412\    : AGCBIT; signal  \SUMA15/\  : AGCBIT;
  signal  \54413\    : AGCBIT;
  signal  \54414\    : AGCBIT; signal  \CI16/\    : AGCBIT;
  signal  \54415\    : AGCBIT; signal  \SUMB15/\  : AGCBIT;
  signal  \54417\    : AGCBIT;
  signal  \54418\    : AGCBIT;
  signal  \54419\    : AGCBIT;
  signal  \54420\    : AGCBIT; signal  \A15/\     : AGCBIT;
  signal \$54420\    : AGCBIT;
  signal  \54421\    : AGCBIT;
  signal  \54422\    : AGCBIT;
  signal \&54423\    : AGCBIT;
  signal  \54424\    : AGCBIT;
  signal  \54425\    : AGCBIT;
  signal  \54426\    : AGCBIT; signal  \L15/\     : AGCBIT;
  signal \$54426\    : AGCBIT;
  signal  \54427\    : AGCBIT;
  signal  \54429\    : AGCBIT;
  signal  \54430\    : AGCBIT;
  signal \$54430\    : AGCBIT;
  signal  \54431\    : AGCBIT;
  signal  \54432\    : AGCBIT;
  signal \&54433\    : AGCBIT;
  signal  \54434\    : AGCBIT;
  signal  \54435\    : AGCBIT; signal  \Z15/\     : AGCBIT;
  signal \$54435\    : AGCBIT;
  signal  \54436\    : AGCBIT;
  signal  \54437\    : AGCBIT;
  signal  \54438\    : AGCBIT;
  signal  \54439\    : AGCBIT;
  signal \$54439\    : AGCBIT;
  signal  \54440\    : AGCBIT;
  signal  \54441\    : AGCBIT;
  signal  \54442\    : AGCBIT;
  signal  \54443\    : AGCBIT;
  signal  \54444\    : AGCBIT;
  signal  \54445\    : AGCBIT;
  signal  \54446\    : AGCBIT;
  signal \&54447\    : AGCBIT;
  signal  \54448\    : AGCBIT; signal  \G15/\     : AGCBIT;
  signal \$54448\    : AGCBIT;
  signal  \54449\    : AGCBIT; signal  \G15\      : AGCBIT;
  signal  \54451\    : AGCBIT;
  signal  \54452\    : AGCBIT; signal  \WL15\     : AGCBIT;
  signal \&54453\    : AGCBIT;
  signal  \54454\    : AGCBIT; signal  \WL15/\    : AGCBIT;
  signal  \54457\    : AGCBIT; signal  \RL15/\    : AGCBIT;
  signal \&54458\    : AGCBIT;
  signal  \54461\    : AGCBIT; signal  \PIPAY-/\  : AGCBIT;
  signal \&54462\    : AGCBIT;
  signal \&54463\    : AGCBIT;
  signal  \34101\    : AGCBIT; signal  \G01A/\    : AGCBIT;
  signal  \34102\    : AGCBIT;
  signal  \34103\    : AGCBIT;
  signal  \34104\    : AGCBIT;
  signal  \34105\    : AGCBIT;
  signal  \34106\    : AGCBIT;
  signal  \34107\    : AGCBIT;
  signal  \34108\    : AGCBIT; signal  \PA03\     : AGCBIT;
  signal \&34109\    : AGCBIT;
  signal  \34110\    : AGCBIT; signal  \PA03/\    : AGCBIT;
  signal  \34111\    : AGCBIT;
  signal  \34112\    : AGCBIT;
  signal  \34113\    : AGCBIT;
  signal  \34114\    : AGCBIT;
  signal  \34115\    : AGCBIT;
  signal  \34116\    : AGCBIT;
  signal  \34117\    : AGCBIT;
  signal  \34118\    : AGCBIT; signal  \PA06\     : AGCBIT;
  signal \&34119\    : AGCBIT;
  signal  \34120\    : AGCBIT; signal  \PA06/\    : AGCBIT;
  signal  \34121\    : AGCBIT;
  signal  \34122\    : AGCBIT;
  signal  \34123\    : AGCBIT;
  signal  \34124\    : AGCBIT;
  signal  \34125\    : AGCBIT;
  signal  \34126\    : AGCBIT;
  signal  \34127\    : AGCBIT;
  signal  \34128\    : AGCBIT;
  signal  \34129\    : AGCBIT; signal  \PA09\     : AGCBIT;
  signal \&34130\    : AGCBIT;
  signal  \34131\    : AGCBIT; signal  \PA09/\    : AGCBIT;
  signal  \34132\    : AGCBIT;
  signal  \34133\    : AGCBIT;
  signal  \34134\    : AGCBIT;
  signal  \34135\    : AGCBIT;
  signal  \34136\    : AGCBIT;
  signal  \34137\    : AGCBIT;
  signal  \34138\    : AGCBIT;
  signal  \34139\    : AGCBIT;
  signal  \34140\    : AGCBIT; signal  \PA12\     : AGCBIT;
  signal \&34141\    : AGCBIT;
  signal  \34142\    : AGCBIT;
  signal  \34143\    : AGCBIT; signal  \PA12/\    : AGCBIT;
  signal  \34144\    : AGCBIT;
  signal  \34145\    : AGCBIT;
  signal  \34146\    : AGCBIT; signal  \G16A/\    : AGCBIT;
  signal  \34147\    : AGCBIT;
  signal  \34148\    : AGCBIT;
  signal  \34149\    : AGCBIT;
  signal  \34150\    : AGCBIT;
  signal  \34151\    : AGCBIT; signal  \PA15\     : AGCBIT;
  signal \&34152\    : AGCBIT;
  signal  \34153\    : AGCBIT; signal  \PA15/\    : AGCBIT;
  signal  \34154\    : AGCBIT;
  signal  \34155\    : AGCBIT; signal  \GNZRO\    : AGCBIT;
  signal \&34156\    : AGCBIT;
  signal \&34157\    : AGCBIT;
  signal \&34158\    : AGCBIT;
  signal \&34159\    : AGCBIT;
  signal  \34201\    : AGCBIT;
  signal  \34202\    : AGCBIT;
  signal  \34203\    : AGCBIT;
  signal  \34204\    : AGCBIT;
  signal  \34205\    : AGCBIT; signal  \EXTPLS\   : AGCBIT;
  signal  \34206\    : AGCBIT; signal  \RELPLS\   : AGCBIT;
  signal \&34207\    : AGCBIT;
  signal \&34208\    : AGCBIT;
  signal  \34209\    : AGCBIT;
  signal \$34209\    : AGCBIT;
  signal  \34210\    : AGCBIT;
  signal  \34211\    : AGCBIT;
  signal  \34212\    : AGCBIT; signal  \RADRZ\    : AGCBIT;
  signal  \34213\    : AGCBIT; signal  \RADRG\    : AGCBIT;
  signal \&34214\    : AGCBIT;
  signal  \34215\    : AGCBIT; signal  \INHPLS\   : AGCBIT;
  signal  \34216\    : AGCBIT;
  signal \&34217\    : AGCBIT;
  signal  \34218\    : AGCBIT; signal  \GEQZRO/\  : AGCBIT;
  signal  \34219\    : AGCBIT;
  signal  \34220\    : AGCBIT;
  signal  \34221\    : AGCBIT; signal  \EAD09\    : AGCBIT;
  signal  \34222\    : AGCBIT; signal  \EAD10\    : AGCBIT;
  signal  \34223\    : AGCBIT; signal  \EAD11\    : AGCBIT;
  signal  \34224\    : AGCBIT; signal  \EAD09/\   : AGCBIT;
  signal  \34225\    : AGCBIT; signal  \EAD10/\   : AGCBIT;
  signal  \34226\    : AGCBIT; signal  \EAD11/\   : AGCBIT;
  signal  \34227\    : AGCBIT;
  signal  \34228\    : AGCBIT;
  signal  \34229\    : AGCBIT;
  signal  \34230\    : AGCBIT;
  signal  \34231\    : AGCBIT; signal  \PB09\     : AGCBIT;
  signal \&34232\    : AGCBIT;
  signal  \34233\    : AGCBIT; signal  \PB09/\    : AGCBIT;
  signal  \34234\    : AGCBIT;
  signal  \34235\    : AGCBIT;
  signal  \34236\    : AGCBIT; signal  \PB15\     : AGCBIT;
  signal  \34237\    : AGCBIT; signal  \PB15/\    : AGCBIT;
  signal  \34238\    : AGCBIT;
  signal  \34239\    : AGCBIT;
  signal  \34240\    : AGCBIT; signal  \PC15\     : AGCBIT;
  signal \&34241\    : AGCBIT;
  signal  \34242\    : AGCBIT; signal  \PC15/\    : AGCBIT;
  signal \&34243\    : AGCBIT;
  signal \&34244\    : AGCBIT;
  signal  \34245\    : AGCBIT;
  signal \$34245\    : AGCBIT;
  signal  \34246\    : AGCBIT;
  signal  \34247\    : AGCBIT;
  signal  \34248\    : AGCBIT;
  signal \&34250\    : AGCBIT;
  signal  \34251\    : AGCBIT; signal  \PALE\     : AGCBIT;
  signal \&34252\    : AGCBIT;
  signal  \34253\    : AGCBIT; signal  \BRXP3\    : AGCBIT;
  signal \&34254\    : AGCBIT;
  signal  \34301\    : AGCBIT; signal  \G01ED\    : AGCBIT;
  signal  \34302\    : AGCBIT;
  signal  \34303\    : AGCBIT;
  signal \$34303\    : AGCBIT;
  signal  \34304\    : AGCBIT;
  signal  \34306\    : AGCBIT; signal  \S08\      : AGCBIT;
  signal  \34307\    : AGCBIT; signal  \S08/\     : AGCBIT;
  signal  \34309\    : AGCBIT; signal  \G02ED\    : AGCBIT;
  signal  \34310\    : AGCBIT;
  signal  \34311\    : AGCBIT;
  signal \$34311\    : AGCBIT;
  signal  \34312\    : AGCBIT;
  signal  \34314\    : AGCBIT; signal  \S09\      : AGCBIT;
  signal  \34315\    : AGCBIT; signal  \S09/\     : AGCBIT;
  signal  \34317\    : AGCBIT; signal  \G03ED\    : AGCBIT;
  signal  \34318\    : AGCBIT;
  signal  \34319\    : AGCBIT;
  signal \$34319\    : AGCBIT;
  signal  \34320\    : AGCBIT;
  signal  \34322\    : AGCBIT; signal  \S10\      : AGCBIT;
  signal  \34323\    : AGCBIT; signal  \S10/\     : AGCBIT;
  signal  \34325\    : AGCBIT; signal  \G04ED\    : AGCBIT;
  signal  \34326\    : AGCBIT;
  signal  \34327\    : AGCBIT;
  signal \$34327\    : AGCBIT;
  signal  \34328\    : AGCBIT;
  signal  \34329\    : AGCBIT; signal  \T12A\     : AGCBIT;
  signal  \34330\    : AGCBIT; signal  \S11\      : AGCBIT;
  signal  \34331\    : AGCBIT; signal  \S11/\     : AGCBIT;
  signal  \34333\    : AGCBIT; signal  \G05ED\    : AGCBIT;
  signal  \34334\    : AGCBIT;
  signal  \34335\    : AGCBIT;
  signal \$34335\    : AGCBIT;
  signal  \34336\    : AGCBIT;
  signal  \34338\    : AGCBIT; signal  \S12\      : AGCBIT;
  signal  \34339\    : AGCBIT; signal  \S12/\     : AGCBIT;
  signal  \34340\    : AGCBIT; signal  \SHIFT/\   : AGCBIT;
  signal  \34341\    : AGCBIT; signal  \G06ED\    : AGCBIT;
  signal  \34342\    : AGCBIT; signal  \G07ED\    : AGCBIT;
  signal  \34343\    : AGCBIT;
  signal  \34344\    : AGCBIT;
  signal  \34345\    : AGCBIT;
  signal  \34346\    : AGCBIT;
  signal  \34347\    : AGCBIT;
  signal  \34348\    : AGCBIT; signal  \CYR/\     : AGCBIT;
  signal \$34348\    : AGCBIT;
  signal  \34349\    : AGCBIT;
  signal  \34350\    : AGCBIT; signal  \SR/\      : AGCBIT;
  signal \$34350\    : AGCBIT;
  signal  \34351\    : AGCBIT;
  signal  \34352\    : AGCBIT; signal  \CYL/\     : AGCBIT;
  signal \$34352\    : AGCBIT;
  signal  \34353\    : AGCBIT;
  signal  \34354\    : AGCBIT; signal  \EDOP/\    : AGCBIT;
  signal \$34354\    : AGCBIT;
  signal  \34355\    : AGCBIT;
  signal  \34356\    : AGCBIT;
  signal \&34357\    : AGCBIT;
  signal  \34358\    : AGCBIT; signal  \GINH\     : AGCBIT;
  signal  \34362\    : AGCBIT; signal  \SHIFT\    : AGCBIT;
  signal  \34401\    : AGCBIT;
  signal  \34402\    : AGCBIT;
  signal \$34402\    : AGCBIT;
  signal  \34403\    : AGCBIT;
  signal  \34404\    : AGCBIT; signal  \S01\      : AGCBIT;
  signal  \34406\    : AGCBIT; signal  \S01/\     : AGCBIT;
  signal  \34408\    : AGCBIT;
  signal  \34409\    : AGCBIT;
  signal \$34409\    : AGCBIT;
  signal  \34410\    : AGCBIT;
  signal  \34411\    : AGCBIT; signal  \S02\      : AGCBIT;
  signal  \34413\    : AGCBIT; signal  \S02/\     : AGCBIT;
  signal  \34415\    : AGCBIT;
  signal  \34416\    : AGCBIT;
  signal \$34416\    : AGCBIT;
  signal  \34417\    : AGCBIT;
  signal  \34418\    : AGCBIT; signal  \S03\      : AGCBIT;
  signal  \34420\    : AGCBIT; signal  \S03/\     : AGCBIT;
  signal  \34422\    : AGCBIT;
  signal  \34423\    : AGCBIT;
  signal \$34423\    : AGCBIT;
  signal  \34424\    : AGCBIT;
  signal  \34425\    : AGCBIT; signal  \S04\      : AGCBIT;
  signal  \34427\    : AGCBIT; signal  \S04/\     : AGCBIT;
  signal  \34429\    : AGCBIT;
  signal  \34430\    : AGCBIT;
  signal \$34430\    : AGCBIT;
  signal  \34431\    : AGCBIT;
  signal  \34432\    : AGCBIT; signal  \S05\      : AGCBIT;
  signal  \34434\    : AGCBIT; signal  \S05/\     : AGCBIT;
  signal  \34436\    : AGCBIT;
  signal  \34437\    : AGCBIT;
  signal \$34437\    : AGCBIT;
  signal  \34438\    : AGCBIT;
  signal  \34439\    : AGCBIT; signal  \S06\      : AGCBIT;
  signal  \34441\    : AGCBIT; signal  \S06/\     : AGCBIT;
  signal  \34443\    : AGCBIT;
  signal  \34444\    : AGCBIT;
  signal \$34444\    : AGCBIT;
  signal  \34445\    : AGCBIT;
  signal  \34446\    : AGCBIT; signal  \WGA/\     : AGCBIT;
  signal  \34447\    : AGCBIT; signal  \S07\      : AGCBIT;
  signal  \34449\    : AGCBIT; signal  \S07/\     : AGCBIT;
  signal \&34450\    : AGCBIT;
  signal \&34451\    : AGCBIT;
  signal \&34452\    : AGCBIT;
  signal \&34453\    : AGCBIT;
  signal  \34462\    : AGCBIT;
  signal  \34463\    : AGCBIT; signal  \L02A/\    : AGCBIT;
  signal  \34464\    : AGCBIT;
  signal  \34465\    : AGCBIT; signal  \L15A/\    : AGCBIT;
  signal  \34466\    : AGCBIT; signal  \G01A\     : AGCBIT;
  signal  \34467\    : AGCBIT;
  signal  \41101\    : AGCBIT;
  signal  \41102\    : AGCBIT;
  signal  \41103\    : AGCBIT;
  signal \$41103\    : AGCBIT;
  signal  \41104\    : AGCBIT;
  signal \$41104\    : AGCBIT;
  signal  \41105\    : AGCBIT; signal  \MSTRTP\   : AGCBIT;
  signal \&41106\    : AGCBIT;
  signal  \41107\    : AGCBIT;
  signal \$41107\    : AGCBIT;
  signal  \41108\    : AGCBIT;
  signal \$41108\    : AGCBIT;
  signal  \41109\    : AGCBIT;
  signal \$41109\    : AGCBIT;
  signal  \41110\    : AGCBIT;
  signal \$41110\    : AGCBIT;
  signal  \41111\    : AGCBIT;
  signal  \41112\    : AGCBIT;
  signal  \41113\    : AGCBIT;
  signal \&41114\    : AGCBIT;
  signal \&41115\    : AGCBIT;
  signal \&41116\    : AGCBIT;
  signal  \41117\    : AGCBIT; signal  \CKTAL/\   : AGCBIT;
  signal  \41118\    : AGCBIT; signal  \ALGA\     : AGCBIT;
  signal  \41119\    : AGCBIT;
  signal \&41120\    : AGCBIT;
  signal  \41121\    : AGCBIT;
  signal \$41121\    : AGCBIT;
  signal  \41122\    : AGCBIT;
  signal \$41122\    : AGCBIT;
  signal  \41123\    : AGCBIT;
  signal \$41123\    : AGCBIT;
  signal  \41124\    : AGCBIT;
  signal \$41124\    : AGCBIT;
  signal  \41125\    : AGCBIT;
  signal  \41126\    : AGCBIT;
  signal \&41127\    : AGCBIT;
  signal \&41128\    : AGCBIT;
  signal  \41129\    : AGCBIT;
  signal  \41130\    : AGCBIT;
  signal  \41131\    : AGCBIT; signal  \G16SW/\   : AGCBIT;
  signal \&41132\    : AGCBIT;
  signal \&41133\    : AGCBIT;
  signal  \41134\    : AGCBIT; signal  \CTPLS/\   : AGCBIT;
  signal \&41135\    : AGCBIT;
  signal \&41136\    : AGCBIT;
  signal  \41137\    : AGCBIT;
  signal  \41138\    : AGCBIT;
  signal \$41138\    : AGCBIT;
  signal  \41139\    : AGCBIT;
  signal \$41139\    : AGCBIT;
  signal  \41140\    : AGCBIT;
  signal  \41141\    : AGCBIT;
  signal \$41141\    : AGCBIT;
  signal  \41142\    : AGCBIT;
  signal \$41142\    : AGCBIT;
  signal  \41143\    : AGCBIT;
  signal \&41144\    : AGCBIT;
  signal \&41145\    : AGCBIT;
  signal  \41146\    : AGCBIT;
  signal  \41147\    : AGCBIT; signal  \DOFILT\   : AGCBIT;
  signal  \41148\    : AGCBIT;
  signal  \41149\    : AGCBIT;
  signal \$41149\    : AGCBIT;
  signal  \41150\    : AGCBIT;
  signal \$41150\    : AGCBIT;
  signal  \41151\    : AGCBIT;
  signal  \41152\    : AGCBIT;
  signal \$41152\    : AGCBIT;
  signal  \41153\    : AGCBIT;
  signal \$41153\    : AGCBIT;
  signal  \41154\    : AGCBIT; signal  \DLKPLS\   : AGCBIT;
  signal  \41201\    : AGCBIT;
  signal  \41202\    : AGCBIT;
  signal  \41203\    : AGCBIT;
  signal \$41203\    : AGCBIT;
  signal  \41204\    : AGCBIT;
  signal \$41204\    : AGCBIT;
  signal  \41205\    : AGCBIT;
  signal  \41206\    : AGCBIT;
  signal \&41207\    : AGCBIT;
  signal \&41208\    : AGCBIT;
  signal  \41209\    : AGCBIT;
  signal  \41210\    : AGCBIT;
  signal  \41211\    : AGCBIT;
  signal \$41211\    : AGCBIT;
  signal  \41212\    : AGCBIT;
  signal \$41212\    : AGCBIT;
  signal  \41213\    : AGCBIT;
  signal  \41214\    : AGCBIT;
  signal \$41214\    : AGCBIT;
  signal  \41215\    : AGCBIT;
  signal \$41215\    : AGCBIT;
  signal \&41216\    : AGCBIT;
  signal \&41217\    : AGCBIT;
  signal  \41218\    : AGCBIT;
  signal  \41219\    : AGCBIT; signal  \SYNC4/\   : AGCBIT;
  signal  \41220\    : AGCBIT;
  signal  \41221\    : AGCBIT; signal  \SYNC14/\  : AGCBIT;
  signal \&41222\    : AGCBIT;
  signal \&41223\    : AGCBIT;
  signal  \41224\    : AGCBIT;
  signal  \41225\    : AGCBIT;
  signal \$41225\    : AGCBIT;
  signal  \41226\    : AGCBIT; signal  \AGCWAR\   : AGCBIT;
  signal \$41226\    : AGCBIT;
  signal  \41227\    : AGCBIT; signal  \WARN\     : AGCBIT;
  signal  \41228\    : AGCBIT; signal  \CGCWAR\   : AGCBIT;
  signal  \41229\    : AGCBIT;
  signal  \41230\    : AGCBIT; signal  \TMPCAU\   : AGCBIT;
  signal \&41231\    : AGCBIT;
  signal  \41232\    : AGCBIT;
  signal \$41232\    : AGCBIT;
  signal  \41233\    : AGCBIT; signal  \OSCALM\   : AGCBIT;
  signal \$41233\    : AGCBIT;
  signal  \41234\    : AGCBIT;
  signal \$41234\    : AGCBIT;
  signal  \41235\    : AGCBIT;
  signal \$41235\    : AGCBIT;
  signal  \41236\    : AGCBIT; signal  \SBYEXT\   : AGCBIT;
  signal  \41237\    : AGCBIT;
  signal \$41237\    : AGCBIT;
  signal  \41238\    : AGCBIT;
  signal \$41238\    : AGCBIT;
  signal  \41239\    : AGCBIT;
  signal  \41240\    : AGCBIT; signal  \RESTRT\   : AGCBIT;
  signal  \41241\    : AGCBIT; signal  \F08B/\    : AGCBIT;
  signal  \41242\    : AGCBIT; signal  \CON3\     : AGCBIT;
  signal  \41243\    : AGCBIT; signal  \SCADBL\   : AGCBIT;
  signal  \41245\    : AGCBIT;
  signal  \41246\    : AGCBIT; signal  \STRT1\    : AGCBIT;
  signal \$41246\    : AGCBIT;
  signal  \41247\    : AGCBIT;
  signal \$41247\    : AGCBIT;
  signal  \42101\    : AGCBIT; signal  \ROP/\     : AGCBIT;
  signal \&42102\    : AGCBIT;
  signal  \42103\    : AGCBIT;
  signal  \42104\    : AGCBIT;
  signal \$42104\    : AGCBIT;
  signal  \42105\    : AGCBIT;
  signal \$42105\    : AGCBIT;
  signal  \42106\    : AGCBIT;
  signal  \42107\    : AGCBIT;
  signal \$42107\    : AGCBIT;
  signal \&42108\    : AGCBIT;
  signal  \42109\    : AGCBIT;
  signal \$42109\    : AGCBIT;
  signal  \42110\    : AGCBIT;
  signal  \42111\    : AGCBIT;
  signal \$42111\    : AGCBIT;
  signal  \42112\    : AGCBIT;
  signal \$42112\    : AGCBIT;
  signal  \42113\    : AGCBIT;
  signal  \42114\    : AGCBIT;
  signal  \42115\    : AGCBIT;
  signal  \42116\    : AGCBIT; signal  \SETAB/\   : AGCBIT;
  signal  \42117\    : AGCBIT; signal  \SETCD/\   : AGCBIT;
  signal \&42118\    : AGCBIT;
  signal \&42119\    : AGCBIT;
  signal \&42120\    : AGCBIT;
  signal \&42121\    : AGCBIT;
  signal  \42122\    : AGCBIT; signal  \SBFSET\   : AGCBIT;
  signal  \42123\    : AGCBIT;
  signal \$42123\    : AGCBIT;
  signal  \42124\    : AGCBIT; signal  \STBF\     : AGCBIT;
  signal \$42124\    : AGCBIT;
  signal  \42125\    : AGCBIT;
  signal  \42126\    : AGCBIT;
  signal \$42126\    : AGCBIT;
  signal  \42127\    : AGCBIT;
  signal \$42127\    : AGCBIT;
  signal  \42128\    : AGCBIT;
  signal  \42129\    : AGCBIT;
  signal  \42130\    : AGCBIT;
  signal  \42131\    : AGCBIT;
  signal  \42132\    : AGCBIT;
  signal \&42133\    : AGCBIT;
  signal \&42134\    : AGCBIT;
  signal  \42135\    : AGCBIT;
  signal  \42136\    : AGCBIT;
  signal  \42137\    : AGCBIT;
  signal  \42138\    : AGCBIT;
  signal \&42139\    : AGCBIT;
  signal \&42140\    : AGCBIT;
  signal \&42141\    : AGCBIT;
  signal \&42142\    : AGCBIT;
  signal  \42143\    : AGCBIT; signal  \TPGF\     : AGCBIT;
  signal  \42144\    : AGCBIT;
  signal  \42145\    : AGCBIT;
  signal \$42145\    : AGCBIT;
  signal  \42146\    : AGCBIT; signal  \STRGAT\   : AGCBIT;
  signal \$42146\    : AGCBIT;
  signal  \42147\    : AGCBIT;
  signal  \42148\    : AGCBIT;
  signal \&42149\    : AGCBIT;
  signal  \42150\    : AGCBIT;
  signal \$42150\    : AGCBIT;
  signal  \42151\    : AGCBIT;
  signal \$42151\    : AGCBIT;
  signal \&42152\    : AGCBIT;
  signal  \42154\    : AGCBIT;
  signal  \42155\    : AGCBIT;
  signal \$42155\    : AGCBIT;
  signal  \42156\    : AGCBIT;
  signal \$42156\    : AGCBIT;
  signal  \42157\    : AGCBIT; signal  \WHOMPA\   : AGCBIT;
  signal  \42201\    : AGCBIT;
  signal  \42202\    : AGCBIT;
  signal \$42202\    : AGCBIT;
  signal  \42203\    : AGCBIT;
  signal \$42203\    : AGCBIT;
  signal  \42204\    : AGCBIT;
  signal  \42205\    : AGCBIT;
  signal \$42205\    : AGCBIT;
  signal  \42206\    : AGCBIT;
  signal \$42206\    : AGCBIT;
  signal \&42207\    : AGCBIT;
  signal \&42208\    : AGCBIT;
  signal  \42209\    : AGCBIT;
  signal \$42209\    : AGCBIT;
  signal  \42210\    : AGCBIT;
  signal \$42210\    : AGCBIT;
  signal  \42211\    : AGCBIT;
  signal  \42212\    : AGCBIT;
  signal \$42212\    : AGCBIT;
  signal  \42213\    : AGCBIT;
  signal \$42213\    : AGCBIT;
  signal  \42214\    : AGCBIT;
  signal  \42215\    : AGCBIT;
  signal  \42216\    : AGCBIT;
  signal  \42217\    : AGCBIT;
  signal  \42218\    : AGCBIT;
  signal \$42218\    : AGCBIT;
  signal  \42219\    : AGCBIT; signal  \RSTK/\    : AGCBIT;
  signal \$42219\    : AGCBIT;
  signal  \42220\    : AGCBIT;
  signal \$42220\    : AGCBIT;
  signal  \42221\    : AGCBIT;
  signal \$42221\    : AGCBIT;
  signal \&42222\    : AGCBIT;
  signal \&42223\    : AGCBIT;
  signal  \42224\    : AGCBIT;
  signal  \42225\    : AGCBIT; signal  \FNERAS/\  : AGCBIT;
  signal \$42225\    : AGCBIT;
  signal  \42226\    : AGCBIT;
  signal \$42226\    : AGCBIT;
  signal  \42227\    : AGCBIT;
  signal  \42228\    : AGCBIT;
  signal \$42228\    : AGCBIT;
  signal  \42229\    : AGCBIT;
  signal \$42229\    : AGCBIT;
  signal \&42230\    : AGCBIT;
  signal \&42231\    : AGCBIT;
  signal  \42232\    : AGCBIT;
  signal  \42233\    : AGCBIT;
  signal  \42234\    : AGCBIT;
  signal \$42234\    : AGCBIT;
  signal  \42235\    : AGCBIT;
  signal \$42235\    : AGCBIT;
  signal \&42236\    : AGCBIT;
  signal \&42237\    : AGCBIT;
  signal  \42238\    : AGCBIT;
  signal \$42238\    : AGCBIT;
  signal  \42239\    : AGCBIT;
  signal \$42239\    : AGCBIT;
  signal  \42240\    : AGCBIT;
  signal  \42241\    : AGCBIT; signal  \REDRST\   : AGCBIT;
  signal  \42242\    : AGCBIT;
  signal \$42242\    : AGCBIT;
  signal  \42243\    : AGCBIT;
  signal \$42243\    : AGCBIT;
  signal  \42244\    : AGCBIT;
  signal  \42245\    : AGCBIT; signal  \SBESET\   : AGCBIT;
  signal  \42246\    : AGCBIT;
  signal \$42246\    : AGCBIT;
  signal  \42247\    : AGCBIT; signal  \STBE\     : AGCBIT;
  signal \$42247\    : AGCBIT;
  signal  \42248\    : AGCBIT; signal  \TPGE\     : AGCBIT;
  signal  \42249\    : AGCBIT; signal  \TPARG/\   : AGCBIT;
  signal \&42250\    : AGCBIT;
  signal \&42251\    : AGCBIT;
  signal  \42252\    : AGCBIT; signal  \ERAS/\    : AGCBIT;
  signal  \42254\    : AGCBIT; signal  \ERAS\     : AGCBIT;
  signal \&42255\    : AGCBIT;
  signal \&42256\    : AGCBIT;
  signal  \42257\    : AGCBIT; signal  \NOTEST/\  : AGCBIT;
  signal  \42301\    : AGCBIT; signal  \XB0\      : AGCBIT;
  signal  \42302\    : AGCBIT; signal  \XB0/\     : AGCBIT;
  signal \&42306\    : AGCBIT;
  signal  \42307\    : AGCBIT; signal  \XB1\      : AGCBIT;
  signal  \42308\    : AGCBIT; signal  \XB1/\     : AGCBIT;
  signal \&42311\    : AGCBIT;
  signal  \42312\    : AGCBIT; signal  \XB2\      : AGCBIT;
  signal  \42313\    : AGCBIT; signal  \XB2/\     : AGCBIT;
  signal \&42316\    : AGCBIT;
  signal  \42317\    : AGCBIT; signal  \XB3\      : AGCBIT;
  signal  \42318\    : AGCBIT; signal  \XB3/\     : AGCBIT;
  signal \&42321\    : AGCBIT;
  signal  \42322\    : AGCBIT; signal  \XB4\      : AGCBIT;
  signal  \42323\    : AGCBIT; signal  \XB4/\     : AGCBIT;
  signal \&42326\    : AGCBIT;
  signal  \42327\    : AGCBIT; signal  \XB5\      : AGCBIT;
  signal  \42328\    : AGCBIT; signal  \XB5/\     : AGCBIT;
  signal \&42331\    : AGCBIT;
  signal  \42332\    : AGCBIT; signal  \XB6\      : AGCBIT;
  signal  \42333\    : AGCBIT; signal  \XB6/\     : AGCBIT;
  signal \&42336\    : AGCBIT;
  signal  \42337\    : AGCBIT; signal  \XB7\      : AGCBIT;
  signal  \42339\    : AGCBIT; signal  \XB7/\     : AGCBIT;
  signal \&42341\    : AGCBIT;
  signal  \42342\    : AGCBIT; signal  \YB0\      : AGCBIT;
  signal  \42343\    : AGCBIT; signal  \YB0/\     : AGCBIT;
  signal \&42345\    : AGCBIT;
  signal  \42346\    : AGCBIT; signal  \YB1\      : AGCBIT;
  signal  \42347\    : AGCBIT; signal  \YB1/\     : AGCBIT;
  signal \&42348\    : AGCBIT;
  signal  \42349\    : AGCBIT; signal  \YB2\      : AGCBIT;
  signal  \42350\    : AGCBIT; signal  \YB2/\     : AGCBIT;
  signal \&42351\    : AGCBIT;
  signal  \42352\    : AGCBIT; signal  \YB3\      : AGCBIT;
  signal  \42353\    : AGCBIT; signal  \YB3/\     : AGCBIT;
  signal \&42354\    : AGCBIT;
  signal  \42355\    : AGCBIT; signal  \RILP1\    : AGCBIT;
  signal  \42356\    : AGCBIT; signal  \RILP1/\   : AGCBIT;
  signal  \42357\    : AGCBIT; signal  \CXB1/\    : AGCBIT;
  signal  \42401\    : AGCBIT; signal  \XT0\      : AGCBIT;
  signal  \42402\    : AGCBIT; signal  \XT0/\     : AGCBIT;
  signal \&42404\    : AGCBIT;
  signal  \42405\    : AGCBIT; signal  \XT1\      : AGCBIT;
  signal  \42406\    : AGCBIT; signal  \XT1/\     : AGCBIT;
  signal \&42408\    : AGCBIT;
  signal  \42409\    : AGCBIT; signal  \XT2\      : AGCBIT;
  signal  \42410\    : AGCBIT; signal  \XT2/\     : AGCBIT;
  signal \&42412\    : AGCBIT;
  signal  \42413\    : AGCBIT; signal  \XT3\      : AGCBIT;
  signal  \42414\    : AGCBIT; signal  \XT3/\     : AGCBIT;
  signal \&42416\    : AGCBIT;
  signal  \42417\    : AGCBIT; signal  \XT4\      : AGCBIT;
  signal  \42418\    : AGCBIT; signal  \XT4/\     : AGCBIT;
  signal \&42420\    : AGCBIT;
  signal  \42421\    : AGCBIT; signal  \XT5\      : AGCBIT;
  signal  \42423\    : AGCBIT; signal  \XT5/\     : AGCBIT;
  signal \&42424\    : AGCBIT;
  signal  \42425\    : AGCBIT; signal  \XT6\      : AGCBIT;
  signal  \42426\    : AGCBIT; signal  \RB1\      : AGCBIT;
  signal  \42427\    : AGCBIT; signal  \XT6/\     : AGCBIT;
  signal \&42428\    : AGCBIT;
  signal  \42429\    : AGCBIT; signal  \XT7\      : AGCBIT;
  signal  \42431\    : AGCBIT; signal  \XT7/\     : AGCBIT;
  signal \&42432\    : AGCBIT;
  signal  \42433\    : AGCBIT;
  signal \&42434\    : AGCBIT;
  signal  \42435\    : AGCBIT;
  signal  \42436\    : AGCBIT;
  signal  \42437\    : AGCBIT;
  signal  \42438\    : AGCBIT;
  signal  \42439\    : AGCBIT;
  signal  \42440\    : AGCBIT;
  signal \&42441\    : AGCBIT;
  signal  \42442\    : AGCBIT;
  signal  \42443\    : AGCBIT;
  signal \&42444\    : AGCBIT;
  signal  \42445\    : AGCBIT;
  signal \&42446\    : AGCBIT;
  signal \&42447\    : AGCBIT;
  signal  \42448\    : AGCBIT;
  signal  \42449\    : AGCBIT; signal  \RSCG/\    : AGCBIT;
  signal  \42451\    : AGCBIT;
  signal  \42452\    : AGCBIT; signal  \WSCG/\    : AGCBIT;
  signal  \42454\    : AGCBIT; signal  \R1C\      : AGCBIT;
  signal \&42457\    : AGCBIT;
  signal  \42459\    : AGCBIT; signal  \NOTEST\   : AGCBIT;
  signal  \35101\    : AGCBIT;
  signal  \35102\    : AGCBIT; signal  \FB16/\    : AGCBIT;
  signal \$35102\    : AGCBIT;
  signal  \35104\    : AGCBIT; signal  \FB16\     : AGCBIT;
  signal \$35104\    : AGCBIT;
  signal  \35105\    : AGCBIT; signal  \BK16\     : AGCBIT;
  signal \&35106\    : AGCBIT;
  signal  \35107\    : AGCBIT;
  signal  \35108\    : AGCBIT; signal  \FB14/\    : AGCBIT;
  signal \$35108\    : AGCBIT;
  signal  \35110\    : AGCBIT; signal  \FB14\     : AGCBIT;
  signal \$35110\    : AGCBIT;
  signal  \35111\    : AGCBIT;
  signal  \35113\    : AGCBIT;
  signal  \35114\    : AGCBIT; signal  \FB13/\    : AGCBIT;
  signal \$35114\    : AGCBIT;
  signal  \35115\    : AGCBIT; signal  \FB13\     : AGCBIT;
  signal \$35115\    : AGCBIT;
  signal  \35116\    : AGCBIT;
  signal \&35117\    : AGCBIT;
  signal  \35118\    : AGCBIT;
  signal  \35119\    : AGCBIT; signal  \FB12/\    : AGCBIT;
  signal \$35119\    : AGCBIT;
  signal  \35120\    : AGCBIT; signal  \FB12\     : AGCBIT;
  signal \$35120\    : AGCBIT;
  signal  \35121\    : AGCBIT;
  signal \&35122\    : AGCBIT;
  signal  \35123\    : AGCBIT;
  signal  \35124\    : AGCBIT; signal  \FB11/\    : AGCBIT;
  signal \$35124\    : AGCBIT;
  signal  \35125\    : AGCBIT; signal  \FB11\     : AGCBIT;
  signal \$35125\    : AGCBIT;
  signal  \35126\    : AGCBIT;
  signal \&35127\    : AGCBIT;
  signal  \35128\    : AGCBIT;
  signal  \35129\    : AGCBIT;
  signal  \35130\    : AGCBIT; signal  \EB11/\    : AGCBIT;
  signal \$35130\    : AGCBIT;
  signal  \35131\    : AGCBIT; signal  \EB11\     : AGCBIT;
  signal \$35131\    : AGCBIT;
  signal  \35132\    : AGCBIT;
  signal  \35133\    : AGCBIT; signal  \BBK3\     : AGCBIT;
  signal \&35134\    : AGCBIT;
  signal  \35135\    : AGCBIT;
  signal  \35136\    : AGCBIT;
  signal  \35137\    : AGCBIT; signal  \EB10/\    : AGCBIT;
  signal \$35137\    : AGCBIT;
  signal  \35138\    : AGCBIT; signal  \EB10\     : AGCBIT;
  signal \$35138\    : AGCBIT;
  signal  \35139\    : AGCBIT;
  signal  \35140\    : AGCBIT; signal  \BBK2\     : AGCBIT;
  signal \&35141\    : AGCBIT;
  signal \&35142\    : AGCBIT;
  signal  \35143\    : AGCBIT;
  signal  \35144\    : AGCBIT;
  signal  \35145\    : AGCBIT; signal  \EB9/\     : AGCBIT;
  signal \$35145\    : AGCBIT;
  signal  \35146\    : AGCBIT; signal  \EB9\      : AGCBIT;
  signal \$35146\    : AGCBIT;
  signal  \35147\    : AGCBIT;
  signal  \35148\    : AGCBIT; signal  \BBK1\     : AGCBIT;
  signal \&35149\    : AGCBIT;
  signal \&35150\    : AGCBIT;
  signal  \35151\    : AGCBIT;
  signal  \35152\    : AGCBIT;
  signal  \35153\    : AGCBIT;
  signal  \35154\    : AGCBIT;
  signal  \35155\    : AGCBIT;
  signal  \35156\    : AGCBIT;
  signal  \35157\    : AGCBIT;
  signal  \35158\    : AGCBIT;
  signal  \35201\    : AGCBIT;
  signal  \35203\    : AGCBIT;
  signal  \35204\    : AGCBIT;
  signal  \35205\    : AGCBIT; signal  \F11/\     : AGCBIT;
  signal  \35206\    : AGCBIT; signal  \F11\      : AGCBIT;
  signal  \35207\    : AGCBIT; signal  \F13\      : AGCBIT;
  signal  \35208\    : AGCBIT; signal  \F12/\     : AGCBIT;
  signal  \35209\    : AGCBIT; signal  \F12\      : AGCBIT;
  signal  \35210\    : AGCBIT; signal  \F13/\     : AGCBIT;
  signal  \35211\    : AGCBIT;
  signal  \35212\    : AGCBIT;
  signal  \35213\    : AGCBIT; signal  \F16\      : AGCBIT;
  signal \&35214\    : AGCBIT;
  signal  \35215\    : AGCBIT; signal  \F14\      : AGCBIT;
  signal  \35216\    : AGCBIT; signal  \F15\      : AGCBIT;
  signal  \35217\    : AGCBIT; signal  \F14/\     : AGCBIT;
  signal  \35218\    : AGCBIT; signal  \F15/\     : AGCBIT;
  signal  \35219\    : AGCBIT; signal  \F16/\     : AGCBIT;
  signal  \35220\    : AGCBIT;
  signal  \35221\    : AGCBIT;
  signal  \35222\    : AGCBIT;
  signal \$35222\    : AGCBIT;
  signal  \35223\    : AGCBIT;
  signal \$35223\    : AGCBIT;
  signal  \35224\    : AGCBIT;
  signal \$35224\    : AGCBIT;
  signal  \35225\    : AGCBIT;
  signal \$35225\    : AGCBIT;
  signal  \35226\    : AGCBIT; signal  \PRPOR3\   : AGCBIT;
  signal  \35227\    : AGCBIT; signal  \PRPOR4\   : AGCBIT;
  signal \&35228\    : AGCBIT;
  signal  \35229\    : AGCBIT;
  signal \&35230\    : AGCBIT;
  signal  \35231\    : AGCBIT;
  signal  \35232\    : AGCBIT; signal  \RPTAD6\   : AGCBIT;
  signal  \35233\    : AGCBIT; signal  \RPTA12\   : AGCBIT;
  signal  \35234\    : AGCBIT;
  signal \$35234\    : AGCBIT;
  signal  \35235\    : AGCBIT; signal  \RUPTOR/\  : AGCBIT;
  signal \$35235\    : AGCBIT;
  signal  \35236\    : AGCBIT;
  signal \&35237\    : AGCBIT;
  signal  \35238\    : AGCBIT;
  signal  \35239\    : AGCBIT; signal  \MINC/\    : AGCBIT;
  signal \$35239\    : AGCBIT;
  signal  \35240\    : AGCBIT; signal  \MINC\     : AGCBIT;
  signal \$35240\    : AGCBIT;
  signal  \35241\    : AGCBIT;
  signal \&35242\    : AGCBIT;
  signal  \35243\    : AGCBIT;
  signal  \35244\    : AGCBIT; signal  \PCDU/\    : AGCBIT;
  signal \$35244\    : AGCBIT;
  signal  \35245\    : AGCBIT; signal  \PCDU\     : AGCBIT;
  signal \$35245\    : AGCBIT;
  signal  \35246\    : AGCBIT;
  signal \&35247\    : AGCBIT;
  signal  \35248\    : AGCBIT;
  signal  \35249\    : AGCBIT; signal  \MCDU/\    : AGCBIT;
  signal \$35249\    : AGCBIT;
  signal  \35250\    : AGCBIT; signal  \MCDU\     : AGCBIT;
  signal \$35250\    : AGCBIT;
  signal \&35251\    : AGCBIT;
  signal  \35301\    : AGCBIT; signal  \WOVR/\    : AGCBIT;
  signal  \35302\    : AGCBIT;
  signal  \35303\    : AGCBIT;
  signal  \35304\    : AGCBIT; signal  \KRPTA/\   : AGCBIT;
  signal  \35306\    : AGCBIT;
  signal  \35307\    : AGCBIT; signal  \T6RPT\    : AGCBIT;
  signal  \35308\    : AGCBIT;
  signal \$35308\    : AGCBIT;
  signal  \35309\    : AGCBIT;
  signal \$35309\    : AGCBIT;
  signal  \35310\    : AGCBIT;
  signal  \35311\    : AGCBIT;
  signal  \35312\    : AGCBIT;
  signal \$35312\    : AGCBIT;
  signal  \35313\    : AGCBIT;
  signal \$35313\    : AGCBIT;
  signal  \35314\    : AGCBIT;
  signal  \35315\    : AGCBIT;
  signal  \35316\    : AGCBIT;
  signal  \35317\    : AGCBIT;
  signal \$35317\    : AGCBIT;
  signal  \35318\    : AGCBIT;
  signal \$35318\    : AGCBIT;
  signal  \35319\    : AGCBIT;
  signal  \35320\    : AGCBIT;
  signal  \35321\    : AGCBIT;
  signal  \35322\    : AGCBIT;
  signal  \35323\    : AGCBIT;
  signal \$35323\    : AGCBIT;
  signal  \35324\    : AGCBIT;
  signal  \35325\    : AGCBIT;
  signal  \35326\    : AGCBIT;
  signal \$35326\    : AGCBIT;
  signal  \35327\    : AGCBIT; signal  \KY1RST\   : AGCBIT;
  signal  \35328\    : AGCBIT;
  signal \$35328\    : AGCBIT;
  signal  \35329\    : AGCBIT;
  signal \$35329\    : AGCBIT;
  signal  \35330\    : AGCBIT;
  signal  \35331\    : AGCBIT;
  signal  \35332\    : AGCBIT;
  signal  \35333\    : AGCBIT; signal  \KY2RST\   : AGCBIT;
  signal  \35334\    : AGCBIT;
  signal \$35334\    : AGCBIT;
  signal  \35335\    : AGCBIT;
  signal \$35335\    : AGCBIT;
  signal  \35336\    : AGCBIT;
  signal  \35339\    : AGCBIT;
  signal  \35340\    : AGCBIT;
  signal \$35340\    : AGCBIT;
  signal  \35341\    : AGCBIT;
  signal \$35341\    : AGCBIT;
  signal  \35342\    : AGCBIT;
  signal  \35343\    : AGCBIT;
  signal  \35344\    : AGCBIT; signal  \PRPOR1\   : AGCBIT;
  signal  \35345\    : AGCBIT; signal  \DRPRST\   : AGCBIT;
  signal  \35346\    : AGCBIT;
  signal \$35346\    : AGCBIT;
  signal  \35347\    : AGCBIT; signal  \DNRPTA\   : AGCBIT;
  signal \$35347\    : AGCBIT;
  signal  \35348\    : AGCBIT; signal  \PRPOR2\   : AGCBIT;
  signal  \35349\    : AGCBIT; signal  \RRPA1/\   : AGCBIT;
  signal \&35350\    : AGCBIT;
  signal  \35351\    : AGCBIT;
  signal  \35352\    : AGCBIT; signal  \RPTAD3\   : AGCBIT;
  signal \&35353\    : AGCBIT;
  signal  \35354\    : AGCBIT;
  signal  \35355\    : AGCBIT; signal  \RPTAD4\   : AGCBIT;
  signal \&35356\    : AGCBIT;
  signal  \35357\    : AGCBIT;
  signal  \35358\    : AGCBIT; signal  \RPTAD5\   : AGCBIT;
  signal \&35359\    : AGCBIT;
  signal \&35360\    : AGCBIT;
  signal  \35401\    : AGCBIT;
  signal \&35403\    : AGCBIT;
  signal \&35404\    : AGCBIT;
  signal  \35405\    : AGCBIT;
  signal \&35406\    : AGCBIT;
  signal \&35407\    : AGCBIT;
  signal  \35408\    : AGCBIT;
  signal \&35409\    : AGCBIT;
  signal \&35410\    : AGCBIT;
  signal  \35411\    : AGCBIT;
  signal \&35412\    : AGCBIT;
  signal \&35413\    : AGCBIT;
  signal  \35414\    : AGCBIT;
  signal  \35415\    : AGCBIT;
  signal  \35416\    : AGCBIT;
  signal  \35417\    : AGCBIT;
  signal  \35418\    : AGCBIT;
  signal  \35419\    : AGCBIT;
  signal  \35420\    : AGCBIT;
  signal \&35421\    : AGCBIT;
  signal \&35422\    : AGCBIT;
  signal  \35423\    : AGCBIT;
  signal  \35424\    : AGCBIT;
  signal  \35425\    : AGCBIT;
  signal  \35426\    : AGCBIT;
  signal  \35427\    : AGCBIT;
  signal  \35428\    : AGCBIT;
  signal \&35429\    : AGCBIT;
  signal  \35430\    : AGCBIT;
  signal  \35431\    : AGCBIT;
  signal  \35432\    : AGCBIT;
  signal  \35433\    : AGCBIT;
  signal  \35434\    : AGCBIT;
  signal  \35435\    : AGCBIT;
  signal \&35436\    : AGCBIT;
  signal  \35437\    : AGCBIT;
  signal  \35438\    : AGCBIT;
  signal  \35439\    : AGCBIT;
  signal  \35440\    : AGCBIT;
  signal \&35441\    : AGCBIT;
  signal  \35442\    : AGCBIT;
  signal  \35443\    : AGCBIT;
  signal  \35444\    : AGCBIT;
  signal  \35445\    : AGCBIT;
  signal  \35446\    : AGCBIT;
  signal  \35447\    : AGCBIT;
  signal  \35448\    : AGCBIT;
  signal \&35449\    : AGCBIT;
  signal  \35450\    : AGCBIT;
  signal  \35451\    : AGCBIT;
  signal  \35452\    : AGCBIT;
  signal  \35453\    : AGCBIT;
  signal  \35454\    : AGCBIT;
  signal  \35455\    : AGCBIT;
  signal  \35456\    : AGCBIT;
  signal \&35457\    : AGCBIT;
  signal \&35458\    : AGCBIT;
  signal \&35460\    : AGCBIT;
  signal  \43101\    : AGCBIT;
  signal  \43102\    : AGCBIT;
  signal \$43102\    : AGCBIT;
  signal  \43103\    : AGCBIT;
  signal \$43103\    : AGCBIT;
  signal  \43104\    : AGCBIT;
  signal  \43105\    : AGCBIT; signal  \RC+X+P\   : AGCBIT;
  signal \&43106\    : AGCBIT;
  signal  \43107\    : AGCBIT;
  signal  \43108\    : AGCBIT;
  signal \$43108\    : AGCBIT;
  signal  \43109\    : AGCBIT;
  signal \$43109\    : AGCBIT;
  signal  \43110\    : AGCBIT;
  signal  \43111\    : AGCBIT; signal  \RC-X-P\   : AGCBIT;
  signal \&43112\    : AGCBIT;
  signal  \43113\    : AGCBIT;
  signal  \43114\    : AGCBIT;
  signal \$43114\    : AGCBIT;
  signal  \43115\    : AGCBIT;
  signal \$43115\    : AGCBIT;
  signal  \43116\    : AGCBIT;
  signal  \43117\    : AGCBIT; signal  \RC-X+P\   : AGCBIT;
  signal \&43118\    : AGCBIT;
  signal  \43119\    : AGCBIT;
  signal  \43120\    : AGCBIT;
  signal \$43120\    : AGCBIT;
  signal  \43121\    : AGCBIT;
  signal \$43121\    : AGCBIT;
  signal  \43122\    : AGCBIT;
  signal  \43123\    : AGCBIT; signal  \RC+X-P\   : AGCBIT;
  signal \&43124\    : AGCBIT;
  signal  \43125\    : AGCBIT;
  signal  \43126\    : AGCBIT;
  signal \$43126\    : AGCBIT;
  signal  \43127\    : AGCBIT;
  signal \$43127\    : AGCBIT;
  signal  \43128\    : AGCBIT;
  signal  \43129\    : AGCBIT; signal  \RC+X+Y\   : AGCBIT;
  signal \&43130\    : AGCBIT;
  signal  \43131\    : AGCBIT;
  signal  \43132\    : AGCBIT;
  signal \$43132\    : AGCBIT;
  signal  \43133\    : AGCBIT;
  signal \$43133\    : AGCBIT;
  signal  \43134\    : AGCBIT;
  signal  \43135\    : AGCBIT; signal  \RC-X-Y\   : AGCBIT;
  signal \&43136\    : AGCBIT;
  signal  \43137\    : AGCBIT;
  signal  \43138\    : AGCBIT;
  signal \$43138\    : AGCBIT;
  signal  \43139\    : AGCBIT;
  signal \$43139\    : AGCBIT;
  signal  \43140\    : AGCBIT;
  signal  \43141\    : AGCBIT; signal  \RC-X+Y\   : AGCBIT;
  signal \&43142\    : AGCBIT;
  signal  \43143\    : AGCBIT;
  signal  \43144\    : AGCBIT;
  signal \$43144\    : AGCBIT;
  signal  \43145\    : AGCBIT;
  signal \$43145\    : AGCBIT;
  signal  \43146\    : AGCBIT;
  signal  \43147\    : AGCBIT; signal  \RC+X-Y\   : AGCBIT;
  signal \&43148\    : AGCBIT;
  signal  \43149\    : AGCBIT; signal  \WCH05/\   : AGCBIT;
  signal  \43151\    : AGCBIT;
  signal  \43152\    : AGCBIT;
  signal  \43153\    : AGCBIT;
  signal  \43154\    : AGCBIT; signal  \CCH05\    : AGCBIT;
  signal  \43156\    : AGCBIT;
  signal  \43157\    : AGCBIT;
  signal \$43157\    : AGCBIT;
  signal  \43158\    : AGCBIT;
  signal \$43158\    : AGCBIT;
  signal  \43159\    : AGCBIT; signal  \CH1208\   : AGCBIT;
  signal  \43160\    : AGCBIT; signal  \TVCNAB\   : AGCBIT;
  signal  \43201\    : AGCBIT;
  signal  \43202\    : AGCBIT;
  signal \$43202\    : AGCBIT;
  signal  \43203\    : AGCBIT;
  signal \$43203\    : AGCBIT;
  signal  \43204\    : AGCBIT;
  signal  \43205\    : AGCBIT; signal  \RC+Y-R\   : AGCBIT;
  signal  \43206\    : AGCBIT;
  signal  \43207\    : AGCBIT; signal  \WCH06/\   : AGCBIT;
  signal  \43209\    : AGCBIT;
  signal  \43210\    : AGCBIT;
  signal  \43211\    : AGCBIT; signal  \CCH06\    : AGCBIT;
  signal  \43213\    : AGCBIT;
  signal  \43214\    : AGCBIT; signal  \RCH06/\   : AGCBIT;
  signal  \43216\    : AGCBIT;
  signal  \43217\    : AGCBIT; signal  \RCH05/\   : AGCBIT;
  signal  \43219\    : AGCBIT;
  signal  \43220\    : AGCBIT;
  signal \$43220\    : AGCBIT;
  signal  \43221\    : AGCBIT;
  signal \$43221\    : AGCBIT;
  signal  \43222\    : AGCBIT;
  signal  \43223\    : AGCBIT; signal  \RC-Y+R\   : AGCBIT;
  signal  \43224\    : AGCBIT;
  signal  \43225\    : AGCBIT;
  signal \$43225\    : AGCBIT;
  signal  \43226\    : AGCBIT;
  signal \$43226\    : AGCBIT;
  signal  \43227\    : AGCBIT; signal  \CH1207\   : AGCBIT;
  signal  \43228\    : AGCBIT; signal  \OT1207\   : AGCBIT;
  signal  \43229\    : AGCBIT; signal  \OT1207/\  : AGCBIT;
  signal  \43230\    : AGCBIT;
  signal  \43231\    : AGCBIT;
  signal \$43231\    : AGCBIT;
  signal  \43232\    : AGCBIT;
  signal \$43232\    : AGCBIT;
  signal  \43233\    : AGCBIT;
  signal  \43234\    : AGCBIT; signal  \RC-Y-R\   : AGCBIT;
  signal  \43235\    : AGCBIT;
  signal  \43236\    : AGCBIT;
  signal \$43236\    : AGCBIT;
  signal  \43237\    : AGCBIT;
  signal \$43237\    : AGCBIT;
  signal  \43238\    : AGCBIT;
  signal  \43239\    : AGCBIT; signal  \RC+Y+R\   : AGCBIT;
  signal  \43240\    : AGCBIT;
  signal  \43241\    : AGCBIT;
  signal \$43241\    : AGCBIT;
  signal  \43242\    : AGCBIT;
  signal \$43242\    : AGCBIT;
  signal  \43243\    : AGCBIT;
  signal  \43244\    : AGCBIT; signal  \RC+Z-R\   : AGCBIT;
  signal  \43245\    : AGCBIT;
  signal  \43246\    : AGCBIT;
  signal \$43246\    : AGCBIT;
  signal  \43247\    : AGCBIT;
  signal \$43247\    : AGCBIT;
  signal  \43248\    : AGCBIT;
  signal  \43249\    : AGCBIT; signal  \RC-Z+R\   : AGCBIT;
  signal  \43250\    : AGCBIT;
  signal  \43251\    : AGCBIT;
  signal \$43251\    : AGCBIT;
  signal  \43252\    : AGCBIT;
  signal \$43252\    : AGCBIT;
  signal  \43253\    : AGCBIT;
  signal  \43254\    : AGCBIT; signal  \RC-Z-R\   : AGCBIT;
  signal  \43255\    : AGCBIT;
  signal  \43256\    : AGCBIT;
  signal \$43256\    : AGCBIT;
  signal  \43257\    : AGCBIT;
  signal \$43257\    : AGCBIT;
  signal  \43258\    : AGCBIT;
  signal  \43259\    : AGCBIT; signal  \RC+Z+R\   : AGCBIT;
  signal  \43301\    : AGCBIT;
  signal  \43302\    : AGCBIT; signal  \ZOPCDU\   : AGCBIT;
  signal  \43303\    : AGCBIT;
  signal \$43303\    : AGCBIT;
  signal  \43304\    : AGCBIT;
  signal \$43304\    : AGCBIT;
  signal  \43305\    : AGCBIT;
  signal  \43306\    : AGCBIT;
  signal  \43307\    : AGCBIT;
  signal \$43307\    : AGCBIT;
  signal  \43308\    : AGCBIT;
  signal \$43308\    : AGCBIT;
  signal  \43309\    : AGCBIT;
  signal  \43310\    : AGCBIT; signal  \ENEROP\   : AGCBIT;
  signal  \43311\    : AGCBIT;
  signal  \43312\    : AGCBIT; signal  \STARON\   : AGCBIT;
  signal  \43313\    : AGCBIT;
  signal \$43313\    : AGCBIT;
  signal  \43314\    : AGCBIT;
  signal \$43314\    : AGCBIT;
  signal  \43315\    : AGCBIT;
  signal  \43316\    : AGCBIT;
  signal  \43317\    : AGCBIT;
  signal \$43317\    : AGCBIT;
  signal  \43318\    : AGCBIT;
  signal \$43318\    : AGCBIT;
  signal  \43319\    : AGCBIT;
  signal  \43320\    : AGCBIT; signal  \COARSE\   : AGCBIT;
  signal  \43321\    : AGCBIT;
  signal  \43322\    : AGCBIT; signal  \ZIMCDU\   : AGCBIT;
  signal  \43323\    : AGCBIT;
  signal \$43323\    : AGCBIT;
  signal  \43324\    : AGCBIT;
  signal \$43324\    : AGCBIT;
  signal  \43325\    : AGCBIT;
  signal  \43326\    : AGCBIT;
  signal  \43327\    : AGCBIT;
  signal \$43327\    : AGCBIT;
  signal  \43328\    : AGCBIT;
  signal \$43328\    : AGCBIT;
  signal  \43329\    : AGCBIT;
  signal  \43330\    : AGCBIT; signal  \ENERIM\   : AGCBIT;
  signal  \43331\    : AGCBIT; signal  \CH1209\   : AGCBIT;
  signal  \43332\    : AGCBIT; signal  \S4BTAK\   : AGCBIT;
  signal  \43333\    : AGCBIT;
  signal \$43333\    : AGCBIT;
  signal  \43334\    : AGCBIT;
  signal \$43334\    : AGCBIT;
  signal  \43335\    : AGCBIT;
  signal  \43336\    : AGCBIT;
  signal  \43337\    : AGCBIT;
  signal \$43337\    : AGCBIT;
  signal  \43338\    : AGCBIT;
  signal \$43338\    : AGCBIT;
  signal  \43339\    : AGCBIT; signal  \CH1210\   : AGCBIT;
  signal  \43340\    : AGCBIT; signal  \ZEROPT\   : AGCBIT;
  signal  \43341\    : AGCBIT; signal  \CH1211\   : AGCBIT;
  signal  \43342\    : AGCBIT; signal  \DISDAC\   : AGCBIT;
  signal  \43343\    : AGCBIT;
  signal \$43343\    : AGCBIT;
  signal  \43344\    : AGCBIT;
  signal \$43344\    : AGCBIT;
  signal  \43345\    : AGCBIT;
  signal  \43346\    : AGCBIT; signal  \WCH12/\   : AGCBIT;
  signal  \43349\    : AGCBIT;
  signal  \43350\    : AGCBIT;
  signal  \43351\    : AGCBIT;
  signal  \43352\    : AGCBIT; signal  \CCH12\    : AGCBIT;
  signal  \43355\    : AGCBIT;
  signal  \43356\    : AGCBIT; signal  \RCH12/\   : AGCBIT;
  signal  \43401\    : AGCBIT; signal  \ISSWAR\   : AGCBIT;
  signal  \43402\    : AGCBIT;
  signal  \43403\    : AGCBIT;
  signal \$43403\    : AGCBIT;
  signal  \43404\    : AGCBIT;
  signal \$43404\    : AGCBIT;
  signal  \43405\    : AGCBIT;
  signal  \43406\    : AGCBIT;
  signal \&43407\    : AGCBIT;
  signal \&43408\    : AGCBIT;
  signal  \43409\    : AGCBIT;
  signal \$43409\    : AGCBIT;
  signal  \43410\    : AGCBIT;
  signal \$43410\    : AGCBIT;
  signal  \43411\    : AGCBIT;
  signal  \43412\    : AGCBIT; signal  \COMACT\   : AGCBIT;
  signal  \43413\    : AGCBIT; signal  \UPLACT\   : AGCBIT;
  signal  \43414\    : AGCBIT;
  signal  \43415\    : AGCBIT;
  signal \$43415\    : AGCBIT;
  signal  \43416\    : AGCBIT;
  signal \$43416\    : AGCBIT;
  signal  \43417\    : AGCBIT;
  signal  \43418\    : AGCBIT;
  signal \&43419\    : AGCBIT;
  signal \&43420\    : AGCBIT;
  signal  \43421\    : AGCBIT;
  signal \$43421\    : AGCBIT;
  signal  \43422\    : AGCBIT;
  signal \$43422\    : AGCBIT;
  signal  \43423\    : AGCBIT;
  signal  \43424\    : AGCBIT; signal  \TMPOUT\   : AGCBIT;
  signal \&43425\    : AGCBIT;
  signal \&43426\    : AGCBIT;
  signal  \43427\    : AGCBIT; signal  \KYRLS\    : AGCBIT;
  signal  \43428\    : AGCBIT;
  signal  \43429\    : AGCBIT;
  signal \$43429\    : AGCBIT;
  signal  \43430\    : AGCBIT;
  signal \$43430\    : AGCBIT;
  signal  \43431\    : AGCBIT;
  signal  \43432\    : AGCBIT;
  signal  \43433\    : AGCBIT;
  signal \$43433\    : AGCBIT;
  signal  \43434\    : AGCBIT;
  signal \$43434\    : AGCBIT;
  signal  \43435\    : AGCBIT; signal  \VNFLSH\   : AGCBIT;
  signal  \43436\    : AGCBIT;
  signal \&43437\    : AGCBIT;
  signal \&43438\    : AGCBIT;
  signal \&43439\    : AGCBIT;
  signal \&43440\    : AGCBIT;
  signal  \43441\    : AGCBIT; signal  \OPEROR\   : AGCBIT;
  signal  \43442\    : AGCBIT;
  signal  \43443\    : AGCBIT;
  signal \$43443\    : AGCBIT;
  signal  \43444\    : AGCBIT;
  signal \$43444\    : AGCBIT;
  signal  \43445\    : AGCBIT;
  signal  \43446\    : AGCBIT;
  signal  \43447\    : AGCBIT;
  signal \$43447\    : AGCBIT;
  signal  \43448\    : AGCBIT;
  signal \$43448\    : AGCBIT;
  signal  \43449\    : AGCBIT; signal  \CH1212\   : AGCBIT;
  signal  \43450\    : AGCBIT; signal  \MROLGT\   : AGCBIT;
  signal  \43451\    : AGCBIT; signal  \S4BSEQ\   : AGCBIT;
  signal  \43452\    : AGCBIT; signal  \CH1213\   : AGCBIT;
  signal  \43453\    : AGCBIT;
  signal \$43453\    : AGCBIT;
  signal  \43454\    : AGCBIT;
  signal \$43454\    : AGCBIT;
  signal  \43455\    : AGCBIT;
  signal  \43456\    : AGCBIT;
  signal  \43457\    : AGCBIT;
  signal \$43457\    : AGCBIT;
  signal  \43458\    : AGCBIT;
  signal \$43458\    : AGCBIT;
  signal  \43459\    : AGCBIT; signal  \CH1214\   : AGCBIT;
  signal  \43460\    : AGCBIT; signal  \S4BOFF\   : AGCBIT;
  signal  \44101\    : AGCBIT;
  signal  \44102\    : AGCBIT;
  signal  \44103\    : AGCBIT; signal  \CHOR01/\  : AGCBIT;
  signal  \44104\    : AGCBIT;
  signal  \44105\    : AGCBIT;
  signal  \44106\    : AGCBIT; signal  \CHOR02/\  : AGCBIT;
  signal  \44107\    : AGCBIT;
  signal  \44108\    : AGCBIT;
  signal  \44109\    : AGCBIT; signal  \CHOR03/\  : AGCBIT;
  signal  \44110\    : AGCBIT;
  signal  \44111\    : AGCBIT;
  signal  \44112\    : AGCBIT; signal  \CHOR04/\  : AGCBIT;
  signal  \44113\    : AGCBIT;
  signal  \44114\    : AGCBIT;
  signal  \44115\    : AGCBIT; signal  \CHOR05/\  : AGCBIT;
  signal  \44116\    : AGCBIT;
  signal  \44117\    : AGCBIT;
  signal  \44118\    : AGCBIT; signal  \CHOR06/\  : AGCBIT;
  signal  \44119\    : AGCBIT;
  signal  \44120\    : AGCBIT;
  signal  \44121\    : AGCBIT; signal  \CHOR07/\  : AGCBIT;
  signal  \44122\    : AGCBIT;
  signal  \44123\    : AGCBIT;
  signal  \44124\    : AGCBIT; signal  \CHOR08/\  : AGCBIT;
  signal  \44125\    : AGCBIT;
  signal  \44126\    : AGCBIT;
  signal  \44127\    : AGCBIT; signal  \CHOR09/\  : AGCBIT;
  signal  \44128\    : AGCBIT;
  signal  \44129\    : AGCBIT; signal  \CHOR10/\  : AGCBIT;
  signal  \44130\    : AGCBIT;
  signal  \44131\    : AGCBIT;
  signal  \44132\    : AGCBIT; signal  \CHOR11/\  : AGCBIT;
  signal  \44133\    : AGCBIT;
  signal  \44134\    : AGCBIT;
  signal  \44135\    : AGCBIT; signal  \CHOR12/\  : AGCBIT;
  signal  \44136\    : AGCBIT;
  signal  \44137\    : AGCBIT;
  signal  \44138\    : AGCBIT; signal  \CHOR13/\  : AGCBIT;
  signal  \44139\    : AGCBIT;
  signal  \44140\    : AGCBIT;
  signal  \44141\    : AGCBIT; signal  \CHOR14/\  : AGCBIT;
  signal  \44142\    : AGCBIT;
  signal  \44143\    : AGCBIT;
  signal  \44144\    : AGCBIT; signal  \CHOR16/\  : AGCBIT;
  signal  \44145\    : AGCBIT;
  signal  \44146\    : AGCBIT; signal  \RCH30/\   : AGCBIT;
  signal  \44149\    : AGCBIT;
  signal  \44150\    : AGCBIT; signal  \RCH31/\   : AGCBIT;
  signal  \44153\    : AGCBIT;
  signal  \44154\    : AGCBIT; signal  \RCH32/\   : AGCBIT;
  signal  \44157\    : AGCBIT;
  signal  \44158\    : AGCBIT; signal  \RCH33/\   : AGCBIT;
  signal  \44201\    : AGCBIT;
  signal  \44202\    : AGCBIT;
  signal  \44203\    : AGCBIT;
  signal  \44204\    : AGCBIT;
  signal  \44205\    : AGCBIT;
  signal  \44206\    : AGCBIT;
  signal \&44207\    : AGCBIT;
  signal  \44208\    : AGCBIT;
  signal  \44209\    : AGCBIT;
  signal \$44209\    : AGCBIT;
  signal  \44210\    : AGCBIT;
  signal \$44210\    : AGCBIT;
  signal  \44211\    : AGCBIT; signal  \TRP31A\   : AGCBIT;
  signal  \44212\    : AGCBIT;
  signal \$44212\    : AGCBIT;
  signal  \44213\    : AGCBIT;
  signal \$44213\    : AGCBIT;
  signal  \44214\    : AGCBIT;
  signal  \44215\    : AGCBIT;
  signal  \44216\    : AGCBIT;
  signal  \44217\    : AGCBIT;
  signal  \44218\    : AGCBIT;
  signal  \44219\    : AGCBIT;
  signal  \44220\    : AGCBIT;
  signal  \44221\    : AGCBIT;
  signal \&44222\    : AGCBIT;
  signal  \44223\    : AGCBIT;
  signal  \44224\    : AGCBIT;
  signal \$44224\    : AGCBIT;
  signal  \44225\    : AGCBIT;
  signal \$44225\    : AGCBIT;
  signal  \44226\    : AGCBIT; signal  \TRP31B\   : AGCBIT;
  signal  \44227\    : AGCBIT;
  signal  \44228\    : AGCBIT;
  signal \$44228\    : AGCBIT;
  signal  \44229\    : AGCBIT;
  signal \$44229\    : AGCBIT;
  signal  \44230\    : AGCBIT;
  signal  \44231\    : AGCBIT; signal  \HNDRPT\   : AGCBIT;
  signal  \44232\    : AGCBIT;
  signal  \44233\    : AGCBIT;
  signal  \44234\    : AGCBIT;
  signal  \44235\    : AGCBIT;
  signal  \44236\    : AGCBIT; signal  \CH3201\   : AGCBIT;
  signal  \44237\    : AGCBIT; signal  \CH3206\   : AGCBIT;
  signal  \44238\    : AGCBIT; signal  \CH3202\   : AGCBIT;
  signal  \44239\    : AGCBIT; signal  \CH3207\   : AGCBIT;
  signal  \44240\    : AGCBIT; signal  \CH3203\   : AGCBIT;
  signal  \44241\    : AGCBIT; signal  \CH3208\   : AGCBIT;
  signal  \44242\    : AGCBIT; signal  \CH3204\   : AGCBIT;
  signal  \44243\    : AGCBIT; signal  \CH3209\   : AGCBIT;
  signal  \44244\    : AGCBIT; signal  \CH3205\   : AGCBIT;
  signal  \44245\    : AGCBIT; signal  \CH3210\   : AGCBIT;
  signal \&44246\    : AGCBIT;
  signal \&44247\    : AGCBIT;
  signal  \44248\    : AGCBIT;
  signal \&44249\    : AGCBIT;
  signal  \44250\    : AGCBIT;
  signal  \44251\    : AGCBIT;
  signal \$44251\    : AGCBIT;
  signal  \44252\    : AGCBIT;
  signal \$44252\    : AGCBIT;
  signal  \44253\    : AGCBIT; signal  \TRP32\    : AGCBIT;
  signal  \44254\    : AGCBIT;
  signal \$44254\    : AGCBIT;
  signal  \44255\    : AGCBIT;
  signal \$44255\    : AGCBIT;
  signal  \44256\    : AGCBIT;
  signal  \44257\    : AGCBIT; signal  \CH3316\   : AGCBIT;
  signal  \44258\    : AGCBIT; signal  \CH3314\   : AGCBIT;
  signal  \44259\    : AGCBIT; signal  \CH3313\   : AGCBIT;
  signal  \44301\    : AGCBIT;
  signal  \44302\    : AGCBIT;
  signal \$44302\    : AGCBIT;
  signal  \44303\    : AGCBIT;
  signal \$44303\    : AGCBIT;
  signal  \44304\    : AGCBIT;
  signal  \44305\    : AGCBIT; signal  \RLYB01\   : AGCBIT;
  signal \&44306\    : AGCBIT;
  signal  \44307\    : AGCBIT;
  signal  \44308\    : AGCBIT;
  signal \$44308\    : AGCBIT;
  signal  \44309\    : AGCBIT;
  signal \$44309\    : AGCBIT;
  signal  \44310\    : AGCBIT;
  signal  \44311\    : AGCBIT; signal  \RLYB02\   : AGCBIT;
  signal \&44312\    : AGCBIT;
  signal  \44313\    : AGCBIT;
  signal  \44314\    : AGCBIT;
  signal \$44314\    : AGCBIT;
  signal  \44315\    : AGCBIT;
  signal \$44315\    : AGCBIT;
  signal  \44316\    : AGCBIT;
  signal  \44317\    : AGCBIT; signal  \RLYB03\   : AGCBIT;
  signal \&44318\    : AGCBIT;
  signal  \44319\    : AGCBIT;
  signal  \44320\    : AGCBIT;
  signal \$44320\    : AGCBIT;
  signal  \44321\    : AGCBIT;
  signal \$44321\    : AGCBIT;
  signal  \44322\    : AGCBIT;
  signal  \44323\    : AGCBIT; signal  \RLYB04\   : AGCBIT;
  signal \&44324\    : AGCBIT;
  signal  \44325\    : AGCBIT;
  signal  \44326\    : AGCBIT;
  signal \$44326\    : AGCBIT;
  signal  \44327\    : AGCBIT;
  signal \$44327\    : AGCBIT;
  signal  \44328\    : AGCBIT;
  signal  \44329\    : AGCBIT; signal  \RLYB05\   : AGCBIT;
  signal \&44330\    : AGCBIT;
  signal  \44331\    : AGCBIT;
  signal  \44332\    : AGCBIT;
  signal \$44332\    : AGCBIT;
  signal  \44333\    : AGCBIT;
  signal \$44333\    : AGCBIT;
  signal  \44334\    : AGCBIT;
  signal  \44335\    : AGCBIT; signal  \RLYB06\   : AGCBIT;
  signal \&44336\    : AGCBIT;
  signal  \44337\    : AGCBIT;
  signal  \44338\    : AGCBIT;
  signal \$44338\    : AGCBIT;
  signal  \44339\    : AGCBIT;
  signal \$44339\    : AGCBIT;
  signal  \44340\    : AGCBIT;
  signal  \44341\    : AGCBIT; signal  \RLYB07\   : AGCBIT;
  signal \&44342\    : AGCBIT;
  signal  \44343\    : AGCBIT;
  signal  \44344\    : AGCBIT;
  signal \$44344\    : AGCBIT;
  signal  \44345\    : AGCBIT;
  signal \$44345\    : AGCBIT;
  signal  \44346\    : AGCBIT;
  signal  \44347\    : AGCBIT; signal  \RLYB08\   : AGCBIT;
  signal \&44348\    : AGCBIT;
  signal  \44349\    : AGCBIT;
  signal  \44350\    : AGCBIT;
  signal \$44350\    : AGCBIT;
  signal  \44351\    : AGCBIT;
  signal \$44351\    : AGCBIT;
  signal  \44352\    : AGCBIT;
  signal  \44353\    : AGCBIT; signal  \RLYB09\   : AGCBIT;
  signal \&44354\    : AGCBIT;
  signal  \44355\    : AGCBIT;
  signal  \44356\    : AGCBIT;
  signal \$44356\    : AGCBIT;
  signal  \44357\    : AGCBIT;
  signal \$44357\    : AGCBIT;
  signal  \44358\    : AGCBIT;
  signal  \44359\    : AGCBIT; signal  \RLYB10\   : AGCBIT;
  signal \&44360\    : AGCBIT;
  signal  \44401\    : AGCBIT;
  signal  \44402\    : AGCBIT;
  signal \$44402\    : AGCBIT;
  signal  \44403\    : AGCBIT;
  signal \$44403\    : AGCBIT;
  signal  \44404\    : AGCBIT;
  signal  \44405\    : AGCBIT; signal  \RLYB11\   : AGCBIT;
  signal \&44406\    : AGCBIT;
  signal  \44407\    : AGCBIT;
  signal  \44408\    : AGCBIT;
  signal \$44408\    : AGCBIT;
  signal  \44409\    : AGCBIT;
  signal \$44409\    : AGCBIT;
  signal  \44410\    : AGCBIT;
  signal  \44411\    : AGCBIT; signal  \RYWD12\   : AGCBIT;
  signal \&44412\    : AGCBIT;
  signal  \44413\    : AGCBIT;
  signal  \44414\    : AGCBIT;
  signal \$44414\    : AGCBIT;
  signal  \44415\    : AGCBIT;
  signal \$44415\    : AGCBIT;
  signal  \44416\    : AGCBIT;
  signal  \44417\    : AGCBIT; signal  \RYWD13\   : AGCBIT;
  signal \&44418\    : AGCBIT;
  signal  \44419\    : AGCBIT;
  signal  \44420\    : AGCBIT;
  signal \$44420\    : AGCBIT;
  signal  \44421\    : AGCBIT;
  signal \$44421\    : AGCBIT;
  signal  \44422\    : AGCBIT;
  signal  \44423\    : AGCBIT; signal  \RYWD14\   : AGCBIT;
  signal \&44424\    : AGCBIT;
  signal  \44425\    : AGCBIT;
  signal  \44426\    : AGCBIT;
  signal \$44426\    : AGCBIT;
  signal  \44427\    : AGCBIT;
  signal \$44427\    : AGCBIT;
  signal  \44428\    : AGCBIT;
  signal  \44429\    : AGCBIT; signal  \RYWD16\   : AGCBIT;
  signal \&44430\    : AGCBIT;
  signal  \44431\    : AGCBIT;
  signal  \44432\    : AGCBIT; signal  \WCH10/\   : AGCBIT;
  signal  \44435\    : AGCBIT;
  signal  \44436\    : AGCBIT;
  signal  \44437\    : AGCBIT; signal  \CCH10\    : AGCBIT;
  signal  \44440\    : AGCBIT;
  signal  \44441\    : AGCBIT; signal  \RCH10/\   : AGCBIT;
  signal  \44444\    : AGCBIT;
  signal  \44445\    : AGCBIT; signal  \WCH11/\   : AGCBIT;
  signal  \44448\    : AGCBIT;
  signal  \44449\    : AGCBIT;
  signal  \44450\    : AGCBIT; signal  \CCH11\    : AGCBIT;
  signal  \44453\    : AGCBIT;
  signal  \44454\    : AGCBIT; signal  \RCH11/\   : AGCBIT;
  signal \&44461\    : AGCBIT;
  signal  \44462\    : AGCBIT; signal  \XBC\      : AGCBIT;
  signal  \45101\    : AGCBIT;
  signal \$45101\    : AGCBIT;
  signal  \45102\    : AGCBIT;
  signal \$45102\    : AGCBIT;
  signal  \45103\    : AGCBIT; signal  \CH1501\   : AGCBIT;
  signal  \45104\    : AGCBIT;
  signal  \45105\    : AGCBIT;
  signal \$45105\    : AGCBIT;
  signal  \45106\    : AGCBIT;
  signal \$45106\    : AGCBIT;
  signal  \45107\    : AGCBIT; signal  \CH1502\   : AGCBIT;
  signal  \45108\    : AGCBIT;
  signal  \45109\    : AGCBIT;
  signal \$45109\    : AGCBIT;
  signal  \45110\    : AGCBIT;
  signal \$45110\    : AGCBIT;
  signal  \45111\    : AGCBIT; signal  \CH1503\   : AGCBIT;
  signal  \45112\    : AGCBIT;
  signal  \45113\    : AGCBIT;
  signal \$45113\    : AGCBIT;
  signal  \45114\    : AGCBIT;
  signal \$45114\    : AGCBIT;
  signal  \45115\    : AGCBIT; signal  \CH1504\   : AGCBIT;
  signal  \45116\    : AGCBIT;
  signal  \45117\    : AGCBIT;
  signal \$45117\    : AGCBIT;
  signal  \45118\    : AGCBIT;
  signal \$45118\    : AGCBIT;
  signal  \45119\    : AGCBIT; signal  \CH1505\   : AGCBIT;
  signal  \45120\    : AGCBIT;
  signal  \45121\    : AGCBIT;
  signal  \45122\    : AGCBIT;
  signal  \45123\    : AGCBIT;
  signal  \45124\    : AGCBIT; signal  \RCH15/\   : AGCBIT;
  signal \&45125\    : AGCBIT;
  signal  \45126\    : AGCBIT;
  signal  \45127\    : AGCBIT;
  signal  \45128\    : AGCBIT; signal  \TPOR/\    : AGCBIT;
  signal  \45129\    : AGCBIT;
  signal \$45129\    : AGCBIT;
  signal  \45130\    : AGCBIT;
  signal \$45130\    : AGCBIT;
  signal  \45131\    : AGCBIT; signal  \KYRPT1\   : AGCBIT;
  signal \&45132\    : AGCBIT;
  signal  \45133\    : AGCBIT;
  signal  \45134\    : AGCBIT;
  signal  \45135\    : AGCBIT;
  signal \$45135\    : AGCBIT;
  signal  \45136\    : AGCBIT;
  signal \$45136\    : AGCBIT;
  signal  \45137\    : AGCBIT;
  signal  \45138\    : AGCBIT;
  signal \$45138\    : AGCBIT;
  signal  \45139\    : AGCBIT;
  signal \$45139\    : AGCBIT;
  signal  \45140\    : AGCBIT; signal  \CH1311\   : AGCBIT;
  signal  \45141\    : AGCBIT;
  signal  \45142\    : AGCBIT;
  signal \$45142\    : AGCBIT;
  signal  \45143\    : AGCBIT;
  signal  \45144\    : AGCBIT;
  signal \$45144\    : AGCBIT;
  signal  \45145\    : AGCBIT;
  signal \$45145\    : AGCBIT;
  signal  \45146\    : AGCBIT;
  signal \$45146\    : AGCBIT;
  signal  \45147\    : AGCBIT;
  signal  \45148\    : AGCBIT; signal  \SBY\      : AGCBIT;
  signal  \45149\    : AGCBIT;
  signal  \45150\    : AGCBIT;
  signal \$45150\    : AGCBIT;
  signal  \45151\    : AGCBIT;
  signal \$45151\    : AGCBIT;
  signal  \45152\    : AGCBIT;
  signal  \45153\    : AGCBIT; signal  \STNDBY/\  : AGCBIT;
  signal  \45154\    : AGCBIT;
  signal \$45154\    : AGCBIT;
  signal  \45155\    : AGCBIT; signal  \STNDBY\   : AGCBIT;
  signal \$45155\    : AGCBIT;
  signal  \45156\    : AGCBIT;
  signal  \45157\    : AGCBIT; signal  \SBYLIT\   : AGCBIT;
  signal  \45159\    : AGCBIT; signal  \F17A/\    : AGCBIT;
  signal \&45160\    : AGCBIT;
  signal  \45201\    : AGCBIT;
  signal \$45201\    : AGCBIT;
  signal  \45202\    : AGCBIT;
  signal \$45202\    : AGCBIT;
  signal  \45203\    : AGCBIT; signal  \CH1601\   : AGCBIT;
  signal  \45204\    : AGCBIT;
  signal  \45205\    : AGCBIT;
  signal \$45205\    : AGCBIT;
  signal  \45206\    : AGCBIT;
  signal \$45206\    : AGCBIT;
  signal  \45207\    : AGCBIT; signal  \CH1602\   : AGCBIT;
  signal  \45208\    : AGCBIT;
  signal  \45209\    : AGCBIT;
  signal \$45209\    : AGCBIT;
  signal  \45210\    : AGCBIT;
  signal \$45210\    : AGCBIT;
  signal  \45211\    : AGCBIT; signal  \CH1603\   : AGCBIT;
  signal  \45212\    : AGCBIT;
  signal  \45213\    : AGCBIT;
  signal \$45213\    : AGCBIT;
  signal  \45214\    : AGCBIT;
  signal \$45214\    : AGCBIT;
  signal  \45215\    : AGCBIT; signal  \CH1604\   : AGCBIT;
  signal  \45216\    : AGCBIT;
  signal  \45217\    : AGCBIT;
  signal \$45217\    : AGCBIT;
  signal  \45218\    : AGCBIT;
  signal \$45218\    : AGCBIT;
  signal  \45219\    : AGCBIT; signal  \CH1605\   : AGCBIT;
  signal  \45220\    : AGCBIT;
  signal  \45221\    : AGCBIT;
  signal  \45222\    : AGCBIT;
  signal  \45223\    : AGCBIT;
  signal  \45224\    : AGCBIT; signal  \ERRST\    : AGCBIT;
  signal  \45225\    : AGCBIT;
  signal \$45225\    : AGCBIT;
  signal  \45226\    : AGCBIT;
  signal \$45226\    : AGCBIT;
  signal  \45227\    : AGCBIT; signal  \CH1606\   : AGCBIT;
  signal  \45228\    : AGCBIT;
  signal  \45229\    : AGCBIT;
  signal \$45229\    : AGCBIT;
  signal  \45230\    : AGCBIT;
  signal \$45230\    : AGCBIT;
  signal  \45231\    : AGCBIT; signal  \CH1607\   : AGCBIT;
  signal  \45232\    : AGCBIT;
  signal  \45233\    : AGCBIT;
  signal  \45234\    : AGCBIT;
  signal  \45235\    : AGCBIT;
  signal  \45236\    : AGCBIT; signal  \RCH16/\   : AGCBIT;
  signal \&45238\    : AGCBIT;
  signal  \45239\    : AGCBIT;
  signal  \45240\    : AGCBIT;
  signal  \45241\    : AGCBIT;
  signal \$45241\    : AGCBIT;
  signal  \45242\    : AGCBIT;
  signal \$45242\    : AGCBIT;
  signal \&45243\    : AGCBIT;
  signal  \45244\    : AGCBIT; signal  \KYRPT2\   : AGCBIT;
  signal  \45245\    : AGCBIT;
  signal  \45246\    : AGCBIT;
  signal  \45247\    : AGCBIT;
  signal \$45247\    : AGCBIT;
  signal  \45248\    : AGCBIT;
  signal \$45248\    : AGCBIT;
  signal  \45249\    : AGCBIT;
  signal  \45250\    : AGCBIT;
  signal  \45251\    : AGCBIT;
  signal \$45251\    : AGCBIT;
  signal  \45252\    : AGCBIT;
  signal \$45252\    : AGCBIT;
  signal  \45254\    : AGCBIT; signal  \MKRPT\    : AGCBIT;
  signal  \45255\    : AGCBIT;
  signal  \45256\    : AGCBIT;
  signal  \45257\    : AGCBIT;
  signal \$45257\    : AGCBIT;
  signal  \45258\    : AGCBIT;
  signal \$45258\    : AGCBIT;
  signal  \45261\    : AGCBIT; signal  \F17B/\    : AGCBIT;
  signal  \45262\    : AGCBIT; signal  \TEMPIN/\  : AGCBIT;
  signal  \45301\    : AGCBIT;
  signal  \45302\    : AGCBIT;
  signal \$45302\    : AGCBIT;
  signal  \45303\    : AGCBIT;
  signal \$45303\    : AGCBIT;
  signal  \45304\    : AGCBIT; signal  \CH1304\   : AGCBIT;
  signal  \45305\    : AGCBIT;
  signal  \45306\    : AGCBIT;
  signal  \45307\    : AGCBIT;
  signal \$45307\    : AGCBIT;
  signal  \45308\    : AGCBIT;
  signal \$45308\    : AGCBIT;
  signal  \45309\    : AGCBIT; signal  \CH1303\   : AGCBIT;
  signal  \45310\    : AGCBIT;
  signal  \45311\    : AGCBIT;
  signal  \45312\    : AGCBIT;
  signal  \45313\    : AGCBIT;
  signal \$45313\    : AGCBIT;
  signal  \45314\    : AGCBIT;
  signal \$45314\    : AGCBIT;
  signal  \45315\    : AGCBIT; signal  \CH1302\   : AGCBIT;
  signal  \45316\    : AGCBIT;
  signal  \45317\    : AGCBIT;
  signal \$45317\    : AGCBIT;
  signal  \45318\    : AGCBIT;
  signal \$45318\    : AGCBIT;
  signal  \45319\    : AGCBIT; signal  \CH1301\   : AGCBIT;
  signal  \45320\    : AGCBIT;
  signal \$45320\    : AGCBIT;
  signal  \45321\    : AGCBIT;
  signal \$45321\    : AGCBIT;
  signal  \45322\    : AGCBIT;
  signal  \45323\    : AGCBIT;
  signal  \45324\    : AGCBIT;
  signal  \45325\    : AGCBIT;
  signal  \45326\    : AGCBIT;
  signal  \45327\    : AGCBIT;
  signal  \45328\    : AGCBIT; signal  \RRRANG\   : AGCBIT;
  signal  \45329\    : AGCBIT; signal  \RRRARA\   : AGCBIT;
  signal  \45330\    : AGCBIT; signal  \LRXVEL\   : AGCBIT;
  signal  \45331\    : AGCBIT; signal  \LRYVEL\   : AGCBIT;
  signal  \45332\    : AGCBIT; signal  \LRZVEL\   : AGCBIT;
  signal  \45333\    : AGCBIT; signal  \LRRANG\   : AGCBIT;
  signal  \45334\    : AGCBIT;
  signal  \45335\    : AGCBIT;
  signal  \45336\    : AGCBIT;
  signal  \45337\    : AGCBIT;
  signal \$45337\    : AGCBIT;
  signal  \45338\    : AGCBIT;
  signal \$45338\    : AGCBIT;
  signal  \45339\    : AGCBIT;
  signal  \45340\    : AGCBIT;
  signal \$45340\    : AGCBIT;
  signal  \45341\    : AGCBIT;
  signal \$45341\    : AGCBIT;
  signal  \45342\    : AGCBIT; signal  \RADRPT\   : AGCBIT;
  signal \&45343\    : AGCBIT;
  signal  \45344\    : AGCBIT;
  signal  \45345\    : AGCBIT; signal  \RRSYNC\   : AGCBIT;
  signal  \45346\    : AGCBIT; signal  \LRSYNC\   : AGCBIT;
  signal  \45347\    : AGCBIT;
  signal  \45348\    : AGCBIT;
  signal  \45349\    : AGCBIT;
  signal  \45350\    : AGCBIT;
  signal  \45351\    : AGCBIT;
  signal  \45352\    : AGCBIT; signal  \RNRADP\   : AGCBIT;
  signal  \45353\    : AGCBIT;
  signal  \45354\    : AGCBIT;
  signal  \45355\    : AGCBIT;
  signal  \45356\    : AGCBIT;
  signal  \45357\    : AGCBIT;
  signal  \45358\    : AGCBIT; signal  \RNRADM\   : AGCBIT;
  signal  \45359\    : AGCBIT; signal  \TPORA/\   : AGCBIT;
  signal  \45360\    : AGCBIT; signal  \HERB\     : AGCBIT;
  signal  \45401\    : AGCBIT; signal  \F10AS0\   : AGCBIT;
  signal  \45402\    : AGCBIT;
  signal \$45402\    : AGCBIT;
  signal  \45403\    : AGCBIT;
  signal \$45403\    : AGCBIT;
  signal  \45404\    : AGCBIT;
  signal  \45405\    : AGCBIT;
  signal \$45405\    : AGCBIT;
  signal \&45406\    : AGCBIT;
  signal  \45407\    : AGCBIT;
  signal \$45407\    : AGCBIT;
  signal  \45408\    : AGCBIT;
  signal \$45408\    : AGCBIT;
  signal  \45409\    : AGCBIT;
  signal \$45409\    : AGCBIT;
  signal  \45410\    : AGCBIT;
  signal \$45410\    : AGCBIT;
  signal  \45411\    : AGCBIT;
  signal \$45411\    : AGCBIT;
  signal  \45412\    : AGCBIT;
  signal \$45412\    : AGCBIT;
  signal \&45413\    : AGCBIT;
  signal  \45414\    : AGCBIT;
  signal \$45414\    : AGCBIT;
  signal  \45415\    : AGCBIT;
  signal \$45415\    : AGCBIT;
  signal  \45416\    : AGCBIT;
  signal \$45416\    : AGCBIT;
  signal  \45417\    : AGCBIT;
  signal \$45417\    : AGCBIT;
  signal  \45418\    : AGCBIT;
  signal \$45418\    : AGCBIT;
  signal  \45419\    : AGCBIT;
  signal \$45419\    : AGCBIT;
  signal \&45420\    : AGCBIT;
  signal  \45421\    : AGCBIT;
  signal \$45421\    : AGCBIT;
  signal  \45422\    : AGCBIT;
  signal \$45422\    : AGCBIT;
  signal  \45423\    : AGCBIT;
  signal \$45423\    : AGCBIT;
  signal  \45424\    : AGCBIT;
  signal \$45424\    : AGCBIT;
  signal  \45425\    : AGCBIT;
  signal \$45425\    : AGCBIT;
  signal  \45426\    : AGCBIT;
  signal \$45426\    : AGCBIT;
  signal \&45427\    : AGCBIT;
  signal  \45428\    : AGCBIT;
  signal \$45428\    : AGCBIT;
  signal  \45429\    : AGCBIT;
  signal \$45429\    : AGCBIT;
  signal  \45430\    : AGCBIT;
  signal \$45430\    : AGCBIT;
  signal  \45431\    : AGCBIT;
  signal \$45431\    : AGCBIT;
  signal  \45432\    : AGCBIT;
  signal \$45432\    : AGCBIT;
  signal \&45433\    : AGCBIT;
  signal  \45434\    : AGCBIT; signal  \CNTOF9\   : AGCBIT;
  signal \&45435\    : AGCBIT;
  signal \&45436\    : AGCBIT;
  signal  \45437\    : AGCBIT; signal  \CH11\     : AGCBIT;
  signal \&45438\    : AGCBIT;
  signal \&45439\    : AGCBIT;
  signal  \45440\    : AGCBIT; signal  \CH12\     : AGCBIT;
  signal \&45441\    : AGCBIT;
  signal  \45442\    : AGCBIT; signal  \CH13\     : AGCBIT;
  signal \&45443\    : AGCBIT;
  signal  \45444\    : AGCBIT; signal  \CH14\     : AGCBIT;
  signal \&45445\    : AGCBIT;
  signal  \45446\    : AGCBIT; signal  \CH16\     : AGCBIT;
  signal  \45447\    : AGCBIT;
  signal  \45448\    : AGCBIT; signal  \END\      : AGCBIT;
  signal  \45449\    : AGCBIT; signal  \DLKRPT\   : AGCBIT;
  signal \$45449\    : AGCBIT;
  signal  \45450\    : AGCBIT;
  signal \$45450\    : AGCBIT;
  signal  \45451\    : AGCBIT;
  signal \$45451\    : AGCBIT;
  signal  \45452\    : AGCBIT;
  signal \$45452\    : AGCBIT;
  signal  \45453\    : AGCBIT;
  signal  \45454\    : AGCBIT;
  signal \$45454\    : AGCBIT;
  signal  \45455\    : AGCBIT;
  signal \$45455\    : AGCBIT;
  signal  \45456\    : AGCBIT; signal  \CH3312\   : AGCBIT;
  signal \&45458\    : AGCBIT;
  signal  \46101\    : AGCBIT;
  signal  \46102\    : AGCBIT; signal  \SH3MS/\   : AGCBIT;
  signal \$46102\    : AGCBIT;
  signal  \46103\    : AGCBIT;
  signal \$46103\    : AGCBIT;
  signal  \46104\    : AGCBIT;
  signal  \46105\    : AGCBIT;
  signal  \46106\    : AGCBIT;
  signal  \46107\    : AGCBIT;
  signal  \46108\    : AGCBIT;
  signal  \46109\    : AGCBIT; signal  \ALT0\     : AGCBIT;
  signal  \46110\    : AGCBIT; signal  \ALT1\     : AGCBIT;
  signal  \46111\    : AGCBIT; signal  \ALRT0\    : AGCBIT;
  signal  \46112\    : AGCBIT; signal  \ALRT1\    : AGCBIT;
  signal  \46113\    : AGCBIT;
  signal  \46114\    : AGCBIT;
  signal \$46114\    : AGCBIT;
  signal  \46115\    : AGCBIT;
  signal \$46115\    : AGCBIT;
  signal  \46116\    : AGCBIT; signal  \CH1402\   : AGCBIT;
  signal  \46117\    : AGCBIT;
  signal  \46118\    : AGCBIT;
  signal \$46118\    : AGCBIT;
  signal  \46119\    : AGCBIT;
  signal \$46119\    : AGCBIT;
  signal  \46120\    : AGCBIT; signal  \CH1403\   : AGCBIT;
  signal  \46121\    : AGCBIT;
  signal  \46122\    : AGCBIT;
  signal  \46123\    : AGCBIT;
  signal  \46124\    : AGCBIT;
  signal \$46124\    : AGCBIT;
  signal  \46125\    : AGCBIT;
  signal \$46125\    : AGCBIT;
  signal  \46126\    : AGCBIT;
  signal  \46127\    : AGCBIT;
  signal \$46127\    : AGCBIT;
  signal  \46128\    : AGCBIT;
  signal \$46128\    : AGCBIT;
  signal  \46129\    : AGCBIT; signal  \ALTM\     : AGCBIT;
  signal  \46130\    : AGCBIT;
  signal \$46130\    : AGCBIT;
  signal  \46131\    : AGCBIT;
  signal \$46131\    : AGCBIT;
  signal  \46132\    : AGCBIT; signal  \ALTSNC\   : AGCBIT;
  signal  \46133\    : AGCBIT;
  signal  \46134\    : AGCBIT;
  signal  \46135\    : AGCBIT;
  signal \$46135\    : AGCBIT;
  signal  \46136\    : AGCBIT;
  signal \$46136\    : AGCBIT;
  signal  \46137\    : AGCBIT;
  signal  \46138\    : AGCBIT;
  signal \$46138\    : AGCBIT;
  signal  \46139\    : AGCBIT;
  signal \$46139\    : AGCBIT;
  signal  \46140\    : AGCBIT;
  signal  \46141\    : AGCBIT;
  signal \$46141\    : AGCBIT;
  signal  \46142\    : AGCBIT;
  signal \$46142\    : AGCBIT;
  signal  \46143\    : AGCBIT; signal  \OTLNKM\   : AGCBIT;
  signal  \46144\    : AGCBIT;
  signal  \46145\    : AGCBIT; signal  \CH1401\   : AGCBIT;
  signal  \46146\    : AGCBIT;
  signal  \46147\    : AGCBIT; signal  \OTLNK0\   : AGCBIT;
  signal  \46148\    : AGCBIT;
  signal  \46149\    : AGCBIT; signal  \OTLNK1\   : AGCBIT;
  signal  \46150\    : AGCBIT;
  signal  \46151\    : AGCBIT;
  signal  \46152\    : AGCBIT; signal  \F5ASB0\   : AGCBIT;
  signal  \46153\    : AGCBIT; signal  \F5ASB0/\  : AGCBIT;
  signal  \46154\    : AGCBIT; signal  \F5ASB2\   : AGCBIT;
  signal  \46155\    : AGCBIT; signal  \F5ASB2/\  : AGCBIT;
  signal  \46156\    : AGCBIT; signal  \F5BSB2\   : AGCBIT;
  signal  \46157\    : AGCBIT; signal  \F5BSB2/\  : AGCBIT;
  signal  \46158\    : AGCBIT;
  signal  \46159\    : AGCBIT;
  signal  \46160\    : AGCBIT; signal  \T2P\      : AGCBIT;
  signal  \46201\    : AGCBIT;
  signal  \46202\    : AGCBIT;
  signal  \46203\    : AGCBIT; signal  \INLNKM\   : AGCBIT;
  signal  \46204\    : AGCBIT;
  signal  \46205\    : AGCBIT;
  signal  \46206\    : AGCBIT; signal  \INLNKP\   : AGCBIT;
  signal  \46207\    : AGCBIT;
  signal  \46208\    : AGCBIT;
  signal \&46209\    : AGCBIT;
  signal  \46210\    : AGCBIT;
  signal  \46211\    : AGCBIT;
  signal  \46212\    : AGCBIT; signal  \CCH33\    : AGCBIT;
  signal  \46213\    : AGCBIT;
  signal \$46213\    : AGCBIT;
  signal  \46214\    : AGCBIT;
  signal \$46214\    : AGCBIT;
  signal  \46215\    : AGCBIT; signal  \CH3311\   : AGCBIT;
  signal  \46216\    : AGCBIT;
  signal \$46216\    : AGCBIT;
  signal  \46217\    : AGCBIT;
  signal \$46217\    : AGCBIT;
  signal  \46218\    : AGCBIT;
  signal \$46218\    : AGCBIT;
  signal  \46219\    : AGCBIT;
  signal \$46219\    : AGCBIT;
  signal  \46220\    : AGCBIT; signal  \C45R/\    : AGCBIT;
  signal  \46221\    : AGCBIT; signal  \CH3310\   : AGCBIT;
  signal  \46222\    : AGCBIT;
  signal  \46223\    : AGCBIT;
  signal  \46224\    : AGCBIT;
  signal \$46224\    : AGCBIT;
  signal  \46225\    : AGCBIT;
  signal \$46225\    : AGCBIT;
  signal  \46226\    : AGCBIT;
  signal \$46226\    : AGCBIT;
  signal  \46227\    : AGCBIT;
  signal \$46227\    : AGCBIT;
  signal  \46228\    : AGCBIT; signal  \CH1305\   : AGCBIT;
  signal  \46229\    : AGCBIT; signal  \CH1306\   : AGCBIT;
  signal  \46230\    : AGCBIT;
  signal  \46231\    : AGCBIT;
  signal \$46231\    : AGCBIT;
  signal  \46232\    : AGCBIT;
  signal \$46232\    : AGCBIT;
  signal  \46233\    : AGCBIT; signal  \CH1404\   : AGCBIT;
  signal  \46234\    : AGCBIT; signal  \THRSTD\   : AGCBIT;
  signal  \46235\    : AGCBIT;
  signal  \46236\    : AGCBIT;
  signal \$46236\    : AGCBIT;
  signal  \46237\    : AGCBIT;
  signal \$46237\    : AGCBIT;
  signal  \46238\    : AGCBIT; signal  \CH1405\   : AGCBIT;
  signal  \46239\    : AGCBIT; signal  \EMSD\     : AGCBIT;
  signal  \46240\    : AGCBIT;
  signal  \46241\    : AGCBIT;
  signal  \46242\    : AGCBIT;
  signal  \46243\    : AGCBIT;
  signal \$46243\    : AGCBIT;
  signal  \46244\    : AGCBIT;
  signal \$46244\    : AGCBIT;
  signal  \46245\    : AGCBIT;
  signal \$46245\    : AGCBIT;
  signal  \46246\    : AGCBIT;
  signal \$46246\    : AGCBIT;
  signal  \46247\    : AGCBIT; signal  \THRST+\   : AGCBIT;
  signal  \46248\    : AGCBIT; signal  \THRST-\   : AGCBIT;
  signal  \46249\    : AGCBIT;
  signal  \46250\    : AGCBIT;
  signal  \46251\    : AGCBIT;
  signal  \46252\    : AGCBIT;
  signal \$46252\    : AGCBIT;
  signal  \46253\    : AGCBIT;
  signal \$46253\    : AGCBIT;
  signal  \46254\    : AGCBIT; signal  \EMS+\     : AGCBIT;
  signal  \46255\    : AGCBIT;
  signal  \46256\    : AGCBIT;
  signal \$46256\    : AGCBIT;
  signal  \46257\    : AGCBIT;
  signal \$46257\    : AGCBIT;
  signal  \46258\    : AGCBIT; signal  \EMS-\     : AGCBIT;
  signal  \46259\    : AGCBIT;
  signal \&46261\    : AGCBIT;
  signal  \46303\    : AGCBIT; signal  \UPRUPT\   : AGCBIT;
  signal  \46304\    : AGCBIT; signal  \UPL0/\    : AGCBIT;
  signal  \46305\    : AGCBIT; signal  \UPL1/\    : AGCBIT;
  signal  \46306\    : AGCBIT; signal  \XLNK0/\   : AGCBIT;
  signal  \46307\    : AGCBIT; signal  \XLNK1/\   : AGCBIT;
  signal  \46308\    : AGCBIT; signal  \BLKUPL\   : AGCBIT;
  signal  \46309\    : AGCBIT; signal  \F10B/\    : AGCBIT;
  signal  \46310\    : AGCBIT; signal  \T1P\      : AGCBIT;
  signal  \46311\    : AGCBIT; signal  \T3P\      : AGCBIT;
  signal  \46312\    : AGCBIT; signal  \F09B/\    : AGCBIT;
  signal  \46313\    : AGCBIT; signal  \T4P\      : AGCBIT;
  signal  \46314\    : AGCBIT; signal  \F10A/\    : AGCBIT;
  signal  \46315\    : AGCBIT; signal  \T5P\      : AGCBIT;
  signal  \46316\    : AGCBIT; signal  \F06B/\    : AGCBIT;
  signal  \46317\    : AGCBIT; signal  \T6P\      : AGCBIT;
  signal  \46318\    : AGCBIT;
  signal  \46319\    : AGCBIT;
  signal \$46319\    : AGCBIT;
  signal  \46320\    : AGCBIT;
  signal \$46320\    : AGCBIT;
  signal  \46321\    : AGCBIT; signal  \CH1308\   : AGCBIT;
  signal  \46322\    : AGCBIT;
  signal  \46323\    : AGCBIT;
  signal  \46324\    : AGCBIT;
  signal \$46324\    : AGCBIT;
  signal  \46325\    : AGCBIT;
  signal \$46325\    : AGCBIT;
  signal  \46326\    : AGCBIT; signal  \CH1309\   : AGCBIT;
  signal  \46327\    : AGCBIT;
  signal  \46328\    : AGCBIT;
  signal \$46328\    : AGCBIT;
  signal  \46329\    : AGCBIT;
  signal \$46329\    : AGCBIT;
  signal  \46330\    : AGCBIT; signal  \RHCGO\    : AGCBIT;
  signal  \46331\    : AGCBIT;
  signal  \46332\    : AGCBIT;
  signal  \46333\    : AGCBIT;
  signal \$46333\    : AGCBIT;
  signal  \46334\    : AGCBIT;
  signal \$46334\    : AGCBIT;
  signal  \46335\    : AGCBIT;
  signal  \46336\    : AGCBIT;
  signal  \46337\    : AGCBIT;
  signal  \46338\    : AGCBIT;
  signal  \46339\    : AGCBIT; signal  \BMAGXP\   : AGCBIT;
  signal  \46340\    : AGCBIT; signal  \BMAGXM\   : AGCBIT;
  signal  \46341\    : AGCBIT;
  signal  \46342\    : AGCBIT;
  signal \$46342\    : AGCBIT;
  signal  \46343\    : AGCBIT;
  signal \$46343\    : AGCBIT;
  signal  \46344\    : AGCBIT;
  signal  \46345\    : AGCBIT;
  signal  \46346\    : AGCBIT;
  signal  \46347\    : AGCBIT;
  signal  \46348\    : AGCBIT; signal  \BMAGYP\   : AGCBIT;
  signal  \46349\    : AGCBIT; signal  \BMAGYM\   : AGCBIT;
  signal  \46350\    : AGCBIT;
  signal  \46351\    : AGCBIT;
  signal  \46352\    : AGCBIT;
  signal \$46352\    : AGCBIT;
  signal  \46353\    : AGCBIT;
  signal \$46353\    : AGCBIT;
  signal  \46354\    : AGCBIT;
  signal  \46355\    : AGCBIT;
  signal  \46356\    : AGCBIT;
  signal  \46357\    : AGCBIT;
  signal  \46358\    : AGCBIT; signal  \BMAGZP\   : AGCBIT;
  signal  \46359\    : AGCBIT; signal  \BMAGZM\   : AGCBIT;
  signal  \46401\    : AGCBIT;
  signal  \46402\    : AGCBIT;
  signal \$46402\    : AGCBIT;
  signal  \46403\    : AGCBIT;
  signal \$46403\    : AGCBIT;
  signal  \46404\    : AGCBIT; signal  \CH1410\   : AGCBIT;
  signal  \46405\    : AGCBIT; signal  \GYROD\    : AGCBIT;
  signal  \46406\    : AGCBIT;
  signal  \46407\    : AGCBIT;
  signal \$46407\    : AGCBIT;
  signal  \46408\    : AGCBIT;
  signal \$46408\    : AGCBIT;
  signal  \46409\    : AGCBIT; signal  \CH1409\   : AGCBIT;
  signal  \46410\    : AGCBIT;
  signal  \46411\    : AGCBIT;
  signal \$46411\    : AGCBIT;
  signal  \46412\    : AGCBIT;
  signal \$46412\    : AGCBIT;
  signal  \46413\    : AGCBIT; signal  \CH1408\   : AGCBIT;
  signal  \46414\    : AGCBIT;
  signal  \46415\    : AGCBIT;
  signal \$46415\    : AGCBIT;
  signal  \46416\    : AGCBIT;
  signal \$46416\    : AGCBIT;
  signal  \46417\    : AGCBIT; signal  \CH1407\   : AGCBIT;
  signal  \46418\    : AGCBIT;
  signal  \46419\    : AGCBIT;
  signal \$46419\    : AGCBIT;
  signal  \46420\    : AGCBIT;
  signal \$46420\    : AGCBIT;
  signal  \46421\    : AGCBIT; signal  \CH1406\   : AGCBIT;
  signal  \46422\    : AGCBIT;
  signal  \46423\    : AGCBIT;
  signal  \46424\    : AGCBIT; signal  \GYXP\     : AGCBIT;
  signal  \46425\    : AGCBIT; signal  \GYXM\     : AGCBIT;
  signal  \46426\    : AGCBIT; signal  \GYYP\     : AGCBIT;
  signal  \46427\    : AGCBIT; signal  \GYYM\     : AGCBIT;
  signal  \46428\    : AGCBIT;
  signal  \46429\    : AGCBIT;
  signal  \46430\    : AGCBIT;
  signal  \46431\    : AGCBIT;
  signal  \46432\    : AGCBIT; signal  \GYZP\     : AGCBIT;
  signal  \46433\    : AGCBIT; signal  \GYZM\     : AGCBIT;
  signal  \46434\    : AGCBIT; signal  \GYENAB\   : AGCBIT;
  signal  \46435\    : AGCBIT;
  signal  \46436\    : AGCBIT;
  signal  \46437\    : AGCBIT;
  signal  \46438\    : AGCBIT;
  signal  \46439\    : AGCBIT;
  signal  \46440\    : AGCBIT;
  signal \$46440\    : AGCBIT;
  signal  \46441\    : AGCBIT;
  signal \$46441\    : AGCBIT;
  signal  \46442\    : AGCBIT; signal  \GYRSET\   : AGCBIT;
  signal  \46443\    : AGCBIT; signal  \GYRRST\   : AGCBIT;
  signal  \46444\    : AGCBIT;
  signal  \46445\    : AGCBIT; signal  \FF1109/\  : AGCBIT;
  signal \$46445\    : AGCBIT;
  signal  \46446\    : AGCBIT; signal  \FF1109\   : AGCBIT;
  signal \$46446\    : AGCBIT;
  signal  \46447\    : AGCBIT; signal  \CH1109\   : AGCBIT;
  signal  \46448\    : AGCBIT; signal  \W1110\    : AGCBIT;
  signal  \46449\    : AGCBIT; signal  \FF1110/\  : AGCBIT;
  signal \$46449\    : AGCBIT;
  signal  \46450\    : AGCBIT; signal  \FF1110\   : AGCBIT;
  signal \$46450\    : AGCBIT;
  signal  \46451\    : AGCBIT; signal  \CH1110\   : AGCBIT;
  signal  \46452\    : AGCBIT;
  signal  \46453\    : AGCBIT; signal  \FF1111/\  : AGCBIT;
  signal \$46453\    : AGCBIT;
  signal  \46454\    : AGCBIT; signal  \FF1111\   : AGCBIT;
  signal \$46454\    : AGCBIT;
  signal  \46455\    : AGCBIT; signal  \CH1111\   : AGCBIT;
  signal  \46456\    : AGCBIT;
  signal  \46457\    : AGCBIT; signal  \FF1112/\  : AGCBIT;
  signal \$46457\    : AGCBIT;
  signal  \46458\    : AGCBIT; signal  \FF1112\   : AGCBIT;
  signal \$46458\    : AGCBIT;
  signal  \46459\    : AGCBIT; signal  \CH1112\   : AGCBIT;
  signal  \31101\    : AGCBIT;
  signal  \31102\    : AGCBIT;
  signal \$31102\    : AGCBIT;
  signal  \31103\    : AGCBIT;
  signal \$31103\    : AGCBIT;
  signal  \31104\    : AGCBIT;
  signal  \31105\    : AGCBIT;
  signal  \31106\    : AGCBIT;
  signal \$31106\    : AGCBIT;
  signal  \31107\    : AGCBIT;
  signal \$31107\    : AGCBIT;
  signal  \31108\    : AGCBIT; signal  \C32A\     : AGCBIT;
  signal  \31109\    : AGCBIT;
  signal \$31109\    : AGCBIT;
  signal  \31110\    : AGCBIT;
  signal \$31110\    : AGCBIT;
  signal  \31111\    : AGCBIT;
  signal  \31112\    : AGCBIT; signal  \C32R\     : AGCBIT;
  signal  \31113\    : AGCBIT; signal  \C32P\     : AGCBIT;
  signal  \31114\    : AGCBIT; signal  \C32M\     : AGCBIT;
  signal  \31115\    : AGCBIT;
  signal \$31115\    : AGCBIT;
  signal  \31116\    : AGCBIT;
  signal \$31116\    : AGCBIT;
  signal  \31117\    : AGCBIT;
  signal  \31118\    : AGCBIT;
  signal  \31119\    : AGCBIT;
  signal \$31119\    : AGCBIT;
  signal  \31120\    : AGCBIT;
  signal \$31120\    : AGCBIT;
  signal  \31121\    : AGCBIT; signal  \C33A\     : AGCBIT;
  signal  \31122\    : AGCBIT;
  signal  \31123\    : AGCBIT; signal  \CG11\     : AGCBIT;
  signal  \31124\    : AGCBIT;
  signal \$31124\    : AGCBIT;
  signal  \31125\    : AGCBIT;
  signal \$31125\    : AGCBIT;
  signal  \31126\    : AGCBIT; signal  \C33R\     : AGCBIT;
  signal  \31127\    : AGCBIT; signal  \C33P\     : AGCBIT;
  signal  \31128\    : AGCBIT; signal  \C33M\     : AGCBIT;
  signal  \31129\    : AGCBIT;
  signal \$31129\    : AGCBIT;
  signal  \31130\    : AGCBIT;
  signal \$31130\    : AGCBIT;
  signal  \31131\    : AGCBIT;
  signal  \31132\    : AGCBIT;
  signal \$31132\    : AGCBIT;
  signal  \31133\    : AGCBIT;
  signal \$31133\    : AGCBIT;
  signal  \31134\    : AGCBIT; signal  \C24A\     : AGCBIT;
  signal  \31135\    : AGCBIT; signal  \C24R\     : AGCBIT;
  signal  \31136\    : AGCBIT;
  signal \$31136\    : AGCBIT;
  signal  \31137\    : AGCBIT;
  signal \$31137\    : AGCBIT;
  signal  \31138\    : AGCBIT;
  signal  \31139\    : AGCBIT;
  signal \$31139\    : AGCBIT;
  signal  \31140\    : AGCBIT;
  signal \$31140\    : AGCBIT;
  signal  \31141\    : AGCBIT; signal  \C25A\     : AGCBIT;
  signal  \31142\    : AGCBIT; signal  \C25R\     : AGCBIT;
  signal  \31143\    : AGCBIT;
  signal \$31143\    : AGCBIT;
  signal  \31144\    : AGCBIT;
  signal \$31144\    : AGCBIT;
  signal  \31145\    : AGCBIT;
  signal  \31146\    : AGCBIT;
  signal \$31146\    : AGCBIT;
  signal  \31147\    : AGCBIT;
  signal \$31147\    : AGCBIT;
  signal \&31148\    : AGCBIT;
  signal  \31149\    : AGCBIT; signal  \C26A\     : AGCBIT;
  signal  \31150\    : AGCBIT;
  signal \&31151\    : AGCBIT;
  signal  \31152\    : AGCBIT; signal  \CG21\     : AGCBIT;
  signal  \31153\    : AGCBIT; signal  \C26R\     : AGCBIT;
  signal  \31154\    : AGCBIT; signal  \CA3/\     : AGCBIT;
  signal  \31158\    : AGCBIT; signal  \CXB7/\    : AGCBIT;
  signal  \31201\    : AGCBIT;
  signal  \31202\    : AGCBIT;
  signal \$31202\    : AGCBIT;
  signal  \31203\    : AGCBIT;
  signal \$31203\    : AGCBIT;
  signal  \31204\    : AGCBIT;
  signal  \31205\    : AGCBIT;
  signal  \31206\    : AGCBIT;
  signal \$31206\    : AGCBIT;
  signal  \31207\    : AGCBIT;
  signal \$31207\    : AGCBIT;
  signal  \31208\    : AGCBIT; signal  \C34A\     : AGCBIT;
  signal  \31209\    : AGCBIT;
  signal \$31209\    : AGCBIT;
  signal  \31210\    : AGCBIT;
  signal \$31210\    : AGCBIT;
  signal  \31211\    : AGCBIT;
  signal  \31212\    : AGCBIT; signal  \C34R\     : AGCBIT;
  signal  \31213\    : AGCBIT; signal  \C34P\     : AGCBIT;
  signal  \31214\    : AGCBIT; signal  \C34M\     : AGCBIT;
  signal  \31215\    : AGCBIT;
  signal \$31215\    : AGCBIT;
  signal  \31216\    : AGCBIT;
  signal \$31216\    : AGCBIT;
  signal  \31217\    : AGCBIT;
  signal  \31218\    : AGCBIT;
  signal  \31219\    : AGCBIT;
  signal \$31219\    : AGCBIT;
  signal  \31220\    : AGCBIT;
  signal \$31220\    : AGCBIT;
  signal  \31221\    : AGCBIT; signal  \C35A\     : AGCBIT;
  signal  \31222\    : AGCBIT;
  signal  \31223\    : AGCBIT; signal  \CG12\     : AGCBIT;
  signal  \31224\    : AGCBIT;
  signal \$31224\    : AGCBIT;
  signal  \31225\    : AGCBIT;
  signal \$31225\    : AGCBIT;
  signal  \31226\    : AGCBIT; signal  \C35R\     : AGCBIT;
  signal  \31227\    : AGCBIT; signal  \C35P\     : AGCBIT;
  signal  \31228\    : AGCBIT; signal  \C35M\     : AGCBIT;
  signal  \31229\    : AGCBIT;
  signal \$31229\    : AGCBIT;
  signal  \31230\    : AGCBIT;
  signal \$31230\    : AGCBIT;
  signal  \31231\    : AGCBIT;
  signal  \31232\    : AGCBIT;
  signal \$31232\    : AGCBIT;
  signal  \31233\    : AGCBIT;
  signal \$31233\    : AGCBIT;
  signal  \31234\    : AGCBIT; signal  \C27A\     : AGCBIT;
  signal  \31235\    : AGCBIT; signal  \C27R\     : AGCBIT;
  signal  \31236\    : AGCBIT;
  signal \$31236\    : AGCBIT;
  signal  \31237\    : AGCBIT;
  signal \$31237\    : AGCBIT;
  signal  \31238\    : AGCBIT;
  signal  \31239\    : AGCBIT;
  signal \$31239\    : AGCBIT;
  signal  \31240\    : AGCBIT;
  signal \$31240\    : AGCBIT;
  signal  \31241\    : AGCBIT; signal  \C30A\     : AGCBIT;
  signal  \31242\    : AGCBIT; signal  \C30R\     : AGCBIT;
  signal  \31243\    : AGCBIT;
  signal \$31243\    : AGCBIT;
  signal  \31244\    : AGCBIT;
  signal \$31244\    : AGCBIT;
  signal  \31245\    : AGCBIT;
  signal  \31246\    : AGCBIT;
  signal \$31246\    : AGCBIT;
  signal  \31247\    : AGCBIT;
  signal \$31247\    : AGCBIT;
  signal \&31248\    : AGCBIT;
  signal  \31249\    : AGCBIT; signal  \C31A\     : AGCBIT;
  signal  \31250\    : AGCBIT;
  signal \&31251\    : AGCBIT;
  signal  \31252\    : AGCBIT; signal  \CG22\     : AGCBIT;
  signal  \31253\    : AGCBIT; signal  \C31R\     : AGCBIT;
  signal  \31256\    : AGCBIT; signal  \CXB2/\    : AGCBIT;
  signal  \31301\    : AGCBIT;
  signal  \31302\    : AGCBIT;
  signal \$31302\    : AGCBIT;
  signal  \31303\    : AGCBIT;
  signal \$31303\    : AGCBIT;
  signal  \31304\    : AGCBIT;
  signal  \31305\    : AGCBIT;
  signal  \31306\    : AGCBIT;
  signal \$31306\    : AGCBIT;
  signal  \31307\    : AGCBIT;
  signal \$31307\    : AGCBIT;
  signal  \31308\    : AGCBIT; signal  \C36A\     : AGCBIT;
  signal  \31309\    : AGCBIT;
  signal \$31309\    : AGCBIT;
  signal  \31310\    : AGCBIT;
  signal \$31310\    : AGCBIT;
  signal  \31311\    : AGCBIT;
  signal  \31312\    : AGCBIT; signal  \C36R\     : AGCBIT;
  signal  \31313\    : AGCBIT; signal  \C36P\     : AGCBIT;
  signal  \31314\    : AGCBIT; signal  \C36M\     : AGCBIT;
  signal  \31315\    : AGCBIT;
  signal \$31315\    : AGCBIT;
  signal  \31316\    : AGCBIT;
  signal \$31316\    : AGCBIT;
  signal  \31317\    : AGCBIT;
  signal  \31318\    : AGCBIT;
  signal  \31319\    : AGCBIT;
  signal \$31319\    : AGCBIT;
  signal  \31320\    : AGCBIT;
  signal \$31320\    : AGCBIT;
  signal  \31321\    : AGCBIT; signal  \C37A\     : AGCBIT;
  signal  \31322\    : AGCBIT;
  signal  \31323\    : AGCBIT; signal  \CG14\     : AGCBIT;
  signal  \31324\    : AGCBIT;
  signal \$31324\    : AGCBIT;
  signal  \31325\    : AGCBIT;
  signal \$31325\    : AGCBIT;
  signal  \31326\    : AGCBIT; signal  \C37R\     : AGCBIT;
  signal  \31327\    : AGCBIT; signal  \C37P\     : AGCBIT;
  signal  \31328\    : AGCBIT; signal  \C37M\     : AGCBIT;
  signal  \31329\    : AGCBIT;
  signal \$31329\    : AGCBIT;
  signal  \31330\    : AGCBIT;
  signal \$31330\    : AGCBIT;
  signal  \31331\    : AGCBIT;
  signal  \31332\    : AGCBIT;
  signal \$31332\    : AGCBIT;
  signal  \31333\    : AGCBIT;
  signal \$31333\    : AGCBIT;
  signal  \31334\    : AGCBIT; signal  \C50A\     : AGCBIT;
  signal  \31335\    : AGCBIT; signal  \C50R\     : AGCBIT;
  signal  \31336\    : AGCBIT;
  signal \$31336\    : AGCBIT;
  signal  \31337\    : AGCBIT;
  signal \$31337\    : AGCBIT;
  signal  \31338\    : AGCBIT;
  signal  \31339\    : AGCBIT;
  signal \$31339\    : AGCBIT;
  signal  \31340\    : AGCBIT;
  signal \$31340\    : AGCBIT;
  signal  \31341\    : AGCBIT; signal  \C51A\     : AGCBIT;
  signal  \31342\    : AGCBIT; signal  \C51R\     : AGCBIT;
  signal  \31343\    : AGCBIT;
  signal \$31343\    : AGCBIT;
  signal  \31344\    : AGCBIT;
  signal \$31344\    : AGCBIT;
  signal  \31345\    : AGCBIT;
  signal  \31346\    : AGCBIT;
  signal \$31346\    : AGCBIT;
  signal  \31347\    : AGCBIT;
  signal \$31347\    : AGCBIT;
  signal \&31348\    : AGCBIT;
  signal  \31349\    : AGCBIT; signal  \C52A\     : AGCBIT;
  signal  \31350\    : AGCBIT;
  signal \&31351\    : AGCBIT;
  signal  \31352\    : AGCBIT; signal  \CG24\     : AGCBIT;
  signal  \31353\    : AGCBIT; signal  \C52R\     : AGCBIT;
  signal  \31354\    : AGCBIT; signal  \CA4/\     : AGCBIT;
  signal  \31356\    : AGCBIT; signal  \CXB3/\    : AGCBIT;
  signal  \31358\    : AGCBIT; signal  \CA2/\     : AGCBIT;
  signal  \31401\    : AGCBIT;
  signal  \31402\    : AGCBIT;
  signal \$31402\    : AGCBIT;
  signal  \31403\    : AGCBIT;
  signal \$31403\    : AGCBIT;
  signal  \31404\    : AGCBIT;
  signal  \31405\    : AGCBIT;
  signal  \31406\    : AGCBIT;
  signal \$31406\    : AGCBIT;
  signal  \31407\    : AGCBIT;
  signal \$31407\    : AGCBIT;
  signal  \31408\    : AGCBIT; signal  \C40A\     : AGCBIT;
  signal  \31409\    : AGCBIT;
  signal \$31409\    : AGCBIT;
  signal  \31410\    : AGCBIT;
  signal \$31410\    : AGCBIT;
  signal  \31411\    : AGCBIT;
  signal  \31412\    : AGCBIT; signal  \C40R\     : AGCBIT;
  signal  \31413\    : AGCBIT; signal  \C40P\     : AGCBIT;
  signal  \31414\    : AGCBIT; signal  \C40M\     : AGCBIT;
  signal  \31415\    : AGCBIT;
  signal \$31415\    : AGCBIT;
  signal  \31416\    : AGCBIT;
  signal \$31416\    : AGCBIT;
  signal  \31417\    : AGCBIT;
  signal  \31418\    : AGCBIT;
  signal  \31419\    : AGCBIT;
  signal \$31419\    : AGCBIT;
  signal  \31420\    : AGCBIT;
  signal \$31420\    : AGCBIT;
  signal  \31421\    : AGCBIT; signal  \C41A\     : AGCBIT;
  signal  \31422\    : AGCBIT;
  signal  \31423\    : AGCBIT; signal  \CG13\     : AGCBIT;
  signal  \31424\    : AGCBIT;
  signal \$31424\    : AGCBIT;
  signal  \31425\    : AGCBIT;
  signal \$31425\    : AGCBIT;
  signal  \31426\    : AGCBIT; signal  \C41R\     : AGCBIT;
  signal  \31427\    : AGCBIT; signal  \C41P\     : AGCBIT;
  signal  \31428\    : AGCBIT; signal  \C41M\     : AGCBIT;
  signal  \31429\    : AGCBIT;
  signal \$31429\    : AGCBIT;
  signal  \31430\    : AGCBIT;
  signal \$31430\    : AGCBIT;
  signal  \31431\    : AGCBIT;
  signal  \31432\    : AGCBIT;
  signal \$31432\    : AGCBIT;
  signal  \31433\    : AGCBIT;
  signal \$31433\    : AGCBIT;
  signal  \31434\    : AGCBIT; signal  \C53A\     : AGCBIT;
  signal  \31435\    : AGCBIT; signal  \C53R\     : AGCBIT;
  signal  \31436\    : AGCBIT;
  signal \$31436\    : AGCBIT;
  signal  \31437\    : AGCBIT;
  signal \$31437\    : AGCBIT;
  signal  \31438\    : AGCBIT;
  signal  \31439\    : AGCBIT;
  signal \$31439\    : AGCBIT;
  signal  \31440\    : AGCBIT;
  signal \$31440\    : AGCBIT;
  signal  \31441\    : AGCBIT; signal  \C54A\     : AGCBIT;
  signal  \31442\    : AGCBIT; signal  \C54R\     : AGCBIT;
  signal  \31443\    : AGCBIT;
  signal \$31443\    : AGCBIT;
  signal  \31444\    : AGCBIT;
  signal \$31444\    : AGCBIT;
  signal  \31445\    : AGCBIT;
  signal  \31446\    : AGCBIT;
  signal \$31446\    : AGCBIT;
  signal  \31447\    : AGCBIT;
  signal \$31447\    : AGCBIT;
  signal \&31448\    : AGCBIT;
  signal  \31449\    : AGCBIT; signal  \C55A\     : AGCBIT;
  signal  \31450\    : AGCBIT;
  signal \&31451\    : AGCBIT;
  signal  \31452\    : AGCBIT; signal  \CG23\     : AGCBIT;
  signal  \31453\    : AGCBIT; signal  \C55R\     : AGCBIT;
  signal  \31456\    : AGCBIT; signal  \CXB4/\    : AGCBIT;
  signal  \31458\    : AGCBIT; signal  \CA6/\     : AGCBIT;
  signal \&32001\    : AGCBIT;
  signal \&32002\    : AGCBIT;
  signal \&32003\    : AGCBIT;
  signal \&32004\    : AGCBIT;
  signal \&32005\    : AGCBIT;
  signal \&32006\    : AGCBIT;
  signal  \32007\    : AGCBIT;
  signal  \32008\    : AGCBIT; signal  \CAD4\     : AGCBIT;
  signal \&32011\    : AGCBIT;
  signal \&32012\    : AGCBIT;
  signal \&32013\    : AGCBIT;
  signal  \32014\    : AGCBIT; signal  \32004K?\  : AGCBIT;
  signal  \32015\    : AGCBIT;
  signal  \32016\    : AGCBIT;
  signal  \32021\    : AGCBIT;
  signal  \32022\    : AGCBIT;
  signal \&32023\    : AGCBIT;
  signal \&32024\    : AGCBIT;
  signal \&32026\    : AGCBIT;
  signal \&32031\    : AGCBIT;
  signal \&32032\    : AGCBIT;
  signal  \32033\    : AGCBIT;
  signal \&32034\    : AGCBIT;
  signal  \32035\    : AGCBIT; signal  \CAD5\     : AGCBIT;
  signal \&32036\    : AGCBIT;
  signal \&32041\    : AGCBIT;
  signal \&32042\    : AGCBIT;
  signal \&32043\    : AGCBIT;
  signal  \32044\    : AGCBIT;
  signal  \32045\    : AGCBIT; signal  \DINC/\    : AGCBIT;
  signal  \32046\    : AGCBIT; signal  \CAD6\     : AGCBIT;
  signal  \32047\    : AGCBIT; signal  \DINC\     : AGCBIT;
  signal  \32048\    : AGCBIT; signal  \DINCNC/\  : AGCBIT;
  signal \$32048\    : AGCBIT;
  signal  \32049\    : AGCBIT;
  signal  \32050\    : AGCBIT; signal  \50SUM\    : AGCBIT;
  signal  \32051\    : AGCBIT; signal  \CAD1\     : AGCBIT;
  signal  \32052\    : AGCBIT; signal  \CAD2\     : AGCBIT;
  signal \&32053\    : AGCBIT;
  signal \&32054\    : AGCBIT;
  signal \&32055\    : AGCBIT;
  signal  \32056\    : AGCBIT;
  signal  \32058\    : AGCBIT;
  signal  \32059\    : AGCBIT; signal  \SHINC/\   : AGCBIT;
  signal \$32059\    : AGCBIT;
  signal  \32060\    : AGCBIT; signal  \SHINC\    : AGCBIT;
  signal  \32061\    : AGCBIT;
  signal  \32062\    : AGCBIT;
  signal  \32063\    : AGCBIT; signal  \CAD3\     : AGCBIT;
  signal  \32064\    : AGCBIT; signal  \30SUM\    : AGCBIT;
  signal  \32065\    : AGCBIT; signal  \SHANC/\   : AGCBIT;
  signal \$32065\    : AGCBIT;
  signal  \32066\    : AGCBIT; signal  \SHANC\    : AGCBIT;
  signal \&32067\    : AGCBIT;
  signal  \32068\    : AGCBIT;
  signal \&32069\    : AGCBIT;
  signal \&32201\    : AGCBIT;
  signal  \32202\    : AGCBIT;
  signal  \32203\    : AGCBIT;
  signal  \32204\    : AGCBIT;
  signal  \32205\    : AGCBIT;
  signal  \32206\    : AGCBIT;
  signal \$32206\    : AGCBIT;
  signal  \32207\    : AGCBIT;
  signal \$32207\    : AGCBIT;
  signal  \32208\    : AGCBIT; signal  \STORE1\   : AGCBIT;
  signal  \32209\    : AGCBIT; signal  \STORE1/\  : AGCBIT;
  signal  \32210\    : AGCBIT; signal  \STFET1/\  : AGCBIT;
  signal  \32211\    : AGCBIT;
  signal  \32212\    : AGCBIT;
  signal  \32213\    : AGCBIT;
  signal \$32213\    : AGCBIT;
  signal  \32214\    : AGCBIT;
  signal \$32214\    : AGCBIT;
  signal  \32215\    : AGCBIT; signal  \MON/\     : AGCBIT;
  signal  \32216\    : AGCBIT; signal  \FETCH1\   : AGCBIT;
  signal  \32217\    : AGCBIT; signal  \FETCH0\   : AGCBIT;
  signal  \32218\    : AGCBIT;
  signal  \32219\    : AGCBIT; signal  \FETCH0/\  : AGCBIT;
  signal  \32220\    : AGCBIT;
  signal  \32221\    : AGCBIT;
  signal  \32222\    : AGCBIT;
  signal \$32222\    : AGCBIT;
  signal  \32223\    : AGCBIT; signal  \INOTLD\   : AGCBIT;
  signal \$32223\    : AGCBIT;
  signal  \32224\    : AGCBIT;
  signal  \32225\    : AGCBIT;
  signal  \32226\    : AGCBIT;
  signal \$32226\    : AGCBIT;
  signal  \32227\    : AGCBIT; signal  \INOTRD\   : AGCBIT;
  signal \$32227\    : AGCBIT;
  signal  \32228\    : AGCBIT;
  signal \&32229\    : AGCBIT;
  signal \&32230\    : AGCBIT;
  signal  \32231\    : AGCBIT; signal  \MON+CH\   : AGCBIT;
  signal  \32232\    : AGCBIT;
  signal  \32233\    : AGCBIT;
  signal  \32234\    : AGCBIT;
  signal \&32235\    : AGCBIT;
  signal  \32236\    : AGCBIT;
  signal  \32237\    : AGCBIT;
  signal  \32238\    : AGCBIT;
  signal \$32238\    : AGCBIT;
  signal  \32239\    : AGCBIT;
  signal \$32239\    : AGCBIT;
  signal \&32240\    : AGCBIT;
  signal  \32241\    : AGCBIT;
  signal  \32242\    : AGCBIT;
  signal  \32243\    : AGCBIT;
  signal  \32244\    : AGCBIT;
  signal \$32244\    : AGCBIT;
  signal  \32245\    : AGCBIT;
  signal \$32245\    : AGCBIT;
  signal  \32246\    : AGCBIT;
  signal  \32247\    : AGCBIT; signal  \INCSET/\  : AGCBIT;
  signal  \32249\    : AGCBIT; signal  \INKL/\    : AGCBIT;
  signal \&32250\    : AGCBIT;
  signal  \32251\    : AGCBIT; signal  \INKL\     : AGCBIT;
  signal \&32253\    : AGCBIT;
  signal  \32254\    : AGCBIT; signal  \RSSB\     : AGCBIT;
  signal  \32255\    : AGCBIT; signal  \BKTF/\    : AGCBIT;
  signal  \32256\    : AGCBIT; signal  \CHINC/\   : AGCBIT;
  signal \&32257\    : AGCBIT;
  signal \&32258\    : AGCBIT;
  signal  \32259\    : AGCBIT;
  signal  \32501\    : AGCBIT;
  signal  \32502\    : AGCBIT;
  signal \$32502\    : AGCBIT;
  signal  \32503\    : AGCBIT;
  signal \$32503\    : AGCBIT;
  signal  \32504\    : AGCBIT;
  signal  \32505\    : AGCBIT;
  signal  \32506\    : AGCBIT;
  signal \$32506\    : AGCBIT;
  signal  \32507\    : AGCBIT;
  signal \$32507\    : AGCBIT;
  signal  \32508\    : AGCBIT; signal  \C42A\     : AGCBIT;
  signal  \32509\    : AGCBIT;
  signal \$32509\    : AGCBIT;
  signal  \32510\    : AGCBIT;
  signal \$32510\    : AGCBIT;
  signal  \32511\    : AGCBIT;
  signal  \32512\    : AGCBIT; signal  \C42R\     : AGCBIT;
  signal  \32513\    : AGCBIT; signal  \C42P\     : AGCBIT;
  signal  \32514\    : AGCBIT; signal  \C42M\     : AGCBIT;
  signal  \32515\    : AGCBIT;
  signal \$32515\    : AGCBIT;
  signal  \32516\    : AGCBIT;
  signal \$32516\    : AGCBIT;
  signal  \32517\    : AGCBIT;
  signal  \32518\    : AGCBIT;
  signal  \32519\    : AGCBIT;
  signal \$32519\    : AGCBIT;
  signal  \32520\    : AGCBIT;
  signal \$32520\    : AGCBIT;
  signal  \32521\    : AGCBIT; signal  \C43A\     : AGCBIT;
  signal  \32522\    : AGCBIT;
  signal  \32523\    : AGCBIT; signal  \CG15\     : AGCBIT;
  signal  \32524\    : AGCBIT;
  signal \$32524\    : AGCBIT;
  signal  \32525\    : AGCBIT;
  signal \$32525\    : AGCBIT;
  signal  \32526\    : AGCBIT; signal  \C43R\     : AGCBIT;
  signal  \32527\    : AGCBIT; signal  \C43P\     : AGCBIT;
  signal  \32528\    : AGCBIT; signal  \C43M\     : AGCBIT;
  signal  \32529\    : AGCBIT;
  signal \$32529\    : AGCBIT;
  signal  \32530\    : AGCBIT;
  signal \$32530\    : AGCBIT;
  signal  \32531\    : AGCBIT;
  signal  \32532\    : AGCBIT;
  signal \$32532\    : AGCBIT;
  signal  \32533\    : AGCBIT;
  signal \$32533\    : AGCBIT;
  signal  \32534\    : AGCBIT; signal  \C56A\     : AGCBIT;
  signal  \32535\    : AGCBIT; signal  \C56R\     : AGCBIT;
  signal  \32536\    : AGCBIT;
  signal \$32536\    : AGCBIT;
  signal  \32537\    : AGCBIT;
  signal \$32537\    : AGCBIT;
  signal  \32538\    : AGCBIT;
  signal  \32539\    : AGCBIT;
  signal \$32539\    : AGCBIT;
  signal  \32540\    : AGCBIT;
  signal \$32540\    : AGCBIT;
  signal  \32541\    : AGCBIT; signal  \C57A\     : AGCBIT;
  signal  \32542\    : AGCBIT; signal  \C57R\     : AGCBIT;
  signal  \32543\    : AGCBIT;
  signal \$32543\    : AGCBIT;
  signal  \32544\    : AGCBIT;
  signal \$32544\    : AGCBIT;
  signal  \32545\    : AGCBIT;
  signal  \32546\    : AGCBIT;
  signal \$32546\    : AGCBIT;
  signal  \32547\    : AGCBIT;
  signal \$32547\    : AGCBIT;
  signal \&32548\    : AGCBIT;
  signal  \32549\    : AGCBIT; signal  \C60A\     : AGCBIT;
  signal  \32550\    : AGCBIT; signal  \CTROR/\   : AGCBIT;
  signal \&32551\    : AGCBIT;
  signal  \32552\    : AGCBIT; signal  \CTROR\    : AGCBIT;
  signal  \32553\    : AGCBIT; signal  \C60R\     : AGCBIT;
  signal  \32554\    : AGCBIT; signal  \CA5/\     : AGCBIT;
  signal  \32556\    : AGCBIT; signal  \CXB5/\    : AGCBIT;
  signal  \32558\    : AGCBIT; signal  \CHINC\    : AGCBIT;
  signal  \32601\    : AGCBIT;
  signal  \32602\    : AGCBIT;
  signal \$32602\    : AGCBIT;
  signal  \32603\    : AGCBIT;
  signal \$32603\    : AGCBIT;
  signal  \32604\    : AGCBIT;
  signal  \32605\    : AGCBIT;
  signal  \32606\    : AGCBIT;
  signal \$32606\    : AGCBIT;
  signal  \32607\    : AGCBIT;
  signal \$32607\    : AGCBIT;
  signal  \32608\    : AGCBIT; signal  \C44A\     : AGCBIT;
  signal  \32609\    : AGCBIT;
  signal \$32609\    : AGCBIT;
  signal  \32610\    : AGCBIT;
  signal \$32610\    : AGCBIT;
  signal  \32611\    : AGCBIT;
  signal  \32612\    : AGCBIT; signal  \C44R\     : AGCBIT;
  signal  \32613\    : AGCBIT; signal  \C44P\     : AGCBIT;
  signal  \32614\    : AGCBIT; signal  \C44M\     : AGCBIT;
  signal  \32615\    : AGCBIT;
  signal \$32615\    : AGCBIT;
  signal  \32616\    : AGCBIT;
  signal \$32616\    : AGCBIT;
  signal  \32617\    : AGCBIT;
  signal  \32618\    : AGCBIT;
  signal  \32619\    : AGCBIT;
  signal \$32619\    : AGCBIT;
  signal  \32620\    : AGCBIT;
  signal \$32620\    : AGCBIT;
  signal  \32621\    : AGCBIT; signal  \C45A\     : AGCBIT;
  signal  \32622\    : AGCBIT;
  signal  \32623\    : AGCBIT; signal  \CG16\     : AGCBIT;
  signal  \32624\    : AGCBIT;
  signal \$32624\    : AGCBIT;
  signal  \32625\    : AGCBIT;
  signal \$32625\    : AGCBIT;
  signal  \32626\    : AGCBIT; signal  \C45R\     : AGCBIT;
  signal  \32627\    : AGCBIT; signal  \C45P\     : AGCBIT;
  signal  \32628\    : AGCBIT; signal  \C45M\     : AGCBIT;
  signal  \32629\    : AGCBIT;
  signal \$32629\    : AGCBIT;
  signal  \32630\    : AGCBIT;
  signal \$32630\    : AGCBIT;
  signal  \32631\    : AGCBIT;
  signal  \32632\    : AGCBIT;
  signal \$32632\    : AGCBIT;
  signal  \32633\    : AGCBIT;
  signal \$32633\    : AGCBIT;
  signal  \32634\    : AGCBIT; signal  \C46A\     : AGCBIT;
  signal  \32635\    : AGCBIT; signal  \C46R\     : AGCBIT;
  signal  \32636\    : AGCBIT;
  signal \$32636\    : AGCBIT;
  signal  \32637\    : AGCBIT;
  signal \$32637\    : AGCBIT;
  signal  \32638\    : AGCBIT;
  signal  \32639\    : AGCBIT; signal  \C46P\     : AGCBIT;
  signal  \32640\    : AGCBIT; signal  \C46M\     : AGCBIT;
  signal  \32643\    : AGCBIT;
  signal \$32643\    : AGCBIT;
  signal  \32644\    : AGCBIT;
  signal \$32644\    : AGCBIT;
  signal  \32645\    : AGCBIT;
  signal  \32646\    : AGCBIT;
  signal \$32646\    : AGCBIT;
  signal  \32647\    : AGCBIT;
  signal \$32647\    : AGCBIT;
  signal  \32649\    : AGCBIT; signal  \C47A\     : AGCBIT;
  signal  \32650\    : AGCBIT;
  signal  \32652\    : AGCBIT; signal  \CG26\     : AGCBIT;
  signal  \32653\    : AGCBIT; signal  \C47R\     : AGCBIT;
  signal  \32654\    : AGCBIT; signal  \CXB0/\    : AGCBIT;
  signal  \32656\    : AGCBIT; signal  \CXB6/\    : AGCBIT;
  signal  \32658\    : AGCBIT; signal  \RQ/\      : AGCBIT;
  signal  \47101\    : AGCBIT;
  signal  \47102\    : AGCBIT; signal  \DLKCLR\   : AGCBIT;
  signal  \47104\    : AGCBIT;
  signal \$47104\    : AGCBIT;
  signal  \47105\    : AGCBIT; signal  \RDOUT/\   : AGCBIT;
  signal \$47105\    : AGCBIT;
  signal  \47106\    : AGCBIT; signal  \ADVCTR\   : AGCBIT;
  signal  \47107\    : AGCBIT;
  signal  \47108\    : AGCBIT;
  signal  \47109\    : AGCBIT; signal  \1CNT\     : AGCBIT;
  signal \$47109\    : AGCBIT;
  signal  \47110\    : AGCBIT;
  signal \$47110\    : AGCBIT;
  signal  \47111\    : AGCBIT;
  signal \$47111\    : AGCBIT;
  signal  \47112\    : AGCBIT;
  signal \$47112\    : AGCBIT;
  signal  \47113\    : AGCBIT;
  signal \$47113\    : AGCBIT;
  signal  \47114\    : AGCBIT;
  signal \$47114\    : AGCBIT;
  signal  \47115\    : AGCBIT; signal  \DKCTR1/\  : AGCBIT;
  signal  \47116\    : AGCBIT; signal  \DKCTR1\   : AGCBIT;
  signal  \47117\    : AGCBIT;
  signal \$47117\    : AGCBIT;
  signal  \47118\    : AGCBIT;
  signal \$47118\    : AGCBIT;
  signal  \47119\    : AGCBIT;
  signal \$47119\    : AGCBIT;
  signal  \47120\    : AGCBIT;
  signal \$47120\    : AGCBIT;
  signal  \47121\    : AGCBIT;
  signal \$47121\    : AGCBIT;
  signal  \47122\    : AGCBIT;
  signal \$47122\    : AGCBIT;
  signal  \47123\    : AGCBIT; signal  \DKCTR2/\  : AGCBIT;
  signal  \47124\    : AGCBIT; signal  \DKCTR2\   : AGCBIT;
  signal  \47125\    : AGCBIT;
  signal \$47125\    : AGCBIT;
  signal  \47126\    : AGCBIT;
  signal \$47126\    : AGCBIT;
  signal  \47127\    : AGCBIT;
  signal \$47127\    : AGCBIT;
  signal  \47128\    : AGCBIT;
  signal \$47128\    : AGCBIT;
  signal  \47129\    : AGCBIT;
  signal \$47129\    : AGCBIT;
  signal  \47130\    : AGCBIT;
  signal \$47130\    : AGCBIT;
  signal  \47131\    : AGCBIT; signal  \DKCTR3/\  : AGCBIT;
  signal  \47132\    : AGCBIT; signal  \DKCTR3\   : AGCBIT;
  signal  \47133\    : AGCBIT;
  signal \$47133\    : AGCBIT;
  signal  \47134\    : AGCBIT;
  signal \$47134\    : AGCBIT;
  signal  \47135\    : AGCBIT;
  signal \$47135\    : AGCBIT;
  signal  \47136\    : AGCBIT;
  signal \$47136\    : AGCBIT;
  signal  \47137\    : AGCBIT; signal  \DKCTR4\   : AGCBIT;
  signal \$47137\    : AGCBIT;
  signal  \47138\    : AGCBIT; signal  \DKCTR4/\  : AGCBIT;
  signal \$47138\    : AGCBIT;
  signal  \47139\    : AGCBIT; signal  \16CNT\    : AGCBIT;
  signal \$47139\    : AGCBIT;
  signal  \47140\    : AGCBIT;
  signal \$47140\    : AGCBIT;
  signal  \47141\    : AGCBIT;
  signal \$47141\    : AGCBIT;
  signal  \47142\    : AGCBIT; signal  \32CNT\    : AGCBIT;
  signal \$47142\    : AGCBIT;
  signal  \47143\    : AGCBIT; signal  \DKCTR5\   : AGCBIT;
  signal \$47143\    : AGCBIT;
  signal  \47144\    : AGCBIT; signal  \DKCTR5/\  : AGCBIT;
  signal \$47144\    : AGCBIT;
  signal  \47145\    : AGCBIT;
  signal  \47147\    : AGCBIT;
  signal \$47147\    : AGCBIT;
  signal  \47148\    : AGCBIT;
  signal \$47148\    : AGCBIT;
  signal  \47149\    : AGCBIT;
  signal \$47149\    : AGCBIT;
  signal  \47150\    : AGCBIT;
  signal \$47150\    : AGCBIT;
  signal  \47151\    : AGCBIT;
  signal \$47151\    : AGCBIT;
  signal  \47153\    : AGCBIT;
  signal \$47153\    : AGCBIT;
  signal  \47154\    : AGCBIT; signal  \WDORDR\   : AGCBIT;
  signal \$47154\    : AGCBIT;
  signal  \47155\    : AGCBIT;
  signal  \47156\    : AGCBIT;
  signal \$47156\    : AGCBIT;
  signal  \47157\    : AGCBIT;
  signal \$47157\    : AGCBIT;
  signal  \47158\    : AGCBIT; signal  \CH1307\   : AGCBIT;
  signal  \47159\    : AGCBIT; signal  \ORDRBT\   : AGCBIT;
  signal  \47161\    : AGCBIT; signal  \F12B/\    : AGCBIT;
  signal  \47162\    : AGCBIT; signal  \F14H\     : AGCBIT;
  signal  \47201\    : AGCBIT;
  signal  \47202\    : AGCBIT; signal  \WCH13/\   : AGCBIT;
  signal  \47205\    : AGCBIT;
  signal  \47206\    : AGCBIT;
  signal  \47207\    : AGCBIT; signal  \CCH13\    : AGCBIT;
  signal  \47210\    : AGCBIT;
  signal  \47211\    : AGCBIT; signal  \RCH13/\   : AGCBIT;
  signal  \47214\    : AGCBIT;
  signal  \47215\    : AGCBIT; signal  \WCH14/\   : AGCBIT;
  signal  \47218\    : AGCBIT;
  signal  \47219\    : AGCBIT;
  signal  \47220\    : AGCBIT; signal  \CCH14\    : AGCBIT;
  signal  \47223\    : AGCBIT;
  signal  \47224\    : AGCBIT; signal  \RCH14/\   : AGCBIT;
  signal  \47227\    : AGCBIT; signal  \BSYNC/\   : AGCBIT;
  signal  \47228\    : AGCBIT;
  signal  \47229\    : AGCBIT; signal  \LOW0/\    : AGCBIT;
  signal  \47230\    : AGCBIT;
  signal  \47231\    : AGCBIT; signal  \LOW1/\    : AGCBIT;
  signal  \47232\    : AGCBIT;
  signal  \47233\    : AGCBIT; signal  \LOW2/\    : AGCBIT;
  signal  \47234\    : AGCBIT;
  signal  \47235\    : AGCBIT; signal  \LOW3/\    : AGCBIT;
  signal  \47236\    : AGCBIT;
  signal  \47237\    : AGCBIT; signal  \LOW4/\    : AGCBIT;
  signal  \47238\    : AGCBIT;
  signal  \47239\    : AGCBIT; signal  \LOW5/\    : AGCBIT;
  signal  \47240\    : AGCBIT;
  signal  \47241\    : AGCBIT; signal  \LOW6/\    : AGCBIT;
  signal  \47242\    : AGCBIT;
  signal  \47243\    : AGCBIT; signal  \LOW7/\    : AGCBIT;
  signal  \47244\    : AGCBIT;
  signal  \47245\    : AGCBIT;
  signal  \47246\    : AGCBIT;
  signal \$47246\    : AGCBIT;
  signal  \47247\    : AGCBIT;
  signal \$47247\    : AGCBIT;
  signal  \47248\    : AGCBIT;
  signal \$47248\    : AGCBIT;
  signal  \47249\    : AGCBIT;
  signal \$47249\    : AGCBIT;
  signal  \47250\    : AGCBIT;
  signal  \47251\    : AGCBIT;
  signal \&47252\    : AGCBIT;
  signal  \47253\    : AGCBIT; signal  \DATA/\    : AGCBIT;
  signal  \47254\    : AGCBIT;
  signal  \47255\    : AGCBIT; signal  \DKDAT/\   : AGCBIT;
  signal  \47256\    : AGCBIT; signal  \DKDATA\   : AGCBIT;
  signal  \47261\    : AGCBIT; signal  \DKDATB\   : AGCBIT;
  signal  \47262\    : AGCBIT; signal  \FS13/\    : AGCBIT;
  signal  \47301\    : AGCBIT;
  signal  \47302\    : AGCBIT;
  signal \$47302\    : AGCBIT;
  signal  \47303\    : AGCBIT;
  signal \$47303\    : AGCBIT;
  signal  \47304\    : AGCBIT; signal  \WRD1BP\   : AGCBIT;
  signal  \47305\    : AGCBIT;
  signal  \47306\    : AGCBIT;
  signal \$47306\    : AGCBIT;
  signal  \47307\    : AGCBIT;
  signal \$47307\    : AGCBIT;
  signal  \47308\    : AGCBIT; signal  \WRD1B1\   : AGCBIT;
  signal  \47309\    : AGCBIT;
  signal  \47310\    : AGCBIT;
  signal \$47310\    : AGCBIT;
  signal  \47311\    : AGCBIT;
  signal \$47311\    : AGCBIT;
  signal  \47312\    : AGCBIT;
  signal  \47313\    : AGCBIT;
  signal  \47314\    : AGCBIT;
  signal \$47314\    : AGCBIT;
  signal  \47315\    : AGCBIT;
  signal \$47315\    : AGCBIT;
  signal  \47316\    : AGCBIT;
  signal  \47317\    : AGCBIT;
  signal  \47318\    : AGCBIT;
  signal \$47318\    : AGCBIT;
  signal  \47319\    : AGCBIT;
  signal \$47319\    : AGCBIT;
  signal  \47320\    : AGCBIT;
  signal \&47321\    : AGCBIT;
  signal  \47322\    : AGCBIT;
  signal  \47323\    : AGCBIT;
  signal \$47323\    : AGCBIT;
  signal  \47324\    : AGCBIT;
  signal \$47324\    : AGCBIT;
  signal  \47325\    : AGCBIT;
  signal  \47326\    : AGCBIT;
  signal  \47327\    : AGCBIT;
  signal \$47327\    : AGCBIT;
  signal  \47328\    : AGCBIT;
  signal \$47328\    : AGCBIT;
  signal  \47329\    : AGCBIT;
  signal  \47330\    : AGCBIT;
  signal  \47331\    : AGCBIT;
  signal \$47331\    : AGCBIT;
  signal  \47332\    : AGCBIT;
  signal \$47332\    : AGCBIT;
  signal  \47333\    : AGCBIT;
  signal \&47334\    : AGCBIT;
  signal  \47335\    : AGCBIT;
  signal  \47336\    : AGCBIT;
  signal \$47336\    : AGCBIT;
  signal  \47337\    : AGCBIT;
  signal \$47337\    : AGCBIT;
  signal  \47338\    : AGCBIT;
  signal  \47339\    : AGCBIT;
  signal  \47340\    : AGCBIT;
  signal \$47340\    : AGCBIT;
  signal  \47341\    : AGCBIT;
  signal \$47341\    : AGCBIT;
  signal  \47342\    : AGCBIT;
  signal \&47343\    : AGCBIT;
  signal  \47344\    : AGCBIT;
  signal  \47345\    : AGCBIT;
  signal \$47345\    : AGCBIT;
  signal  \47346\    : AGCBIT;
  signal \$47346\    : AGCBIT;
  signal  \47347\    : AGCBIT;
  signal  \47348\    : AGCBIT;
  signal  \47349\    : AGCBIT;
  signal \$47349\    : AGCBIT;
  signal  \47350\    : AGCBIT;
  signal \$47350\    : AGCBIT;
  signal  \47351\    : AGCBIT;
  signal  \47352\    : AGCBIT;
  signal  \47353\    : AGCBIT;
  signal \$47353\    : AGCBIT;
  signal  \47354\    : AGCBIT;
  signal \$47354\    : AGCBIT;
  signal  \47355\    : AGCBIT;
  signal  \47356\    : AGCBIT;
  signal  \47357\    : AGCBIT;
  signal \$47357\    : AGCBIT;
  signal  \47358\    : AGCBIT;
  signal \$47358\    : AGCBIT;
  signal  \47359\    : AGCBIT;
  signal \&47360\    : AGCBIT;
  signal  \47401\    : AGCBIT;
  signal  \47402\    : AGCBIT;
  signal \$47402\    : AGCBIT;
  signal  \47403\    : AGCBIT;
  signal \$47403\    : AGCBIT;
  signal  \47404\    : AGCBIT; signal  \WRD2B2\   : AGCBIT;
  signal  \47405\    : AGCBIT;
  signal  \47406\    : AGCBIT;
  signal \$47406\    : AGCBIT;
  signal  \47407\    : AGCBIT;
  signal \$47407\    : AGCBIT;
  signal  \47408\    : AGCBIT; signal  \WRD2B3\   : AGCBIT;
  signal  \47409\    : AGCBIT;
  signal  \47410\    : AGCBIT;
  signal \$47410\    : AGCBIT;
  signal  \47411\    : AGCBIT;
  signal \$47411\    : AGCBIT;
  signal  \47412\    : AGCBIT;
  signal  \47413\    : AGCBIT;
  signal  \47414\    : AGCBIT;
  signal \$47414\    : AGCBIT;
  signal  \47415\    : AGCBIT;
  signal \$47415\    : AGCBIT;
  signal  \47416\    : AGCBIT;
  signal  \47417\    : AGCBIT;
  signal  \47418\    : AGCBIT;
  signal \$47418\    : AGCBIT;
  signal  \47419\    : AGCBIT;
  signal \$47419\    : AGCBIT;
  signal  \47420\    : AGCBIT;
  signal \&47421\    : AGCBIT;
  signal  \47422\    : AGCBIT;
  signal  \47423\    : AGCBIT;
  signal \$47423\    : AGCBIT;
  signal  \47424\    : AGCBIT;
  signal \$47424\    : AGCBIT;
  signal  \47425\    : AGCBIT;
  signal  \47426\    : AGCBIT;
  signal  \47427\    : AGCBIT;
  signal \$47427\    : AGCBIT;
  signal  \47428\    : AGCBIT;
  signal \$47428\    : AGCBIT;
  signal  \47429\    : AGCBIT;
  signal  \47430\    : AGCBIT;
  signal  \47431\    : AGCBIT;
  signal \$47431\    : AGCBIT;
  signal  \47432\    : AGCBIT;
  signal \$47432\    : AGCBIT;
  signal  \47433\    : AGCBIT;
  signal \&47434\    : AGCBIT;
  signal  \47435\    : AGCBIT;
  signal  \47436\    : AGCBIT;
  signal \$47436\    : AGCBIT;
  signal  \47437\    : AGCBIT;
  signal \$47437\    : AGCBIT;
  signal  \47438\    : AGCBIT;
  signal  \47439\    : AGCBIT;
  signal  \47440\    : AGCBIT;
  signal \$47440\    : AGCBIT;
  signal  \47441\    : AGCBIT;
  signal \$47441\    : AGCBIT;
  signal  \47442\    : AGCBIT;
  signal  \47443\    : AGCBIT;
  signal  \47444\    : AGCBIT;
  signal \$47444\    : AGCBIT;
  signal  \47445\    : AGCBIT;
  signal \$47445\    : AGCBIT;
  signal  \47446\    : AGCBIT;
  signal \&47447\    : AGCBIT;
  signal  \47448\    : AGCBIT;
  signal  \47449\    : AGCBIT;
  signal \$47449\    : AGCBIT;
  signal  \47450\    : AGCBIT;
  signal \$47450\    : AGCBIT;
  signal  \47451\    : AGCBIT;
  signal  \47452\    : AGCBIT;
  signal  \47453\    : AGCBIT;
  signal \$47453\    : AGCBIT;
  signal  \47454\    : AGCBIT;
  signal \$47454\    : AGCBIT;
  signal  \47455\    : AGCBIT;
  signal  \47456\    : AGCBIT;
  signal  \47457\    : AGCBIT;
  signal \$47457\    : AGCBIT;
  signal  \47458\    : AGCBIT;
  signal \$47458\    : AGCBIT;
  signal  \47459\    : AGCBIT;
  signal \&47460\    : AGCBIT;
  signal \&48101\    : AGCBIT;
  signal  \48102\    : AGCBIT;
  signal  \48103\    : AGCBIT;
  signal  \48104\    : AGCBIT;
  signal  \48105\    : AGCBIT;
  signal \&48106\    : AGCBIT;
  signal  \48107\    : AGCBIT;
  signal \$48107\    : AGCBIT;
  signal  \48108\    : AGCBIT; signal  \PIPAFL\   : AGCBIT;
  signal \$48108\    : AGCBIT;
  signal  \48109\    : AGCBIT;
  signal  \48110\    : AGCBIT;
  signal  \48111\    : AGCBIT;
  signal \$48111\    : AGCBIT;
  signal  \48112\    : AGCBIT;
  signal \$48112\    : AGCBIT;
  signal  \48113\    : AGCBIT;
  signal \$48113\    : AGCBIT;
  signal  \48114\    : AGCBIT;
  signal \$48114\    : AGCBIT;
  signal  \48115\    : AGCBIT;
  signal  \48116\    : AGCBIT;
  signal \&48117\    : AGCBIT;
  signal  \48118\    : AGCBIT;
  signal  \48119\    : AGCBIT;
  signal  \48120\    : AGCBIT; signal  \WCH35/\   : AGCBIT;
  signal  \48123\    : AGCBIT;
  signal  \48124\    : AGCBIT; signal  \CCH35\    : AGCBIT;
  signal  \48127\    : AGCBIT; signal  \BOTHX\    : AGCBIT;
  signal  \48128\    : AGCBIT;
  signal  \48129\    : AGCBIT;
  signal  \48130\    : AGCBIT;
  signal  \48131\    : AGCBIT;
  signal  \48132\    : AGCBIT;
  signal  \48133\    : AGCBIT;
  signal \$48133\    : AGCBIT;
  signal  \48134\    : AGCBIT;
  signal \$48134\    : AGCBIT;
  signal  \48135\    : AGCBIT;
  signal  \48136\    : AGCBIT;
  signal  \48137\    : AGCBIT;
  signal \$48137\    : AGCBIT;
  signal  \48138\    : AGCBIT;
  signal \$48138\    : AGCBIT;
  signal  \48139\    : AGCBIT;
  signal  \48140\    : AGCBIT;
  signal  \48141\    : AGCBIT;
  signal  \48142\    : AGCBIT;
  signal  \48143\    : AGCBIT;
  signal \$48143\    : AGCBIT;
  signal  \48144\    : AGCBIT;
  signal \$48144\    : AGCBIT;
  signal  \48145\    : AGCBIT;
  signal  \48146\    : AGCBIT;
  signal  \48147\    : AGCBIT;
  signal \$48147\    : AGCBIT;
  signal  \48148\    : AGCBIT;
  signal \$48148\    : AGCBIT;
  signal  \48149\    : AGCBIT; signal  \NOXM\     : AGCBIT;
  signal \$48149\    : AGCBIT;
  signal  \48150\    : AGCBIT;
  signal \$48150\    : AGCBIT;
  signal  \48151\    : AGCBIT; signal  \NOXP\     : AGCBIT;
  signal \$48151\    : AGCBIT;
  signal  \48152\    : AGCBIT;
  signal \$48152\    : AGCBIT;
  signal  \48153\    : AGCBIT; signal  \MISSX\    : AGCBIT;
  signal \$48153\    : AGCBIT;
  signal  \48154\    : AGCBIT;
  signal \$48154\    : AGCBIT;
  signal  \48155\    : AGCBIT; signal  \PIPXP\    : AGCBIT;
  signal  \48156\    : AGCBIT; signal  \PIPXM\    : AGCBIT;
  signal  \48157\    : AGCBIT; signal  \F18B/\    : AGCBIT;
  signal \&48201\    : AGCBIT;
  signal  \48202\    : AGCBIT; signal  \CH01\     : AGCBIT;
  signal \&48203\    : AGCBIT;
  signal  \48204\    : AGCBIT; signal  \CH02\     : AGCBIT;
  signal \&48205\    : AGCBIT;
  signal  \48206\    : AGCBIT; signal  \CH03\     : AGCBIT;
  signal \&48207\    : AGCBIT;
  signal  \48208\    : AGCBIT; signal  \CH04\     : AGCBIT;
  signal \&48209\    : AGCBIT;
  signal \&48210\    : AGCBIT;
  signal  \48211\    : AGCBIT; signal  \CH05\     : AGCBIT;
  signal \&48212\    : AGCBIT;
  signal  \48213\    : AGCBIT; signal  \CH06\     : AGCBIT;
  signal \&48214\    : AGCBIT;
  signal  \48215\    : AGCBIT; signal  \CH07\     : AGCBIT;
  signal \&48216\    : AGCBIT;
  signal \&48217\    : AGCBIT;
  signal  \48218\    : AGCBIT; signal  \CH08\     : AGCBIT;
  signal  \48219\    : AGCBIT;
  signal  \48220\    : AGCBIT;
  signal  \48221\    : AGCBIT; signal  \WCH34/\   : AGCBIT;
  signal  \48224\    : AGCBIT;
  signal  \48225\    : AGCBIT; signal  \CCH34\    : AGCBIT;
  signal  \48228\    : AGCBIT; signal  \BOTHY\    : AGCBIT;
  signal  \48229\    : AGCBIT;
  signal  \48230\    : AGCBIT;
  signal  \48231\    : AGCBIT;
  signal  \48232\    : AGCBIT;
  signal  \48233\    : AGCBIT;
  signal  \48234\    : AGCBIT;
  signal \$48234\    : AGCBIT;
  signal  \48235\    : AGCBIT;
  signal \$48235\    : AGCBIT;
  signal  \48236\    : AGCBIT;
  signal  \48237\    : AGCBIT;
  signal  \48238\    : AGCBIT;
  signal \$48238\    : AGCBIT;
  signal  \48239\    : AGCBIT;
  signal \$48239\    : AGCBIT;
  signal  \48240\    : AGCBIT;
  signal  \48241\    : AGCBIT;
  signal  \48242\    : AGCBIT;
  signal  \48243\    : AGCBIT;
  signal  \48244\    : AGCBIT;
  signal \$48244\    : AGCBIT;
  signal  \48245\    : AGCBIT;
  signal \$48245\    : AGCBIT;
  signal  \48246\    : AGCBIT;
  signal  \48247\    : AGCBIT;
  signal  \48248\    : AGCBIT;
  signal \$48248\    : AGCBIT;
  signal  \48249\    : AGCBIT;
  signal \$48249\    : AGCBIT;
  signal  \48250\    : AGCBIT; signal  \PIPYP\    : AGCBIT;
  signal  \48251\    : AGCBIT; signal  \PIPYM\    : AGCBIT;
  signal  \48252\    : AGCBIT; signal  \NOYM\     : AGCBIT;
  signal \$48252\    : AGCBIT;
  signal  \48253\    : AGCBIT;
  signal \$48253\    : AGCBIT;
  signal  \48254\    : AGCBIT; signal  \NOYP\     : AGCBIT;
  signal \$48254\    : AGCBIT;
  signal  \48255\    : AGCBIT;
  signal \$48255\    : AGCBIT;
  signal  \48256\    : AGCBIT; signal  \MISSY\    : AGCBIT;
  signal \$48256\    : AGCBIT;
  signal  \48257\    : AGCBIT;
  signal \$48257\    : AGCBIT;
  signal \&48258\    : AGCBIT;
  signal  \48301\    : AGCBIT;
  signal  \48302\    : AGCBIT;
  signal \$48302\    : AGCBIT;
  signal  \48303\    : AGCBIT;
  signal \$48303\    : AGCBIT;
  signal  \48304\    : AGCBIT; signal  \CH1416\   : AGCBIT;
  signal  \48305\    : AGCBIT; signal  \CDUXD\    : AGCBIT;
  signal  \48306\    : AGCBIT;
  signal  \48307\    : AGCBIT;
  signal  \48308\    : AGCBIT; signal  \CDUXDP\   : AGCBIT;
  signal  \48309\    : AGCBIT; signal  \CDUXDM\   : AGCBIT;
  signal  \48310\    : AGCBIT;
  signal  \48311\    : AGCBIT;
  signal  \48312\    : AGCBIT;
  signal \$48312\    : AGCBIT;
  signal  \48313\    : AGCBIT;
  signal \$48313\    : AGCBIT;
  signal  \48314\    : AGCBIT; signal  \CH1414\   : AGCBIT;
  signal  \48315\    : AGCBIT; signal  \CDUYD\    : AGCBIT;
  signal  \48316\    : AGCBIT;
  signal  \48317\    : AGCBIT;
  signal  \48318\    : AGCBIT; signal  \CDUYDP\   : AGCBIT;
  signal  \48319\    : AGCBIT; signal  \CDUYDM\   : AGCBIT;
  signal  \48320\    : AGCBIT;
  signal  \48321\    : AGCBIT;
  signal  \48322\    : AGCBIT;
  signal \$48322\    : AGCBIT;
  signal  \48323\    : AGCBIT; signal  \CH1413\   : AGCBIT;
  signal  \48324\    : AGCBIT;
  signal \$48324\    : AGCBIT;
  signal  \48325\    : AGCBIT; signal  \CDUZD\    : AGCBIT;
  signal  \48326\    : AGCBIT; signal  \CDUZDP\   : AGCBIT;
  signal  \48327\    : AGCBIT;
  signal  \48328\    : AGCBIT;
  signal  \48329\    : AGCBIT; signal  \CDUZDM\   : AGCBIT;
  signal  \48330\    : AGCBIT;
  signal  \48331\    : AGCBIT;
  signal  \48332\    : AGCBIT;
  signal \$48332\    : AGCBIT;
  signal  \48333\    : AGCBIT;
  signal \$48333\    : AGCBIT;
  signal  \48334\    : AGCBIT; signal  \CH1412\   : AGCBIT;
  signal  \48335\    : AGCBIT; signal  \TRUND\    : AGCBIT;
  signal  \48336\    : AGCBIT; signal  \TRNDP\    : AGCBIT;
  signal  \48337\    : AGCBIT;
  signal  \48338\    : AGCBIT;
  signal  \48339\    : AGCBIT; signal  \TRNDM\    : AGCBIT;
  signal  \48340\    : AGCBIT;
  signal  \48341\    : AGCBIT;
  signal  \48342\    : AGCBIT;
  signal \$48342\    : AGCBIT;
  signal  \48343\    : AGCBIT;
  signal \$48343\    : AGCBIT;
  signal  \48344\    : AGCBIT; signal  \CH1411\   : AGCBIT;
  signal  \48345\    : AGCBIT; signal  \SHAFTD\   : AGCBIT;
  signal  \48346\    : AGCBIT;
  signal  \48347\    : AGCBIT;
  signal  \48348\    : AGCBIT; signal  \SHFTDP\   : AGCBIT;
  signal  \48349\    : AGCBIT; signal  \SHFTDM\   : AGCBIT;
  signal  \48350\    : AGCBIT;
  signal  \48351\    : AGCBIT; signal  \POUT/\    : AGCBIT;
  signal  \48353\    : AGCBIT; signal  \MOUT/\    : AGCBIT;
  signal  \48355\    : AGCBIT; signal  \ZOUT/\    : AGCBIT;
  signal  \48357\    : AGCBIT;
  signal  \48358\    : AGCBIT; signal  \T7PHS4/\  : AGCBIT;
  signal  \48359\    : AGCBIT; signal  \T7PHS4\   : AGCBIT;
  signal  \48401\    : AGCBIT;
  signal  \48402\    : AGCBIT;
  signal \$48402\    : AGCBIT;
  signal  \48403\    : AGCBIT; signal  \E5\       : AGCBIT;
  signal \$48403\    : AGCBIT;
  signal  \48404\    : AGCBIT; signal  \CH0705\   : AGCBIT;
  signal  \48405\    : AGCBIT;
  signal  \48406\    : AGCBIT;
  signal \$48406\    : AGCBIT;
  signal  \48407\    : AGCBIT; signal  \E6\       : AGCBIT;
  signal \$48407\    : AGCBIT;
  signal  \48408\    : AGCBIT; signal  \CH0706\   : AGCBIT;
  signal  \48409\    : AGCBIT;
  signal  \48410\    : AGCBIT; signal  \E7/\      : AGCBIT;
  signal \$48410\    : AGCBIT;
  signal  \48411\    : AGCBIT;
  signal \$48411\    : AGCBIT;
  signal  \48412\    : AGCBIT; signal  \CH0707\   : AGCBIT;
  signal  \48413\    : AGCBIT; signal  \CCH07\    : AGCBIT;
  signal  \48414\    : AGCBIT;
  signal  \48415\    : AGCBIT; signal  \WCH07/\   : AGCBIT;
  signal  \48416\    : AGCBIT;
  signal  \48417\    : AGCBIT; signal  \RCH07/\   : AGCBIT;
  signal  \48418\    : AGCBIT;
  signal  \48419\    : AGCBIT;
  signal \$48419\    : AGCBIT;
  signal  \48420\    : AGCBIT;
  signal \$48420\    : AGCBIT;
  signal  \48421\    : AGCBIT; signal  \CH1108\   : AGCBIT;
  signal  \48422\    : AGCBIT; signal  \OT1108\   : AGCBIT;
  signal  \48423\    : AGCBIT;
  signal  \48424\    : AGCBIT;
  signal \$48424\    : AGCBIT;
  signal  \48425\    : AGCBIT;
  signal \$48425\    : AGCBIT;
  signal  \48426\    : AGCBIT; signal  \CH1113\   : AGCBIT;
  signal  \48427\    : AGCBIT; signal  \OT1113\   : AGCBIT;
  signal  \48428\    : AGCBIT;
  signal  \48429\    : AGCBIT;
  signal \$48429\    : AGCBIT;
  signal  \48430\    : AGCBIT;
  signal \$48430\    : AGCBIT;
  signal  \48431\    : AGCBIT; signal  \CH1114\   : AGCBIT;
  signal  \48432\    : AGCBIT; signal  \OT1114\   : AGCBIT;
  signal  \48433\    : AGCBIT;
  signal  \48434\    : AGCBIT;
  signal \$48434\    : AGCBIT;
  signal  \48435\    : AGCBIT;
  signal \$48435\    : AGCBIT;
  signal  \48436\    : AGCBIT; signal  \CH1116\   : AGCBIT;
  signal  \48437\    : AGCBIT; signal  \OT1116\   : AGCBIT;
  signal \&48438\    : AGCBIT;
  signal \&48439\    : AGCBIT;
  signal  \48440\    : AGCBIT; signal  \CH09\     : AGCBIT;
  signal  \48441\    : AGCBIT;
  signal  \48442\    : AGCBIT;
  signal \$48442\    : AGCBIT;
  signal  \48443\    : AGCBIT;
  signal \$48443\    : AGCBIT;
  signal  \48444\    : AGCBIT; signal  \CH1216\   : AGCBIT;
  signal  \48445\    : AGCBIT; signal  \ISSTDC\   : AGCBIT;
  signal  \48446\    : AGCBIT;
  signal  \48447\    : AGCBIT; signal  \T6ON/\    : AGCBIT;
  signal \$48447\    : AGCBIT;
  signal  \48448\    : AGCBIT;
  signal \$48448\    : AGCBIT;
  signal  \48449\    : AGCBIT; signal  \CH1316\   : AGCBIT;
  signal  \48450\    : AGCBIT;
  signal  \48451\    : AGCBIT;
  signal \$48451\    : AGCBIT;
  signal  \48452\    : AGCBIT;
  signal \$48452\    : AGCBIT;
  signal  \48453\    : AGCBIT; signal  \CH1310\   : AGCBIT;
  signal  \48454\    : AGCBIT; signal  \ALTEST\   : AGCBIT;
  signal \&48456\    : AGCBIT;
  signal \&48457\    : AGCBIT;
  signal  \48458\    : AGCBIT; signal  \CH10\     : AGCBIT;
  signal  \49101\    : AGCBIT;
  signal  \49102\    : AGCBIT;
  signal  \49103\    : AGCBIT;
  signal  \49104\    : AGCBIT;
  signal  \49105\    : AGCBIT;
  signal  \49106\    : AGCBIT;
  signal  \49107\    : AGCBIT;
  signal  \49108\    : AGCBIT;
  signal \$49108\    : AGCBIT;
  signal  \49109\    : AGCBIT; signal  \OVNHRP\   : AGCBIT;
  signal  \49110\    : AGCBIT;
  signal  \49111\    : AGCBIT;
  signal  \49112\    : AGCBIT;
  signal \$49112\    : AGCBIT;
  signal  \49113\    : AGCBIT;
  signal  \49114\    : AGCBIT; signal  \WATCHP\   : AGCBIT;
  signal  \49115\    : AGCBIT;
  signal  \49116\    : AGCBIT; signal  \WATCH/\   : AGCBIT;
  signal \$49116\    : AGCBIT;
  signal  \49117\    : AGCBIT; signal  \WATCH\    : AGCBIT;
  signal \&49118\    : AGCBIT;
  signal  \49120\    : AGCBIT;
  signal  \49121\    : AGCBIT; signal  \HIGH0/\   : AGCBIT;
  signal  \49123\    : AGCBIT;
  signal  \49124\    : AGCBIT; signal  \HIGH1/\   : AGCBIT;
  signal  \49126\    : AGCBIT;
  signal  \49127\    : AGCBIT; signal  \HIGH2/\   : AGCBIT;
  signal  \49129\    : AGCBIT;
  signal  \49130\    : AGCBIT; signal  \HIGH3/\   : AGCBIT;
  signal  \49132\    : AGCBIT;
  signal  \49133\    : AGCBIT; signal  \RCHG/\    : AGCBIT;
  signal  \49136\    : AGCBIT;
  signal  \49137\    : AGCBIT; signal  \WCHG/\    : AGCBIT;
  signal  \49140\    : AGCBIT;
  signal  \49141\    : AGCBIT; signal  \CCHG/\    : AGCBIT;
  signal  \49143\    : AGCBIT; signal  \CHWL01/\  : AGCBIT;
  signal  \49145\    : AGCBIT; signal  \CHWL02/\  : AGCBIT;
  signal  \49147\    : AGCBIT; signal  \CHWL03/\  : AGCBIT;
  signal  \49149\    : AGCBIT; signal  \CHWL04/\  : AGCBIT;
  signal  \49151\    : AGCBIT; signal  \CHWL05/\  : AGCBIT;
  signal  \49153\    : AGCBIT; signal  \CHWL06/\  : AGCBIT;
  signal  \49155\    : AGCBIT; signal  \CHWL07/\  : AGCBIT;
  signal  \49157\    : AGCBIT; signal  \CHWL08/\  : AGCBIT;
  signal  \49159\    : AGCBIT; signal  \CHWL09/\  : AGCBIT;
  signal  \49201\    : AGCBIT;
  signal  \49202\    : AGCBIT;
  signal  \49203\    : AGCBIT; signal  \PIPPLS/\  : AGCBIT;
  signal  \49204\    : AGCBIT; signal  \PIPASW\   : AGCBIT;
  signal  \49205\    : AGCBIT; signal  \FS05/\    : AGCBIT;
  signal  \49206\    : AGCBIT; signal  \PIPDAT\   : AGCBIT;
  signal  \49207\    : AGCBIT;
  signal  \49208\    : AGCBIT; signal  \PIPINT\   : AGCBIT;
  signal  \49209\    : AGCBIT; signal  \800SET\   : AGCBIT;
  signal  \49210\    : AGCBIT; signal  \800RST\   : AGCBIT;
  signal  \49211\    : AGCBIT; signal  \3200A\    : AGCBIT;
  signal  \49212\    : AGCBIT; signal  \3200B\    : AGCBIT;
  signal  \49213\    : AGCBIT; signal  \3200C\    : AGCBIT;
  signal  \49214\    : AGCBIT;
  signal  \49215\    : AGCBIT; signal  \3200D\    : AGCBIT;
  signal  \49216\    : AGCBIT;
  signal  \49217\    : AGCBIT; signal  \12KPPS\   : AGCBIT;
  signal  \49218\    : AGCBIT; signal  \RRRST\    : AGCBIT;
  signal  \49219\    : AGCBIT; signal  \LRRST\    : AGCBIT;
  signal  \49220\    : AGCBIT; signal  \25KPPS\   : AGCBIT;
  signal  \49221\    : AGCBIT;
  signal  \49222\    : AGCBIT;
  signal  \49223\    : AGCBIT; signal  \CDUCLK\   : AGCBIT;
  signal  \49224\    : AGCBIT; signal  \SB0/\     : AGCBIT;
  signal  \49226\    : AGCBIT; signal  \SB1/\     : AGCBIT;
  signal  \49228\    : AGCBIT; signal  \SB2/\     : AGCBIT;
  signal  \49230\    : AGCBIT; signal  \F05A/\    : AGCBIT;
  signal  \49232\    : AGCBIT; signal  \F05B/\    : AGCBIT;
  signal  \49234\    : AGCBIT; signal  \F07B/\    : AGCBIT;
  signal  \49235\    : AGCBIT; signal  \CHWL10/\  : AGCBIT;
  signal  \49237\    : AGCBIT; signal  \NISQ\     : AGCBIT;
  signal \&49238\    : AGCBIT;
  signal \&49239\    : AGCBIT;
  signal  \49240\    : AGCBIT;
  signal  \49241\    : AGCBIT; signal  \RCHAT/\   : AGCBIT;
  signal  \49244\    : AGCBIT;
  signal  \49245\    : AGCBIT; signal  \RCHBT/\   : AGCBIT;
  signal  \49248\    : AGCBIT;
  signal  \49249\    : AGCBIT; signal  \ELSNCN\   : AGCBIT;
  signal  \49250\    : AGCBIT; signal  \ELSNCM\   : AGCBIT;
  signal  \49252\    : AGCBIT; signal  \OT1110\   : AGCBIT;
  signal  \49253\    : AGCBIT; signal  \OT1111\   : AGCBIT;
  signal  \49254\    : AGCBIT; signal  \OT1112\   : AGCBIT;
  signal  \49301\    : AGCBIT;
  signal  \49302\    : AGCBIT;
  signal  \49303\    : AGCBIT; signal  \NOZM\     : AGCBIT;
  signal \$49303\    : AGCBIT;
  signal  \49304\    : AGCBIT;
  signal \$49304\    : AGCBIT;
  signal  \49305\    : AGCBIT; signal  \NOZP\     : AGCBIT;
  signal \$49305\    : AGCBIT;
  signal  \49306\    : AGCBIT;
  signal \$49306\    : AGCBIT;
  signal  \49307\    : AGCBIT; signal  \MISSZ\    : AGCBIT;
  signal \$49307\    : AGCBIT;
  signal  \49308\    : AGCBIT;
  signal \$49308\    : AGCBIT;
  signal  \49309\    : AGCBIT; signal  \BOTHZ\    : AGCBIT;
  signal  \49310\    : AGCBIT;
  signal  \49311\    : AGCBIT;
  signal  \49312\    : AGCBIT;
  signal \$49312\    : AGCBIT;
  signal  \49313\    : AGCBIT;
  signal \$49313\    : AGCBIT;
  signal  \49314\    : AGCBIT;
  signal  \49315\    : AGCBIT;
  signal  \49316\    : AGCBIT;
  signal \$49316\    : AGCBIT;
  signal  \49317\    : AGCBIT;
  signal \$49317\    : AGCBIT;
  signal  \49318\    : AGCBIT;
  signal  \49319\    : AGCBIT;
  signal  \49320\    : AGCBIT;
  signal  \49321\    : AGCBIT;
  signal  \49322\    : AGCBIT;
  signal  \49323\    : AGCBIT;
  signal \$49323\    : AGCBIT;
  signal  \49324\    : AGCBIT;
  signal \$49324\    : AGCBIT;
  signal  \49325\    : AGCBIT;
  signal  \49326\    : AGCBIT;
  signal  \49327\    : AGCBIT;
  signal \$49327\    : AGCBIT;
  signal  \49328\    : AGCBIT;
  signal \$49328\    : AGCBIT;
  signal  \49329\    : AGCBIT; signal  \PIPZP\    : AGCBIT;
  signal  \49330\    : AGCBIT; signal  \PIPZM\    : AGCBIT;
  signal  \49331\    : AGCBIT; signal  \CNTRSB/\  : AGCBIT;
  signal  \49332\    : AGCBIT; signal  \RSCT/\    : AGCBIT;
  signal \&49334\    : AGCBIT;
  signal \&49335\    : AGCBIT;
  signal  \49336\    : AGCBIT; signal  \US2SG\    : AGCBIT;
  signal  \49337\    : AGCBIT; signal  \U2BBKG/\  : AGCBIT;
  signal \&49339\    : AGCBIT;
  signal  \49341\    : AGCBIT;
  signal  \49342\    : AGCBIT;
  signal  \49343\    : AGCBIT; signal  \GTSET\    : AGCBIT;
  signal  \49344\    : AGCBIT; signal  \GTSET/\   : AGCBIT;
  signal  \49345\    : AGCBIT; signal  \GTRST\    : AGCBIT;
  signal  \49346\    : AGCBIT; signal  \GTONE\    : AGCBIT;
  signal \&49347\    : AGCBIT;
  signal  \49348\    : AGCBIT; signal  \FS09/\    : AGCBIT;
  signal  \49351\    : AGCBIT;
  signal  \49352\    : AGCBIT; signal  \F09D\     : AGCBIT;
  signal  \49353\    : AGCBIT; signal  \F09A/\    : AGCBIT;
  signal  \49354\    : AGCBIT; signal  \CI\       : AGCBIT;
  signal  \49355\    : AGCBIT;
  signal  \49356\    : AGCBIT;
  signal  \49357\    : AGCBIT; signal  \F07D/\    : AGCBIT;
  signal  \49358\    : AGCBIT; signal  \F07C/\    : AGCBIT;
  signal  \49359\    : AGCBIT;
  signal  \49360\    : AGCBIT; signal  \F7CSB1/\  : AGCBIT;
  signal  \49409\    : AGCBIT; signal  \FLASH\    : AGCBIT;
  signal  \49410\    : AGCBIT; signal  \FLASH/\   : AGCBIT;
  signal  \49411\    : AGCBIT; signal  \ONE\      : AGCBIT;
  signal  \49412\    : AGCBIT;
  signal \$49412\    : AGCBIT;
  signal  \49413\    : AGCBIT; signal  \CDUSTB/\  : AGCBIT;
  signal \$49413\    : AGCBIT;
  signal  \49414\    : AGCBIT; signal  \PHS3/\    : AGCBIT;
  signal  \49418\    : AGCBIT; signal  \F04B/\    : AGCBIT;
  signal  \49419\    : AGCBIT; signal  \IC11/\    : AGCBIT;
  signal  \49420\    : AGCBIT; signal  \F05D\     : AGCBIT;
  signal  \49425\    : AGCBIT; signal  \CHWL11/\  : AGCBIT;
  signal  \49427\    : AGCBIT; signal  \CHWL12/\  : AGCBIT;
  signal  \49429\    : AGCBIT; signal  \CHWL13/\  : AGCBIT;
  signal  \49431\    : AGCBIT; signal  \CHWL14/\  : AGCBIT;
  signal  \49433\    : AGCBIT; signal  \CHWL16/\  : AGCBIT;
  signal \&49435\    : AGCBIT;
  signal \&49436\    : AGCBIT;
  signal \&49437\    : AGCBIT;
  signal \&49438\    : AGCBIT;
  signal \&49439\    : AGCBIT;
  signal \&49440\    : AGCBIT;
  signal \&49441\    : AGCBIT;
  signal \&49442\    : AGCBIT;
  signal \&49443\    : AGCBIT;
  signal  \1A\       : AGCBIT;
  signal  \2A\       : AGCBIT;
  signal  \2B\       : AGCBIT;
  signal  \3A\       : AGCBIT;
  signal  \3B\       : AGCBIT;
  signal  \4A\       : AGCBIT;
  signal  \4B\       : AGCBIT;
  signal  \5A\       : AGCBIT;
  signal  \6A\       : AGCBIT;
  signal  \6B\       : AGCBIT;
  signal \$6B\       : AGCBIT;
  signal  \7A\       : AGCBIT;
  signal  \8A\       : AGCBIT;
  signal  \1B\       : AGCBIT;
  signal \&10A\      : AGCBIT;
  signal \&10B\      : AGCBIT;
  signal  \5B\       : AGCBIT;
  signal  \8B\       : AGCBIT;
  signal  \9A\       : AGCBIT;
  signal  \12A\      : AGCBIT;
  signal  \11A\      : AGCBIT;
  signal  \13A\      : AGCBIT;
  signal  \14A\      : AGCBIT;
  signal  \15A\      : AGCBIT;
  signal  \16A\      : AGCBIT;
  signal  \17A\      : AGCBIT;
  signal  \18A\      : AGCBIT;
  signal  \19A\      : AGCBIT;
  signal  \20A\      : AGCBIT;
  signal  \11B\      : AGCBIT;
  signal \$11B\      : AGCBIT;
  signal  \21B\      : AGCBIT;
  signal  \13B\      : AGCBIT;
  signal \$13B\      : AGCBIT;
  signal  \22B\      : AGCBIT;
  signal  \14B\      : AGCBIT;
  signal \$14B\      : AGCBIT;
  signal  \23B\      : AGCBIT;
  signal  \15B\      : AGCBIT;
  signal \$15B\      : AGCBIT;
  signal  \24B\      : AGCBIT;
  signal  \16B\      : AGCBIT;
  signal \$16B\      : AGCBIT;
  signal  \25B\      : AGCBIT;
  signal  \17B\      : AGCBIT;
  signal \$17B\      : AGCBIT;
  signal  \26B\      : AGCBIT;
  signal  \18B\      : AGCBIT;
  signal \$18B\      : AGCBIT;
  signal  \27B\      : AGCBIT;
  signal  \19B\      : AGCBIT;
  signal \$19B\      : AGCBIT;
  signal  \28B\      : AGCBIT;
  signal  \20B\      : AGCBIT;
  signal \$20B\      : AGCBIT;
  signal  \29B\      : AGCBIT;
  signal  \21A\      : AGCBIT; signal  \MDT01\    : AGCBIT;
  signal  \22A\      : AGCBIT; signal  \MDT02\    : AGCBIT;
  signal  \23A\      : AGCBIT; signal  \MDT03\    : AGCBIT;
  signal  \24A\      : AGCBIT; signal  \MDT04\    : AGCBIT;
  signal  \25A\      : AGCBIT; signal  \MDT05\    : AGCBIT;
  signal  \26A\      : AGCBIT; signal  \MDT06\    : AGCBIT;
  signal  \27A\      : AGCBIT; signal  \MDT07\    : AGCBIT;
  signal  \28A\      : AGCBIT; signal  \MDT08\    : AGCBIT;
  signal  \29A\      : AGCBIT; signal  \MDT09\    : AGCBIT;
  signal  \PULLD01\  : AGCBIT; signal  \DERHI\    : AGCBIT;
  signal  \PULLD02\  : AGCBIT; signal  \DERLO\    : AGCBIT;
  signal  \PULLD03\  : AGCBIT; signal  \MDT10\    : AGCBIT;
  signal  \PULLD04\  : AGCBIT; signal  \MDT11\    : AGCBIT;
  signal  \PULLD05\  : AGCBIT; signal  \MDT12\    : AGCBIT;
  signal  \PULLD06\  : AGCBIT; signal  \MDT13\    : AGCBIT;
  signal  \PULLD07\  : AGCBIT; signal  \MDT14\    : AGCBIT;
  signal  \PULLD08\  : AGCBIT; signal  \MDT15\    : AGCBIT;
  signal  \PULLD09\  : AGCBIT; signal  \MDT16\    : AGCBIT;
  signal  \PULLD10\  : AGCBIT; signal  \MNHSBF\   : AGCBIT;
  signal  \PULLD11\  : AGCBIT; signal  \MNHNC\    : AGCBIT;
  signal  \PULLD12\  : AGCBIT; signal  \MNHRPT\   : AGCBIT;
  signal  \PULLD13\  : AGCBIT; signal  \MTCSAI\   : AGCBIT;
  signal  \PULLD14\  : AGCBIT; signal  \MSTRT\    : AGCBIT;
  signal  \PULLD15\  : AGCBIT; signal  \MSTP\     : AGCBIT;
  signal  \PULLD16\  : AGCBIT; signal  \MSBSTP\   : AGCBIT;
  signal  \PULLD17\  : AGCBIT; signal  \MRDCH\    : AGCBIT;
  signal  \PULLD18\  : AGCBIT; signal  \MLDCH\    : AGCBIT;
  signal  \PULLD19\  : AGCBIT; signal  \MONPAR\   : AGCBIT;
  signal  \PULLD20\  : AGCBIT; signal  \MONWBK\   : AGCBIT;
  signal  \PULLD21\  : AGCBIT; signal  \MLOAD\    : AGCBIT;
  signal  \PULLD22\  : AGCBIT; signal  \MREAD\    : AGCBIT;
  signal  \PULLD23\  : AGCBIT; signal  \NHALGA\   : AGCBIT;
  signal  \PULLD24\  : AGCBIT; signal  \DOSCAL\   : AGCBIT;
  signal  \PULLD25\  : AGCBIT; signal  \DBLTST\   : AGCBIT;
  signal  \PULLD26\  : AGCBIT; signal  \MAMU\     : AGCBIT;
  signal  \PULLU01\  : AGCBIT; signal  \MWL01\    : AGCBIT;
  signal  \PULLU02\  : AGCBIT; signal  \MWL02\    : AGCBIT;
  signal  \PULLU03\  : AGCBIT; signal  \MWL03\    : AGCBIT;
  signal  \PULLU04\  : AGCBIT; signal  \MWL04\    : AGCBIT;
  signal  \PULLU05\  : AGCBIT; signal  \MWL05\    : AGCBIT;
  signal  \PULLU06\  : AGCBIT; signal  \MWL06\    : AGCBIT;
  signal  \PULLU07\  : AGCBIT; signal  \MT01\     : AGCBIT;
  signal  \PULLU08\  : AGCBIT; signal  \MWSG\     : AGCBIT;
  signal  \PULLU09\  : AGCBIT; signal  \MT12\     : AGCBIT;
  signal  \PULLU10\  : AGCBIT; signal  \MWCH\     : AGCBIT;
  signal  \PULLU11\  : AGCBIT; signal  \MRCH\     : AGCBIT;
  signal  \PULLU12\  : AGCBIT; signal  \MPAL/\    : AGCBIT;
  signal  \PULLU13\  : AGCBIT; signal  \MT05\     : AGCBIT;
  signal  \PULLU14\  : AGCBIT; signal  \MTCAL/\   : AGCBIT;
  signal  \PULLU15\  : AGCBIT; signal  \MRPTAL/\  : AGCBIT;
  signal  \PULLU16\  : AGCBIT; signal  \MWATCH/\  : AGCBIT;
  signal  \PULLU17\  : AGCBIT; signal  \MVFAIL/\  : AGCBIT;
  signal  \PULLU18\  : AGCBIT; signal  \MCTRAL/\  : AGCBIT;
  signal  \PULLU19\  : AGCBIT; signal  \MSCAFL/\  : AGCBIT;
  signal  \PULLU20\  : AGCBIT; signal  \MSCDBL/\  : AGCBIT;
  signal  \PULLU21\  : AGCBIT; signal  \GEM01\    : AGCBIT;
  signal  \PULLU22\  : AGCBIT; signal  \GEM02\    : AGCBIT;
  signal  \PULLU23\  : AGCBIT; signal  \GEM03\    : AGCBIT;
  signal  \PULLU24\  : AGCBIT; signal  \GEM04\    : AGCBIT;
  signal  \PULLU25\  : AGCBIT; signal  \GEM05\    : AGCBIT;
  signal  \PULLU26\  : AGCBIT; signal  \GEM06\    : AGCBIT;
  signal  \PULLU27\  : AGCBIT; signal  \GEM07\    : AGCBIT;
  signal  \PULLU28\  : AGCBIT; signal  \GEM08\    : AGCBIT;
  signal  \PULLU29\  : AGCBIT; signal  \GEM09\    : AGCBIT;
  signal  \PULLU30\  : AGCBIT; signal  \GEM10\    : AGCBIT;
  signal  \PULLU31\  : AGCBIT; signal  \GEM11\    : AGCBIT;
  signal  \PULLU32\  : AGCBIT; signal  \GEM12\    : AGCBIT;
  signal  \PULLU33\  : AGCBIT; signal  \GEM13\    : AGCBIT;
  signal  \PULLU34\  : AGCBIT; signal  \GEM14\    : AGCBIT;
  signal  \PULLU35\  : AGCBIT; signal  \GEM16\    : AGCBIT;
  signal  \PULLU36\  : AGCBIT; signal  \GEMP\     : AGCBIT;
  signal  \PULLU37\  : AGCBIT; signal  \SBE\      : AGCBIT;
  signal  \PULLU38\  : AGCBIT; signal  \SBF\      : AGCBIT;
  signal  \PULLU39\  : AGCBIT; signal  \ZID\      : AGCBIT;
  signal  \PULLU40\  : AGCBIT; signal  \REX\      : AGCBIT;
  signal  \PULLU41\  : AGCBIT; signal  \REY\      : AGCBIT;
  signal  \PULLU42\  : AGCBIT; signal  \WEX\      : AGCBIT;
  signal  \PULLU43\  : AGCBIT; signal  \WEY\      : AGCBIT;
  signal  \PULLU44\  : AGCBIT; signal  \CLROPE\   : AGCBIT;
  signal  \PULLU45\  : AGCBIT; signal  \FILTIN\   : AGCBIT;
  signal  \PULLU46\  : AGCBIT; signal  \HIMOD\    : AGCBIT;
  signal  \PULLU47\  : AGCBIT; signal  \IHENV\    : AGCBIT;
  signal  \PULLU48\  : AGCBIT; signal  \IL01\     : AGCBIT;
  signal  \PULLU49\  : AGCBIT; signal  \IL01/\    : AGCBIT;
  signal  \PULLU50\  : AGCBIT; signal  \IL02\     : AGCBIT;
  signal  \PULLU51\  : AGCBIT; signal  \IL02/\    : AGCBIT;
  signal  \PULLU52\  : AGCBIT; signal  \IL03\     : AGCBIT;
  signal  \PULLU53\  : AGCBIT; signal  \IL03/\    : AGCBIT;
  signal  \PULLU54\  : AGCBIT; signal  \IL04\     : AGCBIT;
  signal  \PULLU55\  : AGCBIT; signal  \IL04/\    : AGCBIT;
  signal  \PULLU56\  : AGCBIT; signal  \IL05\     : AGCBIT;
  signal  \PULLU57\  : AGCBIT; signal  \IL05/\    : AGCBIT;
  signal  \PULLU58\  : AGCBIT; signal  \IL06\     : AGCBIT;
  signal  \PULLU59\  : AGCBIT; signal  \IL06/\    : AGCBIT;
  signal  \PULLU60\  : AGCBIT; signal  \IL07\     : AGCBIT;
  signal  \PULLU61\  : AGCBIT; signal  \IL07/\    : AGCBIT;
  signal  \PULLU62\  : AGCBIT; signal  \ILP\      : AGCBIT;
  signal  \PULLU63\  : AGCBIT; signal  \ILP/\     : AGCBIT;
  signal  \PULLU64\  : AGCBIT; signal  \LOMOD\    : AGCBIT;
  signal  \PULLU65\  : AGCBIT; signal  \MBR1\     : AGCBIT;
  signal  \PULLU66\  : AGCBIT; signal  \MBR2\     : AGCBIT;
  signal  \PULLU67\  : AGCBIT; signal  \MGOJAM\   : AGCBIT;
  signal  \PULLU68\  : AGCBIT; signal  \MGP/\     : AGCBIT;
  signal  \PULLU69\  : AGCBIT; signal  \MIIP\     : AGCBIT;
  signal  \PULLU70\  : AGCBIT; signal  \MINHL\    : AGCBIT;
  signal  \PULLU71\  : AGCBIT; signal  \MINKL\    : AGCBIT;
  signal  \PULLU72\  : AGCBIT; signal  \MNISQ\    : AGCBIT;
  signal  \PULLU73\  : AGCBIT; signal  \MON800\   : AGCBIT;
  signal  \PULLU74\  : AGCBIT; signal  \MONWT\    : AGCBIT;
  signal  \PULLU75\  : AGCBIT; signal  \MOSCAL/\  : AGCBIT;
  signal  \PULLU76\  : AGCBIT; signal  \MPIPAL/\  : AGCBIT;
  signal  \PULLU77\  : AGCBIT; signal  \MRAG\     : AGCBIT;
  signal  \PULLU78\  : AGCBIT; signal  \MREQIN\   : AGCBIT;
  signal  \PULLU79\  : AGCBIT; signal  \MRGG\     : AGCBIT;
  signal  \PULLU80\  : AGCBIT; signal  \MRLG\     : AGCBIT;
  signal  \PULLU81\  : AGCBIT; signal  \MRSC\     : AGCBIT;
  signal  \PULLU82\  : AGCBIT; signal  \MRULOG\   : AGCBIT;
  signal  \PULLU83\  : AGCBIT; signal  \MSP\      : AGCBIT;
  signal  \PULLU84\  : AGCBIT; signal  \MSQ10\    : AGCBIT;
  signal  \PULLU85\  : AGCBIT; signal  \MSQ11\    : AGCBIT;
  signal  \PULLU86\  : AGCBIT; signal  \MSQ12\    : AGCBIT;
  signal  \PULLU87\  : AGCBIT; signal  \MSQ13\    : AGCBIT;
  signal  \PULLU88\  : AGCBIT; signal  \MSQ14\    : AGCBIT;
  signal  \PULLU89\  : AGCBIT; signal  \MSQ16\    : AGCBIT;
  signal  \PULLU90\  : AGCBIT; signal  \MSQEXT\   : AGCBIT;
  signal  \PULLU91\  : AGCBIT; signal  \MST1\     : AGCBIT;
  signal  \PULLU92\  : AGCBIT; signal  \MST2\     : AGCBIT;
  signal  \PULLU93\  : AGCBIT; signal  \MST3\     : AGCBIT;
  signal  \PULLU94\  : AGCBIT; signal  \MSTPIT/\  : AGCBIT;
  signal  \PULLU95\  : AGCBIT; signal  \MT02\     : AGCBIT;
  signal  \PULLU96\  : AGCBIT; signal  \MT03\     : AGCBIT;
  signal  \PULLU97\  : AGCBIT; signal  \MT04\     : AGCBIT;
  signal  \PULLU98\  : AGCBIT; signal  \MT06\     : AGCBIT;
  signal  \PULLU99\  : AGCBIT; signal  \MT07\     : AGCBIT;
  signal  \PULLU100\ : AGCBIT; signal  \MT08\     : AGCBIT;
  signal  \PULLU101\ : AGCBIT; signal  \MT09\     : AGCBIT;
  signal  \PULLU102\ : AGCBIT; signal  \MT10\     : AGCBIT;
  signal  \PULLU103\ : AGCBIT; signal  \MT11\     : AGCBIT;
  signal  \PULLU104\ : AGCBIT; signal  \MTCSA/\   : AGCBIT;
  signal  \PULLU105\ : AGCBIT; signal  \MWAG\     : AGCBIT;
  signal  \PULLU106\ : AGCBIT; signal  \MWARNF/\  : AGCBIT;
  signal  \PULLU107\ : AGCBIT; signal  \MWBBEG\   : AGCBIT;
  signal  \PULLU108\ : AGCBIT; signal  \MWBG\     : AGCBIT;
  signal  \PULLU109\ : AGCBIT; signal  \MWEBG\    : AGCBIT;
  signal  \PULLU110\ : AGCBIT; signal  \MWFBG\    : AGCBIT;
  signal  \PULLU111\ : AGCBIT; signal  \MWG\      : AGCBIT;
  signal  \PULLU112\ : AGCBIT; signal  \MWL07\    : AGCBIT;
  signal  \PULLU113\ : AGCBIT; signal  \MWL08\    : AGCBIT;
  signal  \PULLU114\ : AGCBIT; signal  \MWL09\    : AGCBIT;
  signal  \PULLU115\ : AGCBIT; signal  \MWL10\    : AGCBIT;
  signal  \PULLU116\ : AGCBIT; signal  \MWL11\    : AGCBIT;
  signal  \PULLU117\ : AGCBIT; signal  \MWL12\    : AGCBIT;
  signal  \PULLU118\ : AGCBIT; signal  \MWL13\    : AGCBIT;
  signal  \PULLU119\ : AGCBIT; signal  \MWL14\    : AGCBIT;
  signal  \PULLU120\ : AGCBIT; signal  \MWL15\    : AGCBIT;
  signal  \PULLU121\ : AGCBIT; signal  \MWL16\    : AGCBIT;
  signal  \PULLU122\ : AGCBIT; signal  \MWLG\     : AGCBIT;
  signal  \PULLU123\ : AGCBIT; signal  \MWQG\     : AGCBIT;
  signal  \PULLU124\ : AGCBIT; signal  \MWYG\     : AGCBIT;
  signal  \PULLU125\ : AGCBIT; signal  \MWZG\     : AGCBIT;
  signal  \PULLU126\ : AGCBIT; signal  \OUTCOM\   : AGCBIT;
  signal  \PULLU127\ : AGCBIT; signal  \Q2A\      : AGCBIT;
  signal  \PULLU128\ : AGCBIT; signal  \RESETA\   : AGCBIT;
  signal  \PULLU129\ : AGCBIT; signal  \RESETB\   : AGCBIT;
  signal  \PULLU130\ : AGCBIT; signal  \RESETC\   : AGCBIT;
  signal  \PULLU131\ : AGCBIT; signal  \RESETD\   : AGCBIT;
  signal  \PULLU132\ : AGCBIT; signal  \ROPER\    : AGCBIT;
  signal  \PULLU133\ : AGCBIT; signal  \ROPES\    : AGCBIT;
  signal  \PULLU134\ : AGCBIT; signal  \ROPET\    : AGCBIT;
  signal  \PULLU135\ : AGCBIT; signal  \RSTKX/\   : AGCBIT;
  signal  \PULLU136\ : AGCBIT; signal  \RSTKY/\   : AGCBIT;
  signal  \PULLU137\ : AGCBIT; signal  \SBYREL/\  : AGCBIT;
  signal  \PULLU138\ : AGCBIT; signal  \SCAS10\   : AGCBIT;
  signal  \PULLU139\ : AGCBIT; signal  \SCAS17\   : AGCBIT;
  signal  \PULLU140\ : AGCBIT; signal  \SETAB\    : AGCBIT;
  signal  \PULLU141\ : AGCBIT; signal  \SETCD\    : AGCBIT;
  signal  \PULLU142\ : AGCBIT; signal  \SETEK\    : AGCBIT;
  signal  \PULLU143\ : AGCBIT; signal  \STR14\    : AGCBIT;
  signal  \PULLU144\ : AGCBIT; signal  \STR19\    : AGCBIT;
  signal  \PULLU145\ : AGCBIT; signal  \STR210\   : AGCBIT;
  signal  \PULLU146\ : AGCBIT; signal  \STR311\   : AGCBIT;
  signal  \PULLU147\ : AGCBIT; signal  \STR412\   : AGCBIT;
  signal  \PULLU148\ : AGCBIT; signal  \STR58\    : AGCBIT;
  signal  \PULLU149\ : AGCBIT; signal  \STR912\   : AGCBIT;
  signal  \PULLU151\ : AGCBIT; signal  \XB0E\     : AGCBIT;
  signal  \PULLU152\ : AGCBIT; signal  \XB1E\     : AGCBIT;
  signal  \PULLU153\ : AGCBIT; signal  \XB2E\     : AGCBIT;
  signal  \PULLU154\ : AGCBIT; signal  \XB3E\     : AGCBIT;
  signal  \PULLU155\ : AGCBIT; signal  \XB4E\     : AGCBIT;
  signal  \PULLU156\ : AGCBIT; signal  \XB5E\     : AGCBIT;
  signal  \PULLU157\ : AGCBIT; signal  \XB6E\     : AGCBIT;
  signal  \PULLU158\ : AGCBIT; signal  \XB7E\     : AGCBIT;
  signal  \PULLU159\ : AGCBIT; signal  \XT0E\     : AGCBIT;
  signal  \PULLU160\ : AGCBIT; signal  \XT1E\     : AGCBIT;
  signal  \PULLU161\ : AGCBIT; signal  \XT2E\     : AGCBIT;
  signal  \PULLU162\ : AGCBIT; signal  \XT3E\     : AGCBIT;
  signal  \PULLU163\ : AGCBIT; signal  \XT4E\     : AGCBIT;
  signal  \PULLU164\ : AGCBIT; signal  \XT5E\     : AGCBIT;
  signal  \PULLU165\ : AGCBIT; signal  \XT6E\     : AGCBIT;
  signal  \PULLU166\ : AGCBIT; signal  \XT7E\     : AGCBIT;
  signal  \PULLU167\ : AGCBIT; signal  \YB0E\     : AGCBIT;
  signal  \PULLU168\ : AGCBIT; signal  \YB1E\     : AGCBIT;
  signal  \PULLU169\ : AGCBIT; signal  \YB2E\     : AGCBIT;
  signal  \PULLU170\ : AGCBIT; signal  \YB3E\     : AGCBIT;
  signal  \PULLU171\ : AGCBIT; signal  \YT0E\     : AGCBIT;
  signal  \PULLU172\ : AGCBIT; signal  \YT1E\     : AGCBIT;
  signal  \PULLU173\ : AGCBIT; signal  \YT2E\     : AGCBIT;
  signal  \PULLU174\ : AGCBIT; signal  \YT3E\     : AGCBIT;
  signal  \PULLU175\ : AGCBIT; signal  \YT4E\     : AGCBIT;
  signal  \PULLU176\ : AGCBIT; signal  \YT5E\     : AGCBIT;
  signal  \PULLU177\ : AGCBIT; signal  \YT6E\     : AGCBIT;
  signal  \PULLU178\ : AGCBIT; signal  \YT7E\     : AGCBIT;

begin

  -- ***************************
  -- ***                     ***
  -- ***  INPUT assignment.  ***
  -- ***                     ***
  -- ***************************

  \SAP\      <= SAXX( 0); -- Parity from Erasable or Fixed memory to G register.
  \SA01\     <= SAXX( 1); -- LSB of data from Erasable or Fixed memory to G register.
  \SA02\     <= SAXX( 2);
  \SA03\     <= SAXX( 3);
  \SA04\     <= SAXX( 4);
  \SA05\     <= SAXX( 5);
  \SA06\     <= SAXX( 6);
  \SA07\     <= SAXX( 7);
  \SA08\     <= SAXX( 8);
  \SA09\     <= SAXX( 9);
  \SA10\     <= SAXX(10);
  \SA11\     <= SAXX(11);
  \SA12\     <= SAXX(12);
  \SA13\     <= SAXX(13);
  \SA14\     <= SAXX(14);
  \SA16\     <= SAXX(15); -- MSB of data from Erasable or Fixed memory to G register.

  \NHVFAL\    <= INPUTS.\NHVFAL\;
  \MAINRS\    <= INPUTS.\MAINRS\;
  \SBYBUT\    <= INPUTS.\SBYBUT\;
  \IN3212\    <= INPUTS.\IN3212\;
  \CAURST\    <= INPUTS.\CAURST\;
  \IN3213\    <= INPUTS.\IN3213\;
  \NKEY1\     <= INPUTS.\NKEY1\;
  \IN3214\    <= INPUTS.\IN3214\;
  \NKEY2\     <= INPUTS.\NKEY2\;
  \MKEY1\     <= INPUTS.\MKEY1\;
  \NKEY3\     <= INPUTS.\NKEY3\;
  \MKEY2\     <= INPUTS.\MKEY2\;
  \NKEY4\     <= INPUTS.\NKEY4\;
  \MKEY3\     <= INPUTS.\MKEY3\;
  \NKEY5\     <= INPUTS.\NKEY5\;
  \MKEY4\     <= INPUTS.\MKEY4\;
  \NAVRST\    <= INPUTS.\NAVRST\;
  \MKEY5\     <= INPUTS.\MKEY5\;
  \IN3216\    <= INPUTS.\IN3216\;
  \GATEX/\    <= INPUTS.\GATEX/\;
  \GATEY/\    <= INPUTS.\GATEY/\;
  \GATEZ/\    <= INPUTS.\GATEZ/\;
  \SIGNX\     <= INPUTS.\SIGNX\;
  \SIGNY\     <= INPUTS.\SIGNY\;
  \SIGNZ\     <= INPUTS.\SIGNZ\;
  \BMGXP\     <= INPUTS.\BMGXP\;
  \CDUXM\     <= INPUTS.\CDUXM\;
  \DKSTRT\    <= INPUTS.\DKSTRT\;
  \BMGXM\     <= INPUTS.\BMGXM\;
  \CDUYP\     <= INPUTS.\CDUYP\;
  \DKEND\     <= INPUTS.\DKEND\;
  \BMGYP\     <= INPUTS.\BMGYP\;
  \CDUYM\     <= INPUTS.\CDUYM\;
  \DKBSNC\    <= INPUTS.\DKBSNC\;
  \BMGYM\     <= INPUTS.\BMGYM\;
  \CDUZP\     <= INPUTS.\CDUZP\;
  \UPL0\      <= INPUTS.\UPL0\;
  \BMGZP\     <= INPUTS.\BMGZP\;
  \CDUZM\     <= INPUTS.\CDUZM\;
  \UPL1\      <= INPUTS.\UPL1\;
  \BMGZM\     <= INPUTS.\BMGZM\;
  \PIPAX+\    <= INPUTS.\PIPAX+\;
  \RRIN0\     <= INPUTS.\RRIN0\;
  \SHAFTP\    <= INPUTS.\SHAFTP\;
  \PIPAX-\    <= INPUTS.\PIPAX-\;
  \RRIN1\     <= INPUTS.\RRIN1\;
  \SHAFTM\    <= INPUTS.\SHAFTM\;
  \PIPAY+\    <= INPUTS.\PIPAY+\;
  \LRIN0\     <= INPUTS.\LRIN0\;
  \TRNP\      <= INPUTS.\TRNP\;
  \PIPAY-\    <= INPUTS.\PIPAY-\;
  \LRIN1\     <= INPUTS.\LRIN1\;
  \TRNM\      <= INPUTS.\TRNM\;
  \PIPAZ+\    <= INPUTS.\PIPAZ+\;
  \XLNK0\     <= INPUTS.\XLNK0\;
  \CDUXP\     <= INPUTS.\CDUXP\;
  \PIPAZ-\    <= INPUTS.\PIPAZ-\;
  \XLNK1\     <= INPUTS.\XLNK1\;
  \ULLTHR\    <= INPUTS.\ULLTHR\;
  \MNIM+Y\    <= INPUTS.\MNIM+Y\;
  \RRPONA\    <= INPUTS.\RRPONA\;
  \LFTOFF\    <= INPUTS.\LFTOFF\;
  \MNIM-Y\    <= INPUTS.\MNIM-Y\;
  \RRRLSC\    <= INPUTS.\RRRLSC\;
  \GUIREL\    <= INPUTS.\GUIREL\;
  \MNIM+R\    <= INPUTS.\MNIM+R\;
  \MANR+P\    <= INPUTS.\MANR+P\;
  \TRAN+X\    <= INPUTS.\TRAN+X\;
  \MNIM-R\    <= INPUTS.\MNIM-R\;
  \MANR-P\    <= INPUTS.\MANR-P\;
  \TRAN-X\    <= INPUTS.\TRAN-X\;
  \TRST9\     <= INPUTS.\TRST9\;
  \MANR+Y\    <= INPUTS.\MANR+Y\;
  \TRAN+Y\    <= INPUTS.\TRAN+Y\;
  \TRST10\    <= INPUTS.\TRST10\;
  \MANR-Y\    <= INPUTS.\MANR-Y\;
  \TRAN-Y\    <= INPUTS.\TRAN-Y\;
  \HOLFUN\    <= INPUTS.\HOLFUN\;
  \MANR+R\    <= INPUTS.\MANR+R\;
  \TRAN+Z\    <= INPUTS.\TRAN+Z\;
  \FREFUN\    <= INPUTS.\FREFUN\;
  \MANR-R\    <= INPUTS.\MANR-R\;
  \TRAN-Z\    <= INPUTS.\TRAN-Z\;
  \S4BSAB\    <= INPUTS.\S4BSAB\;
  \ISSTOR\    <= INPUTS.\ISSTOR\;
  \OPCDFL\    <= INPUTS.\OPCDFL\;
  \SMSEPR\    <= INPUTS.\SMSEPR\;
  \OPCDEL\    <= INPUTS.\OPCDEL\;
  \MRKRST\    <= INPUTS.\MRKRST\;
  \IN3008\    <= INPUTS.\IN3008\;
  \CDUFAL\    <= INPUTS.\CDUFAL\;
  \ZEROP\     <= INPUTS.\ZEROP\;
  \BLKUPL/\   <= INPUTS.\BLKUPL/\;
  \TEMPIN\    <= INPUTS.\TEMPIN\;
  \MARK\      <= INPUTS.\MARK\;
  \SPSRDY\    <= INPUTS.\SPSRDY\;
  \IMUFAL\    <= INPUTS.\IMUFAL\;
  \OPMSW3\    <= INPUTS.\OPMSW3\;
  \GCAPCL\    <= INPUTS.\GCAPCL\;
  \LEMATT\    <= INPUTS.\LEMATT\;
  \MRKREJ\    <= INPUTS.\MRKREJ\;
  \ROLGOF\    <= INPUTS.\ROLGOF\;
  \IMUOPR\    <= INPUTS.\IMUOPR\;
  \STRPRS\    <= INPUTS.\STRPRS\;
  \PCHGOF\    <= INPUTS.\PCHGOF\;
  \IMUCAG\    <= INPUTS.\IMUCAG\;
  \MNIM+P\    <= INPUTS.\MNIM+P\;
  \LVDAGD\    <= INPUTS.\LVDAGD\;
  \IN3301\    <= INPUTS.\IN3301\;
  \MNIM-P\    <= INPUTS.\MNIM-P\;
  \LRRLSC\    <= INPUTS.\LRRLSC\;
  \CTLSAT\    <= INPUTS.\CTLSAT\;
  \2FSFAL\    <= INPUTS.\2FSFAL\;
  \FLTOUT\    <= INPUTS.\FLTOUT\;
  \OPMSW2\    <= INPUTS.\OPMSW2\;
  \SCAFAL\    <= INPUTS.\SCAFAL\;
  \STRT2\     <= INPUTS.\STRT2\;
  \VFAIL\     <= INPUTS.\VFAIL\;

  -- *****************************
  -- ***                       ***
  -- ***  AGC logic for real!  ***
  -- ***                       ***
  -- *****************************

  -- *************************
  -- ***                   ***
  -- ***  A1 /1 - SCALER.  ***
  -- ***                   ***
  -- *************************

  -- Alias \CHAT05\   
  \=38101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38101\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F10A\     
  \=38102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38102\,
                  I0 =>  \38104\,
                  I1 =>  \38103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38103\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38103\,
                   R => SYSRESET,
                   S => '0' );

  \=38103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38103\,
                  I0 =>  \38102\,
                  I1 =>  \F09A\,
                  I2 =>  \38105\,
                  I3 =>  '0' );

  \:38104\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38104\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38104\,
                   R => SYSRESET,
                   S => '0' );

  \=38104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38104\,
                  I0 =>  \38103\,
                  I1 =>  \38106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38105\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38105\,
                   R => SYSRESET,
                   S => '0' );

  \=38105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38105\,
                  I0 =>  \38103\,
                  I1 =>  \F09A\,
                  I2 =>  \38107\,
                  I3 =>  '0' );

  -- Alias \FS10\     
  \=38106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38106\,
                  I0 =>  \38104\,
                  I1 =>  \38105\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F10B\     
  \=38107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38107\,
                  I0 =>  \38105\,
                  I1 =>  \38106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT06\   
  \=38111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38111\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F11A\     
  \=38112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38112\,
                  I0 =>  \38114\,
                  I1 =>  \38113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38113\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38113\,
                   R => SYSRESET,
                   S => '0' );

  \=38113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38113\,
                  I0 =>  \38112\,
                  I1 =>  \F10A\,
                  I2 =>  \38115\,
                  I3 =>  '0' );

  \:38114\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38114\,
                   R => SYSRESET,
                   S => '0' );

  \=38114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38114\,
                  I0 =>  \38113\,
                  I1 =>  \38116\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38115\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38115\,
                   R => SYSRESET,
                   S => '0' );

  \=38115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38115\,
                  I0 =>  \38113\,
                  I1 =>  \F10A\,
                  I2 =>  \38117\,
                  I3 =>  '0' );

  -- Alias \FS11\     
  \=38116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38116\,
                  I0 =>  \38114\,
                  I1 =>  \38115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F11B\     
  \=38117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38117\,
                  I0 =>  \38115\,
                  I1 =>  \38116\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT07\   
  \=38121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38121\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F12A\     
  \=38122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38122\,
                  I0 =>  \38124\,
                  I1 =>  \38123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38123\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38123\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38123\,
                   R => SYSRESET,
                   S => '0' );

  \=38123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38123\,
                  I0 =>  \38122\,
                  I1 =>  \F11A\,
                  I2 =>  \38125\,
                  I3 =>  '0' );

  \:38124\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38124\,
                   R => SYSRESET,
                   S => '0' );

  \=38124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38124\,
                  I0 =>  \38123\,
                  I1 =>  \38126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38125\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38125\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38125\,
                   R => SYSRESET,
                   S => '0' );

  \=38125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38125\,
                  I0 =>  \38123\,
                  I1 =>  \F11A\,
                  I2 =>  \38127\,
                  I3 =>  '0' );

  -- Alias \FS12\     
  \=38126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38126\,
                  I0 =>  \38124\,
                  I1 =>  \38125\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F12B\     
  \=38127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38127\,
                  I0 =>  \38125\,
                  I1 =>  \38126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT08\   
  \=38131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38131\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F13A\     
  \=38132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38132\,
                  I0 =>  \38134\,
                  I1 =>  \38133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38133\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38133\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38133\,
                   R => SYSRESET,
                   S => '0' );

  \=38133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38133\,
                  I0 =>  \38132\,
                  I1 =>  \F12A\,
                  I2 =>  \38135\,
                  I3 =>  '0' );

  \:38134\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38134\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38134\,
                   R => SYSRESET,
                   S => '0' );

  \=38134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38134\,
                  I0 =>  \38133\,
                  I1 =>  \38136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38135\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38135\,
                   R => SYSRESET,
                   S => '0' );

  \=38135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38135\,
                  I0 =>  \38133\,
                  I1 =>  \F12A\,
                  I2 =>  \38137\,
                  I3 =>  '0' );

  -- Alias \FS13\     
  \=38136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38136\,
                  I0 =>  \38134\,
                  I1 =>  \38135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F13B\     
  \=38137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38137\,
                  I0 =>  \38135\,
                  I1 =>  \38136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT09\   
  \=38141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38141\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F14A\     
  \=38142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38142\,
                  I0 =>  \38144\,
                  I1 =>  \38143\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38143\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38143\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38143\,
                   R => SYSRESET,
                   S => '0' );

  \=38143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38143\,
                  I0 =>  \38142\,
                  I1 =>  \F13A\,
                  I2 =>  \38145\,
                  I3 =>  '0' );

  \:38144\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38144\,
                   R => SYSRESET,
                   S => '0' );

  \=38144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38144\,
                  I0 =>  \38143\,
                  I1 =>  \38146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38145\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38145\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38145\,
                   R => SYSRESET,
                   S => '0' );

  \=38145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38145\,
                  I0 =>  \38143\,
                  I1 =>  \F13A\,
                  I2 =>  \38147\,
                  I3 =>  '0' );

  -- Alias \FS14\     
  \=38146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38146\,
                  I0 =>  \38144\,
                  I1 =>  \38145\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F14B\     
  \=38147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38147\,
                  I0 =>  \38145\,
                  I1 =>  \38146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT10\   
  \=38151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38151\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F15A\     
  \=38152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38152\,
                  I0 =>  \38154\,
                  I1 =>  \38153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38153\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38153\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38153\,
                   R => SYSRESET,
                   S => '0' );

  \=38153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38153\,
                  I0 =>  \38152\,
                  I1 =>  \F14A\,
                  I2 =>  \38155\,
                  I3 =>  '0' );

  \:38154\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38154\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38154\,
                   R => SYSRESET,
                   S => '0' );

  \=38154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38154\,
                  I0 =>  \38153\,
                  I1 =>  \38156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38155\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38155\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38155\,
                   R => SYSRESET,
                   S => '0' );

  \=38155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38155\,
                  I0 =>  \38153\,
                  I1 =>  \F14A\,
                  I2 =>  \38157\,
                  I3 =>  '0' );

  -- Alias \FS15\     
  \=38156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38156\,
                  I0 =>  \38154\,
                  I1 =>  \38155\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F15B\     
  \=38157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38157\,
                  I0 =>  \38155\,
                  I1 =>  \38156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT11\   
  \=38161\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38161\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38164\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F16A\     
  \=38162\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38162\,
                  I0 =>  \38164\,
                  I1 =>  \38163\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38163\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38163\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38163\,
                   R => SYSRESET,
                   S => '0' );

  \=38163\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38163\,
                  I0 =>  \38162\,
                  I1 =>  \F15A\,
                  I2 =>  \38165\,
                  I3 =>  '0' );

  \:38164\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38164\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38164\,
                   R => SYSRESET,
                   S => '0' );

  \=38164\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38164\,
                  I0 =>  \38163\,
                  I1 =>  \38166\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38165\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38165\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38165\,
                   R => SYSRESET,
                   S => '0' );

  \=38165\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38165\,
                  I0 =>  \38163\,
                  I1 =>  \F15A\,
                  I2 =>  \38167\,
                  I3 =>  '0' );

  -- Alias \FS16\     
  \=38166\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38166\,
                  I0 =>  \38164\,
                  I1 =>  \38165\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F16B\     
  \=38167\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38167\,
                  I0 =>  \38165\,
                  I1 =>  \38166\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT12\   
  \=38171\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38171\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38174\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F17A\     
  \=38172\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38172\,
                  I0 =>  \38174\,
                  I1 =>  \38173\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38173\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38173\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38173\,
                   R => SYSRESET,
                   S => '0' );

  \=38173\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38173\,
                  I0 =>  \38172\,
                  I1 =>  \F16A\,
                  I2 =>  \38175\,
                  I3 =>  '0' );

  \:38174\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38174\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38174\,
                   R => SYSRESET,
                   S => '0' );

  \=38174\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38174\,
                  I0 =>  \38173\,
                  I1 =>  \38176\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38175\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38175\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38175\,
                   R => SYSRESET,
                   S => '0' );

  \=38175\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38175\,
                  I0 =>  \38173\,
                  I1 =>  \F16A\,
                  I2 =>  \38177\,
                  I3 =>  '0' );

  -- Alias \FS17\     
  \=38176\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38176\,
                  I0 =>  \38174\,
                  I1 =>  \38175\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F17B\     
  \=38177\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38177\,
                  I0 =>  \38175\,
                  I1 =>  \38176\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS06/\    
  \=38190\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38190\,
                  I0 =>  \FS06\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS07/\    
  \=38191\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38191\,
                  I0 =>  \FS07\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS02A\    
  \=38201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38201\,
                  I0 =>  '0',
                  I1 =>  \38204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F02A\     
  \=38202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38202\,
                  I0 =>  \38204\,
                  I1 =>  \38203\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38203\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38203\,
                   R => SYSRESET,
                   S => '0' );

  \=38203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38203\,
                  I0 =>  \38202\,
                  I1 =>  \FS01/\,
                  I2 =>  \38205\,
                  I3 =>  '0' );

  \:38204\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38204\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38204\,
                   R => SYSRESET,
                   S => '0' );

  \=38204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38204\,
                  I0 =>  \38203\,
                  I1 =>  \38206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38205\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38205\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38205\,
                   R => SYSRESET,
                   S => '0' );

  \=38205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38205\,
                  I0 =>  \38203\,
                  I1 =>  \FS01/\,
                  I2 =>  \38207\,
                  I3 =>  '0' );

  -- Alias \FS02\     
  \=38206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38206\,
                  I0 =>  \38204\,
                  I1 =>  \38205\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F02B\     
  \=38207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38207\,
                  I0 =>  \38205\,
                  I1 =>  \38206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS03A\    
  \=38211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38211\,
                  I0 =>  '0',
                  I1 =>  \38214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F03A\     
  \=38212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38212\,
                  I0 =>  \38214\,
                  I1 =>  \38213\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38213\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38213\,
                   R => SYSRESET,
                   S => '0' );

  \=38213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38213\,
                  I0 =>  \38212\,
                  I1 =>  \F02A\,
                  I2 =>  \38215\,
                  I3 =>  '0' );

  \:38214\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38214\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38214\,
                   R => SYSRESET,
                   S => '0' );

  \=38214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38214\,
                  I0 =>  \38213\,
                  I1 =>  \38216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38215\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38215\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38215\,
                   R => SYSRESET,
                   S => '0' );

  \=38215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38215\,
                  I0 =>  \38213\,
                  I1 =>  \F02A\,
                  I2 =>  \38217\,
                  I3 =>  '0' );

  -- Alias \FS03\     
  \=38216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38216\,
                  I0 =>  \38214\,
                  I1 =>  \38215\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F03B\     
  \=38217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38217\,
                  I0 =>  \38215\,
                  I1 =>  \38216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS04A\    
  \=38221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38221\,
                  I0 =>  '0',
                  I1 =>  \38224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F04A\     
  \=38222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38222\,
                  I0 =>  \38224\,
                  I1 =>  \38223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38223\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38223\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38223\,
                   R => SYSRESET,
                   S => '0' );

  \=38223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38223\,
                  I0 =>  \38222\,
                  I1 =>  \F03A\,
                  I2 =>  \38225\,
                  I3 =>  '0' );

  \:38224\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38224\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38224\,
                   R => SYSRESET,
                   S => '0' );

  \=38224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38224\,
                  I0 =>  \38223\,
                  I1 =>  \38226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38225\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38225\,
                   R => SYSRESET,
                   S => '0' );

  \=38225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38225\,
                  I0 =>  \38223\,
                  I1 =>  \F03A\,
                  I2 =>  \38227\,
                  I3 =>  '0' );

  -- Alias \FS04\     
  \=38226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38226\,
                  I0 =>  \38224\,
                  I1 =>  \38225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F04B\     
  \=38227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38227\,
                  I0 =>  \38225\,
                  I1 =>  \38226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS05A\    
  \=38231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38231\,
                  I0 =>  '0',
                  I1 =>  \38234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F05A\     
  \=38232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38232\,
                  I0 =>  \38234\,
                  I1 =>  \38233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38233\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38233\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38233\,
                   R => SYSRESET,
                   S => '0' );

  \=38233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38233\,
                  I0 =>  \38232\,
                  I1 =>  \F04A\,
                  I2 =>  \38235\,
                  I3 =>  '0' );

  \:38234\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38234\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38234\,
                   R => SYSRESET,
                   S => '0' );

  \=38234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38234\,
                  I0 =>  \38233\,
                  I1 =>  \38236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38235\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38235\,
                   R => SYSRESET,
                   S => '0' );

  \=38235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38235\,
                  I0 =>  \38233\,
                  I1 =>  \F04A\,
                  I2 =>  \38237\,
                  I3 =>  '0' );

  -- Alias \FS05\     
  \=38236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38236\,
                  I0 =>  \38234\,
                  I1 =>  \38235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F05B\     
  \=38237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38237\,
                  I0 =>  \38235\,
                  I1 =>  \38236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT01\   
  \=38241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38241\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F06A\     
  \=38242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38242\,
                  I0 =>  \38244\,
                  I1 =>  \38243\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38243\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38243\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38243\,
                   R => SYSRESET,
                   S => '0' );

  \=38243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38243\,
                  I0 =>  \38242\,
                  I1 =>  \F05A\,
                  I2 =>  \38245\,
                  I3 =>  '0' );

  \:38244\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38244\,
                   R => SYSRESET,
                   S => '0' );

  \=38244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38244\,
                  I0 =>  \38243\,
                  I1 =>  \38246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38245\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38245\,
                   R => SYSRESET,
                   S => '0' );

  \=38245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38245\,
                  I0 =>  \38243\,
                  I1 =>  \F05A\,
                  I2 =>  \38247\,
                  I3 =>  '0' );

  -- Alias \FS06\     
  \=38246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38246\,
                  I0 =>  \38244\,
                  I1 =>  \38245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F06B\     
  \=38247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38247\,
                  I0 =>  \38245\,
                  I1 =>  \38246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT02\   
  \=38251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38251\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07A\     
  \=38252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38252\,
                  I0 =>  \38254\,
                  I1 =>  \38253\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38253\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38253\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38253\,
                   R => SYSRESET,
                   S => '0' );

  \=38253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38253\,
                  I0 =>  \38252\,
                  I1 =>  \F06A\,
                  I2 =>  \38255\,
                  I3 =>  '0' );

  \:38254\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38254\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38254\,
                   R => SYSRESET,
                   S => '0' );

  \=38254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38254\,
                  I0 =>  \38253\,
                  I1 =>  \38256\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38255\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38255\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38255\,
                   R => SYSRESET,
                   S => '0' );

  \=38255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38255\,
                  I0 =>  \38253\,
                  I1 =>  \F06A\,
                  I2 =>  \38257\,
                  I3 =>  '0' );

  -- Alias \FS07\     
  \=38256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38256\,
                  I0 =>  \38254\,
                  I1 =>  \38255\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07B\     
  \=38257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38257\,
                  I0 =>  \38255\,
                  I1 =>  \38256\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT03\   
  \=38261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38261\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38264\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F08A\     
  \=38262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38262\,
                  I0 =>  \38264\,
                  I1 =>  \38263\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38263\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38263\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38263\,
                   R => SYSRESET,
                   S => '0' );

  \=38263\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38263\,
                  I0 =>  \38262\,
                  I1 =>  \F07A\,
                  I2 =>  \38265\,
                  I3 =>  '0' );

  \:38264\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38264\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38264\,
                   R => SYSRESET,
                   S => '0' );

  \=38264\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38264\,
                  I0 =>  \38263\,
                  I1 =>  \38266\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38265\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38265\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38265\,
                   R => SYSRESET,
                   S => '0' );

  \=38265\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38265\,
                  I0 =>  \38263\,
                  I1 =>  \F07A\,
                  I2 =>  \38267\,
                  I3 =>  '0' );

  -- Alias \FS08\     
  \=38266\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38266\,
                  I0 =>  \38264\,
                  I1 =>  \38265\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F08B\     
  \=38267\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38267\,
                  I0 =>  \38265\,
                  I1 =>  \38266\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT04\   
  \=38271\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38271\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38274\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F09A\     
  \=38272\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38272\,
                  I0 =>  \38274\,
                  I1 =>  \38273\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38273\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38273\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38273\,
                   R => SYSRESET,
                   S => '0' );

  \=38273\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38273\,
                  I0 =>  \38272\,
                  I1 =>  \F08A\,
                  I2 =>  \38275\,
                  I3 =>  '0' );

  \:38274\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38274\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38274\,
                   R => SYSRESET,
                   S => '0' );

  \=38274\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38274\,
                  I0 =>  \38273\,
                  I1 =>  \38276\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38275\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38275\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38275\,
                   R => SYSRESET,
                   S => '0' );

  \=38275\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38275\,
                  I0 =>  \38273\,
                  I1 =>  \F08A\,
                  I2 =>  \38277\,
                  I3 =>  '0' );

  -- Alias \FS09\     
  \=38276\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38276\,
                  I0 =>  \38274\,
                  I1 =>  \38275\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F09B\     
  \=38277\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38277\,
                  I0 =>  \38275\,
                  I1 =>  \38276\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS08/\    
  \=38290\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38290\,
                  I0 =>  \FS08\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS07A\    
  \=38291\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38291\,
                  I0 =>  \FS07/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *************************
  -- ***                   ***
  -- ***  A1 /2 - SCALER.  ***
  -- ***                   ***
  -- *************************

  -- Alias \CHAT13\   
  \=38301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38301\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F18A\     
  \=38302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38302\,
                  I0 =>  \38304\,
                  I1 =>  \38303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38303\,
                   R => SYSRESET,
                   S => '0' );

  \=38303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38303\,
                  I0 =>  \38302\,
                  I1 =>  \F17A\,
                  I2 =>  \38305\,
                  I3 =>  '0' );

  \:38304\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38304\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38304\,
                   R => SYSRESET,
                   S => '0' );

  \=38304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38304\,
                  I0 =>  \38303\,
                  I1 =>  \38306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38305\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38305\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38305\,
                   R => SYSRESET,
                   S => '0' );

  \=38305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38305\,
                  I0 =>  \38303\,
                  I1 =>  \F17A\,
                  I2 =>  \38307\,
                  I3 =>  '0' );

  -- Alias \FS18\     
  \=38306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38306\,
                  I0 =>  \38304\,
                  I1 =>  \38305\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F18B\     
  \=38307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38307\,
                  I0 =>  \38305\,
                  I1 =>  \38306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHAT14\   
  \=38311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38311\,
                  I0 =>  \RCHAT/\,
                  I1 =>  \38314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F19A\     
  \=38312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38312\,
                  I0 =>  \38314\,
                  I1 =>  \38313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38313\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38313\,
                   R => SYSRESET,
                   S => '0' );

  \=38313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38313\,
                  I0 =>  \38312\,
                  I1 =>  \F18A\,
                  I2 =>  \38315\,
                  I3 =>  '0' );

  \:38314\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38314\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38314\,
                   R => SYSRESET,
                   S => '0' );

  \=38314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38314\,
                  I0 =>  \38313\,
                  I1 =>  \38316\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38315\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38315\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38315\,
                   R => SYSRESET,
                   S => '0' );

  \=38315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38315\,
                  I0 =>  \38313\,
                  I1 =>  \F18A\,
                  I2 =>  \38317\,
                  I3 =>  '0' );

  -- Alias \FS19\     
  \=38316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38316\,
                  I0 =>  \38314\,
                  I1 =>  \38315\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F19B\     
  \=38317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38317\,
                  I0 =>  \38315\,
                  I1 =>  \38316\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT01\   
  \=38321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38321\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F20A\     
  \=38322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38322\,
                  I0 =>  \38324\,
                  I1 =>  \38323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38323\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38323\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38323\,
                   R => SYSRESET,
                   S => '0' );

  \=38323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38323\,
                  I0 =>  \38322\,
                  I1 =>  \F19A\,
                  I2 =>  \38325\,
                  I3 =>  '0' );

  \:38324\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38324\,
                   R => SYSRESET,
                   S => '0' );

  \=38324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38324\,
                  I0 =>  \38323\,
                  I1 =>  \38326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38325\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38325\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38325\,
                   R => SYSRESET,
                   S => '0' );

  \=38325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38325\,
                  I0 =>  \38323\,
                  I1 =>  \F19A\,
                  I2 =>  \38327\,
                  I3 =>  '0' );

  -- Alias \FS20\     
  \=38326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38326\,
                  I0 =>  \38324\,
                  I1 =>  \38325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F20B\     
  \=38327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38327\,
                  I0 =>  \38325\,
                  I1 =>  \38326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT02\   
  \=38331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38331\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F21A\     
  \=38332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38332\,
                  I0 =>  \38334\,
                  I1 =>  \38333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38333\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38333\,
                   R => SYSRESET,
                   S => '0' );

  \=38333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38333\,
                  I0 =>  \38332\,
                  I1 =>  \F20A\,
                  I2 =>  \38335\,
                  I3 =>  '0' );

  \:38334\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38334\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38334\,
                   R => SYSRESET,
                   S => '0' );

  \=38334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38334\,
                  I0 =>  \38333\,
                  I1 =>  \38336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38335\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38335\,
                   R => SYSRESET,
                   S => '0' );

  \=38335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38335\,
                  I0 =>  \38333\,
                  I1 =>  \F20A\,
                  I2 =>  \38337\,
                  I3 =>  '0' );

  -- Alias \FS21\     
  \=38336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38336\,
                  I0 =>  \38334\,
                  I1 =>  \38335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F21B\     
  \=38337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38337\,
                  I0 =>  \38335\,
                  I1 =>  \38336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT03\   
  \=38341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38341\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F22A\     
  \=38342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38342\,
                  I0 =>  \38344\,
                  I1 =>  \38343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38343\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38343\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38343\,
                   R => SYSRESET,
                   S => '0' );

  \=38343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38343\,
                  I0 =>  \38342\,
                  I1 =>  \F21A\,
                  I2 =>  \38345\,
                  I3 =>  '0' );

  \:38344\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38344\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38344\,
                   R => SYSRESET,
                   S => '0' );

  \=38344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38344\,
                  I0 =>  \38343\,
                  I1 =>  \38346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38345\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38345\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38345\,
                   R => SYSRESET,
                   S => '0' );

  \=38345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38345\,
                  I0 =>  \38343\,
                  I1 =>  \F21A\,
                  I2 =>  \38347\,
                  I3 =>  '0' );

  -- Alias \FS22\     
  \=38346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38346\,
                  I0 =>  \38344\,
                  I1 =>  \38345\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F22B\     
  \=38347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38347\,
                  I0 =>  \38345\,
                  I1 =>  \38346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT04\   
  \=38351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38351\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F23A\     
  \=38352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38352\,
                  I0 =>  \38354\,
                  I1 =>  \38353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38353\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38353\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38353\,
                   R => SYSRESET,
                   S => '0' );

  \=38353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38353\,
                  I0 =>  \38352\,
                  I1 =>  \F22A\,
                  I2 =>  \38355\,
                  I3 =>  '0' );

  \:38354\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38354\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38354\,
                   R => SYSRESET,
                   S => '0' );

  \=38354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38354\,
                  I0 =>  \38353\,
                  I1 =>  \38356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38355\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38355\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38355\,
                   R => SYSRESET,
                   S => '0' );

  \=38355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38355\,
                  I0 =>  \38353\,
                  I1 =>  \F22A\,
                  I2 =>  \38357\,
                  I3 =>  '0' );

  -- Alias \FS23\     
  \=38356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38356\,
                  I0 =>  \38354\,
                  I1 =>  \38355\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F23B\     
  \=38357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38357\,
                  I0 =>  \38355\,
                  I1 =>  \38356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT05\   
  \=38361\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38361\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38364\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F24A\     
  \=38362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38362\,
                  I0 =>  \38364\,
                  I1 =>  \38363\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38363\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38363\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38363\,
                   R => SYSRESET,
                   S => '0' );

  \=38363\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38363\,
                  I0 =>  \38362\,
                  I1 =>  \F23A\,
                  I2 =>  \38365\,
                  I3 =>  '0' );

  \:38364\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38364\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38364\,
                   R => SYSRESET,
                   S => '0' );

  \=38364\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38364\,
                  I0 =>  \38363\,
                  I1 =>  \38366\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38365\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38365\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38365\,
                   R => SYSRESET,
                   S => '0' );

  \=38365\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38365\,
                  I0 =>  \38363\,
                  I1 =>  \F23A\,
                  I2 =>  \38367\,
                  I3 =>  '0' );

  -- Alias \FS24\     
  \=38366\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38366\,
                  I0 =>  \38364\,
                  I1 =>  \38365\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F24B\     
  \=38367\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38367\,
                  I0 =>  \38365\,
                  I1 =>  \38366\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT06\   
  \=38371\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38371\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38374\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F25A\     
  \=38372\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38372\,
                  I0 =>  \38374\,
                  I1 =>  \38373\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38373\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38373\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38373\,
                   R => SYSRESET,
                   S => '0' );

  \=38373\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38373\,
                  I0 =>  \38372\,
                  I1 =>  \F24A\,
                  I2 =>  \38375\,
                  I3 =>  '0' );

  \:38374\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38374\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38374\,
                   R => SYSRESET,
                   S => '0' );

  \=38374\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38374\,
                  I0 =>  \38373\,
                  I1 =>  \38376\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38375\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38375\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38375\,
                   R => SYSRESET,
                   S => '0' );

  \=38375\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38375\,
                  I0 =>  \38373\,
                  I1 =>  \F24A\,
                  I2 =>  \38377\,
                  I3 =>  '0' );

  -- Alias \FS25\     
  \=38376\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38376\,
                  I0 =>  \38374\,
                  I1 =>  \38375\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F25B\     
  \=38377\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38377\,
                  I0 =>  \38375\,
                  I1 =>  \38376\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F18AX\    
  \=38390\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38390\,
                  I0 =>  \F18A/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07A/\    
  \=38391\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38391\,
                  I0 =>  \F07A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT07\   
  \=38401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38401\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38404\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F26A\     
  \=38402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38402\,
                  I0 =>  \38404\,
                  I1 =>  \38403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38403\,
                   R => SYSRESET,
                   S => '0' );

  \=38403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38403\,
                  I0 =>  \38402\,
                  I1 =>  \F25A\,
                  I2 =>  \38405\,
                  I3 =>  '0' );

  \:38404\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38404\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38404\,
                   R => SYSRESET,
                   S => '0' );

  \=38404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38404\,
                  I0 =>  \38403\,
                  I1 =>  \38406\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38405\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38405\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38405\,
                   R => SYSRESET,
                   S => '0' );

  \=38405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38405\,
                  I0 =>  \38403\,
                  I1 =>  \F25A\,
                  I2 =>  \38407\,
                  I3 =>  '0' );

  -- Alias \FS26\     
  \=38406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38406\,
                  I0 =>  \38404\,
                  I1 =>  \38405\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F26B\     
  \=38407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38407\,
                  I0 =>  \38405\,
                  I1 =>  \38406\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT08\   
  \=38411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38411\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38414\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F27A\     
  \=38412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38412\,
                  I0 =>  \38414\,
                  I1 =>  \38413\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38413\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38413\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38413\,
                   R => SYSRESET,
                   S => '0' );

  \=38413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38413\,
                  I0 =>  \38412\,
                  I1 =>  \F26A\,
                  I2 =>  \38415\,
                  I3 =>  '0' );

  \:38414\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38414\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38414\,
                   R => SYSRESET,
                   S => '0' );

  \=38414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38414\,
                  I0 =>  \38413\,
                  I1 =>  \38416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38415\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38415\,
                   R => SYSRESET,
                   S => '0' );

  \=38415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38415\,
                  I0 =>  \38413\,
                  I1 =>  \F26A\,
                  I2 =>  \38417\,
                  I3 =>  '0' );

  -- Alias \FS27\     
  \=38416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38416\,
                  I0 =>  \38414\,
                  I1 =>  \38415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F27B\     
  \=38417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38417\,
                  I0 =>  \38415\,
                  I1 =>  \38416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT09\   
  \=38421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38421\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F28A\     
  \=38422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38422\,
                  I0 =>  \38424\,
                  I1 =>  \38423\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38423\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38423\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38423\,
                   R => SYSRESET,
                   S => '0' );

  \=38423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38423\,
                  I0 =>  \38422\,
                  I1 =>  \F27A\,
                  I2 =>  \38425\,
                  I3 =>  '0' );

  \:38424\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38424\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38424\,
                   R => SYSRESET,
                   S => '0' );

  \=38424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38424\,
                  I0 =>  \38423\,
                  I1 =>  \38426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38425\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38425\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38425\,
                   R => SYSRESET,
                   S => '0' );

  \=38425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38425\,
                  I0 =>  \38423\,
                  I1 =>  \F27A\,
                  I2 =>  \38427\,
                  I3 =>  '0' );

  -- Alias \FS28\     
  \=38426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38426\,
                  I0 =>  \38424\,
                  I1 =>  \38425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F28B\     
  \=38427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38427\,
                  I0 =>  \38425\,
                  I1 =>  \38426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT10\   
  \=38431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38431\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38434\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F29A\     
  \=38432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38432\,
                  I0 =>  \38434\,
                  I1 =>  \38433\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38433\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38433\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38433\,
                   R => SYSRESET,
                   S => '0' );

  \=38433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38433\,
                  I0 =>  \38432\,
                  I1 =>  \F28A\,
                  I2 =>  \38435\,
                  I3 =>  '0' );

  \:38434\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38434\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38434\,
                   R => SYSRESET,
                   S => '0' );

  \=38434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38434\,
                  I0 =>  \38433\,
                  I1 =>  \38436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38435\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38435\,
                   R => SYSRESET,
                   S => '0' );

  \=38435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38435\,
                  I0 =>  \38433\,
                  I1 =>  \F28A\,
                  I2 =>  \38437\,
                  I3 =>  '0' );

  -- Alias \FS29\     
  \=38436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38436\,
                  I0 =>  \38434\,
                  I1 =>  \38435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F29B\     
  \=38437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38437\,
                  I0 =>  \38435\,
                  I1 =>  \38436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT11\   
  \=38441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38441\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38444\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F30A\     
  \=38442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38442\,
                  I0 =>  \38444\,
                  I1 =>  \38443\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38443\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38443\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38443\,
                   R => SYSRESET,
                   S => '0' );

  \=38443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38443\,
                  I0 =>  \38442\,
                  I1 =>  \F29A\,
                  I2 =>  \38445\,
                  I3 =>  '0' );

  \:38444\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38444\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38444\,
                   R => SYSRESET,
                   S => '0' );

  \=38444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38444\,
                  I0 =>  \38443\,
                  I1 =>  \38446\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38445\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38445\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38445\,
                   R => SYSRESET,
                   S => '0' );

  \=38445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38445\,
                  I0 =>  \38443\,
                  I1 =>  \F29A\,
                  I2 =>  \38447\,
                  I3 =>  '0' );

  -- Alias \FS30\     
  \=38446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38446\,
                  I0 =>  \38444\,
                  I1 =>  \38445\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F30B\     
  \=38447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38447\,
                  I0 =>  \38445\,
                  I1 =>  \38446\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT12\   
  \=38451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38451\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F31A\     
  \=38452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38452\,
                  I0 =>  \38454\,
                  I1 =>  \38453\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38453\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38453\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38453\,
                   R => SYSRESET,
                   S => '0' );

  \=38453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38453\,
                  I0 =>  \38452\,
                  I1 =>  \F30A\,
                  I2 =>  \38455\,
                  I3 =>  '0' );

  \:38454\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38454\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38454\,
                   R => SYSRESET,
                   S => '0' );

  \=38454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38454\,
                  I0 =>  \38453\,
                  I1 =>  \38456\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38455\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38455\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38455\,
                   R => SYSRESET,
                   S => '0' );

  \=38455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38455\,
                  I0 =>  \38453\,
                  I1 =>  \F30A\,
                  I2 =>  \38457\,
                  I3 =>  '0' );

  -- Alias \FS31\     
  \=38456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38456\,
                  I0 =>  \38454\,
                  I1 =>  \38455\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F31B\     
  \=38457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38457\,
                  I0 =>  \38455\,
                  I1 =>  \38456\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT13\   
  \=38461\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38461\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38464\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F32A\     
  \=38462\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38462\,
                  I0 =>  \38464\,
                  I1 =>  \38463\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38463\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38463\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38463\,
                   R => SYSRESET,
                   S => '0' );

  \=38463\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38463\,
                  I0 =>  \38462\,
                  I1 =>  \F31A\,
                  I2 =>  \38465\,
                  I3 =>  '0' );

  \:38464\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38464\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38464\,
                   R => SYSRESET,
                   S => '0' );

  \=38464\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38464\,
                  I0 =>  \38463\,
                  I1 =>  \38466\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38465\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38465\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38465\,
                   R => SYSRESET,
                   S => '0' );

  \=38465\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38465\,
                  I0 =>  \38463\,
                  I1 =>  \F31A\,
                  I2 =>  \38467\,
                  I3 =>  '0' );

  -- Alias \FS32\     
  \=38466\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38466\,
                  I0 =>  \38464\,
                  I1 =>  \38465\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F32B\     
  \=38467\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38467\,
                  I0 =>  \38465\,
                  I1 =>  \38466\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHBT14\   
  \=38471\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38471\,
                  I0 =>  \RCHBT/\,
                  I1 =>  \38474\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F33A\     
  \=38472\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38472\,
                  I0 =>  \38474\,
                  I1 =>  \38473\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38473\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38473\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38473\,
                   R => SYSRESET,
                   S => '0' );

  \=38473\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38473\,
                  I0 =>  \38472\,
                  I1 =>  \F32A\,
                  I2 =>  \38475\,
                  I3 =>  '0' );

  \:38474\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38474\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38474\,
                   R => SYSRESET,
                   S => '0' );

  \=38474\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38474\,
                  I0 =>  \38473\,
                  I1 =>  \38476\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:38475\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \38475\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$38475\,
                   R => SYSRESET,
                   S => '0' );

  \=38475\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$38475\,
                  I0 =>  \38473\,
                  I1 =>  \F32A\,
                  I2 =>  \38477\,
                  I3 =>  '0' );

  -- Alias \FS33\     
  \=38476\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38476\,
                  I0 =>  \38474\,
                  I1 =>  \38475\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F33B\     
  \=38477\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38477\,
                  I0 =>  \38475\,
                  I1 =>  \38476\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F18A/\    
  \=38490\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38490\,
                  I0 =>  \F18A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F03B/\    
  \=38491\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \38491\,
                  I0 =>  '0',
                  I1 =>  \F03B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ************************
  -- ***                  ***
  -- ***  A2 /1 - TIMER.  ***
  -- ***                  ***
  -- ************************

  \=37101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37101\,
                  I0 =>  \37105\,
                  I1 =>  \37102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37102\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37102\,
                   R => SYSRESET,
                   S => '0' );

  \=37102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37102\,
                  I0 =>  \37101\,
                  I1 =>  \CLOCK\,
                  I2 =>  \37103\,
                  I3 =>  '0' );

  \:37103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37103\,
                   R => '0',
                   S => SYSRESET );

  \=37103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37103\,
                  I0 =>  \37102\,
                  I1 =>  \CLOCK\,
                  I2 =>  \37104\,
                  I3 =>  '0' );

  -- Alias \PHS2\     
  \=37104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37104\,
                  I0 =>  \37103\,
                  I1 =>  \37106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37105\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37105\,
                   R => '0',
                   S => SYSRESET );

  \=37105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37105\,
                  I0 =>  \37102\,
                  I1 =>  \37106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37106\,
                  I0 =>  \37105\,
                  I1 =>  \37103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37107\,
                  I0 =>  \37101\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PHS4\     
  \=37108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37108\,
                  I0 =>  \37107\,
                  I1 =>  \37103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PHS4/\    
  \=37109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37109\,
                  I0 =>  \37108\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37111\,
                  I0 =>  \37117\,
                  I1 =>  \37112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37112\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37112\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37112\,
                   R => SYSRESET,
                   S => '0' );

  \=37112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37112\,
                  I0 =>  \37111\,
                  I1 =>  \37107\,
                  I2 =>  \37113\,
                  I3 =>  '0' );

  \:37113\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37113\,
                   R => SYSRESET,
                   S => '0' );

  \=37113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37113\,
                  I0 =>  \37112\,
                  I1 =>  \37107\,
                  I2 =>  \37114\,
                  I3 =>  '0' );

  \=37114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37114\,
                  I0 =>  \37113\,
                  I1 =>  \37118\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RINGA/\   
  \=37115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37115\,
                  I0 =>  \37111\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37117\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37117\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37117\,
                   R => '0',
                   S => SYSRESET );

  \=37117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37117\,
                  I0 =>  \37112\,
                  I1 =>  \37118\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37118\,
                  I0 =>  \37117\,
                  I1 =>  \37113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RINGB/\   
  \=37119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37119\,
                  I0 =>  \37114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37121\,
                  I0 =>  \STOP\,
                  I1 =>  \37115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ODDSET/\  
  \=37122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37122\,
                  I0 =>  \37121\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EVNSET\   
  \=37125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37125\,
                  I0 =>  \37119\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EVNSET/\  
  \=37126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37126\,
                  I0 =>  \37125\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RT\       
  \=37129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37129\,
                  I0 =>  \37103\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WT\       
  \=37130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37130\,
                  I0 =>  \37105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WT/\      
  \=37131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37131\,
                  I0 =>  \37130\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TT/\      
  \=37135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37135\,
                  I0 =>  \37130\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MONWT\    
  \=37136\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37136\,
                  I0 =>  \37131\,
                  I1 =>  \37131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CLK\      
  \=37137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37137\,
                  I0 =>  \37131\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Q2A\      
  \=37138\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37138\,
                  I0 =>  \37131\,
                  I1 =>  \37131\,
                  I2 =>  \37131\,
                  I3 =>  '0' );

  \=37139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37139\,
                  I0 =>  \37102\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CT\       
  \=37140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37140\,
                  I0 =>  \37139\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CT/\      
  \=37142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37142\,
                  I0 =>  \37140\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37148\,
                  I0 =>  \37142\,
                  I1 =>  \37149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37149\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37149\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37149\,
                   R => SYSRESET,
                   S => '0' );

  \=37149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37149\,
                  I0 =>  \37154\,
                  I1 =>  \37148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37150\,
                  I0 =>  \37152\,
                  I1 =>  \37149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OVFSTB/\  
  \=37151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37151\,
                  I0 =>  \37149\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37152\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37152\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37152\,
                   R => '0',
                   S => SYSRESET );

  \=37152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37152\,
                  I0 =>  \37150\,
                  I1 =>  \37148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37153\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37153\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37153\,
                   R => SYSRESET,
                   S => '0' );

  \=37153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37153\,
                  I0 =>  \37152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37154\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37154\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37154\,
                   R => '0',
                   S => SYSRESET );

  \=37154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37154\,
                  I0 =>  \37153\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PHS2/\    
  \=37155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37155\,
                  I0 =>  \37104\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ************************
  -- ***                  ***
  -- ***  A2 /2 - TIMER.  ***
  -- ***                  ***
  -- ************************

  \=37201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37201\,
                  I0 =>  \RINGB/\,
                  I1 =>  \37220\,
                  I2 =>  \37216\,
                  I3 =>  '0' );

  \=37202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37202\,
                  I0 =>  \37215\,
                  I1 =>  \37219\,
                  I2 =>  \RINGA/\,
                  I3 =>  '0' );

  -- Alias \P01\      
  \:37203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37203\,
                   R => '0',
                   S => SYSRESET );

  \=37203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37203\,
                  I0 =>  \37201\,
                  I1 =>  \37204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P01/\     
  \=37204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37204\,
                  I0 =>  \37203\,
                  I1 =>  \37202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37205\,
                  I0 =>  \RINGA/\,
                  I1 =>  \37203\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37206\,
                  I0 =>  \37204\,
                  I1 =>  \RINGB/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P02\      
  \:37207\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37207\,
                   R => SYSRESET,
                   S => '0' );

  \=37207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37207\,
                  I0 =>  \37205\,
                  I1 =>  \37208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P02/\     
  \=37208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37208\,
                  I0 =>  \37207\,
                  I1 =>  \37206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37209\,
                  I0 =>  \RINGB/\,
                  I1 =>  \37207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37210\,
                  I0 =>  \37208\,
                  I1 =>  \RINGA/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P03\      
  \:37211\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37211\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37211\,
                   R => SYSRESET,
                   S => '0' );

  \=37211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37211\,
                  I0 =>  \37209\,
                  I1 =>  \37212\,
                  I2 =>  '0',
                  I3 => \&39261\ );

  -- Alias \P03/\     
  \=37212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37212\,
                  I0 =>  \37211\,
                  I1 =>  \37210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37213\,
                  I0 =>  \RINGA/\,
                  I1 =>  \37211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37214\,
                  I0 =>  \37212\,
                  I1 =>  \RINGB/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P04\      
  \:37215\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37215\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37215\,
                   R => SYSRESET,
                   S => '0' );

  \=37215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37215\,
                  I0 =>  \37213\,
                  I1 =>  \37216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P04/\     
  \=37216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37216\,
                  I0 =>  \37215\,
                  I1 =>  \37214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37217\,
                  I0 =>  \RINGB/\,
                  I1 =>  \37215\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37218\,
                  I0 =>  \37216\,
                  I1 =>  \RINGA/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P05\      
  \:37219\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37219\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37219\,
                   R => SYSRESET,
                   S => '0' );

  \=37219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37219\,
                  I0 =>  \37217\,
                  I1 =>  \37220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P05/\     
  \=37220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37220\,
                  I0 =>  \37219\,
                  I1 =>  \37218\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F01D\     
  \=37221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37221\,
                  I0 =>  \37225\,
                  I1 =>  \37222\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F01B\     
  \:37222\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37222\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37222\,
                   R => SYSRESET,
                   S => '0' );

  \=37222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37222\,
                  I0 =>  \37221\,
                  I1 =>  \P01/\,
                  I2 =>  \37223\,
                  I3 =>  '0' );

  -- Alias \F01A\     
  \:37223\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37223\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37223\,
                   R => '0',
                   S => SYSRESET );

  \=37223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37223\,
                  I0 =>  \37222\,
                  I1 =>  \P01/\,
                  I2 =>  \37224\,
                  I3 =>  '0' );

  -- Alias \F01C\     
  \=37224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37224\,
                  I0 =>  \37223\,
                  I1 =>  \37226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS01/\    
  \:37225\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37225\,
                   R => '0',
                   S => SYSRESET );

  \=37225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37225\,
                  I0 =>  \37222\,
                  I1 =>  \37226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS01\     
  \=37226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37226\,
                  I0 =>  \37225\,
                  I1 =>  \37223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \37228\    
  \=37227\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37227\,
                  I0 =>  \SBY\,
                  I1 =>  \ALGA\,
                  I2 =>  \MSTRTP\,
                  I3 =>  '0' );

  -- Alias \GOSET/\   
  \:37228\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37228\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37228\,
                   R => '0',
                   S => SYSRESET );

  \=37228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37228\,
                  I0 =>  \STRT1\,
                  I1 =>  \STRT2\,
                  I2 =>  \37229\,
                  I3 => \&37227\ );

  \=37229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37229\,
                  I0 =>  \37228\,
                  I1 =>  \GOJ1\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37230\,
                  I0 =>  \37228\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37231\,
                  I0 =>  \T12DC/\,
                  I1 =>  \37228\,
                  I2 =>  \EVNSET/\,
                  I3 =>  '0' );

  \=37232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37232\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37233\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37233\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37233\,
                   R => '0',
                   S => SYSRESET );

  \=37233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37233\,
                  I0 =>  \37231\,
                  I1 =>  \37234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STOPA\    
  \=37234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37234\,
                  I0 =>  \37233\,
                  I1 =>  \37232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37235\,
                  I0 =>  \MSTP\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37236\,
                  I0 =>  \T12DC/\,
                  I1 =>  \37235\,
                  I2 =>  \EVNSET/\,
                  I3 =>  '0' );

  \=37237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37237\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \MSTP\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37238\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37238\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37238\,
                   R => '0',
                   S => SYSRESET );

  \=37238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37238\,
                  I0 =>  \37236\,
                  I1 =>  \37239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37239\,
                  I0 =>  \37238\,
                  I1 =>  \37237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GOJAM/\   
  \=37240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37240\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 => \&37241\ );

  -- Alias \37240\    
  \=37241\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37241\,
                  I0 =>  \37234\,
                  I1 =>  \37234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STOP/\    
  \=37242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37242\,
                  I0 =>  \37234\,
                  I1 =>  \37239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STOP\     
  \=37243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37243\,
                  I0 =>  \37242\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSTPIT/\  
  \=37244\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37244\,
                  I0 =>  \37243\,
                  I1 =>  \37243\,
                  I2 =>  \37243\,
                  I3 =>  '0' );

  -- Alias \GOJAM\    
  \=37245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37245\,
                  I0 =>  \37240\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MGOJAM\   
  \=37251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37251\,
                  I0 =>  \37240\,
                  I1 =>  \37240\,
                  I2 =>  \37240\,
                  I3 =>  '0' );

  -- Alias \SB0\      
  \=37255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37255\,
                  I0 =>  \P02/\,
                  I1 =>  \P05\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB1\      
  \=37256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37256\,
                  I0 =>  \P05/\,
                  I1 =>  \P03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB2\      
  \=37257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37257\,
                  I0 =>  \P05/\,
                  I1 =>  \P02\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB4\      
  \=37258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37258\,
                  I0 =>  \P02/\,
                  I1 =>  \P04\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EDSET\    
  \=37259\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37259\,
                  I0 =>  \P02\,
                  I1 =>  \P03/\,
                  I2 =>  \P04\,
                  I3 =>  '0' );

  -- ************************
  -- ***                  ***
  -- ***  A2 /3 - TIMER.  ***
  -- ***                  ***
  -- ************************

  -- Alias \T12\      
  \=37301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37301\,
                  I0 =>  \37302\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T12DC/\   
  \=37302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37302\,
                  I0 =>  \37355\,
                  I1 =>  \GOJAM\,
                  I2 =>  \37303\,
                  I3 =>  '0' );

  \:37303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37303\,
                   R => '0',
                   S => SYSRESET );

  \=37303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37303\,
                  I0 =>  \37302\,
                  I1 =>  \37306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37304\,
                  I0 =>  \37302\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T01DC/\   
  \:37305\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37305\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37305\,
                   R => '0',
                   S => SYSRESET );

  \=37305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37305\,
                  I0 =>  \37304\,
                  I1 =>  \37306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37306\,
                  I0 =>  \37305\,
                  I1 =>  \37310\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \T01\      
  \=37307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37307\,
                  I0 =>  \37305\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37308\,
                  I0 =>  \37305\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T02DC/\   
  \:37309\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37309\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37309\,
                   R => '0',
                   S => SYSRESET );

  \=37309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37309\,
                  I0 =>  \37308\,
                  I1 =>  \37310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37310\,
                  I0 =>  \37309\,
                  I1 =>  \37314\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \T02\      
  \=37311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37311\,
                  I0 =>  \37309\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37312\,
                  I0 =>  \37309\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T03DC/\   
  \:37313\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37313\,
                   R => '0',
                   S => SYSRESET );

  \=37313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37313\,
                  I0 =>  \37312\,
                  I1 =>  \37314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37314\,
                  I0 =>  \37313\,
                  I1 =>  \37318\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \T03\      
  \=37315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37315\,
                  I0 =>  \37313\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37316\,
                  I0 =>  \37313\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37317\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37317\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37317\,
                   R => '0',
                   S => SYSRESET );

  \=37317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37317\,
                  I0 =>  \37316\,
                  I1 =>  \37318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37318\,
                  I0 =>  \37317\,
                  I1 =>  \37322\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \T04\      
  \=37319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37319\,
                  I0 =>  \37317\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37320\,
                  I0 =>  \37317\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37321\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37321\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37321\,
                   R => '0',
                   S => SYSRESET );

  \=37321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37321\,
                  I0 =>  \37320\,
                  I1 =>  \37322\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37322\,
                  I0 =>  \37321\,
                  I1 =>  \37327\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \T05\      
  \=37323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37323\,
                  I0 =>  \37321\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37325\,
                  I0 =>  \37321\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T06DC/\   
  \:37326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37326\,
                   R => '0',
                   S => SYSRESET );

  \=37326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37326\,
                  I0 =>  \37327\,
                  I1 =>  \37325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37327\,
                  I0 =>  \GOJAM\,
                  I1 =>  \37331\,
                  I2 =>  \37326\,
                  I3 =>  '0' );

  -- Alias \T06\      
  \=37328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37328\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37329\,
                  I0 =>  \ODDSET/\,
                  I1 =>  \37326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T07DC/\   
  \:37330\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37330\,
                   R => '0',
                   S => SYSRESET );

  \=37330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37330\,
                  I0 =>  \37331\,
                  I1 =>  \37329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37331\,
                  I0 =>  \GOJAM\,
                  I1 =>  \37335\,
                  I2 =>  \37330\,
                  I3 =>  '0' );

  -- Alias \T07\      
  \=37332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37332\,
                  I0 =>  \ODDSET/\,
                  I1 =>  \37330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37333\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T08DC/\   
  \:37334\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37334\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37334\,
                   R => '0',
                   S => SYSRESET );

  \=37334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37334\,
                  I0 =>  \37335\,
                  I1 =>  \37333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37335\,
                  I0 =>  \GOJAM\,
                  I1 =>  \37339\,
                  I2 =>  \37334\,
                  I3 =>  '0' );

  -- Alias \T08\      
  \=37336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37336\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37337\,
                  I0 =>  \ODDSET/\,
                  I1 =>  \37334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T09DC/\   
  \:37338\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37338\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37338\,
                   R => '0',
                   S => SYSRESET );

  \=37338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37338\,
                  I0 =>  \37339\,
                  I1 =>  \37337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37339\,
                  I0 =>  \37343\,
                  I1 =>  \GOJAM\,
                  I2 =>  \37338\,
                  I3 =>  '0' );

  -- Alias \T09\      
  \=37340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37340\,
                  I0 =>  \ODDSET/\,
                  I1 =>  \37338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37341\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T10DC/\   
  \:37342\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37342\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37342\,
                   R => '0',
                   S => SYSRESET );

  \=37342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37342\,
                  I0 =>  \37343\,
                  I1 =>  \37341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37343\,
                  I0 =>  \37348\,
                  I1 =>  \GOJAM\,
                  I2 =>  \37342\,
                  I3 =>  '0' );

  -- Alias \T10\      
  \=37344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37344\,
                  I0 =>  \37342\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37345\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37345\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37345\,
                   R => SYSRESET,
                   S => '0' );

  \=37345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37345\,
                  I0 =>  \37342\,
                  I1 =>  \ODDSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37346\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \37346\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37346\,
                   R => SYSRESET,
                   S => '0' );

  \=37346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37346\,
                  I0 =>  \37343\,
                  I1 =>  \EVNSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:37347\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \37347\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$37347\,
                   R => '0',
                   S => SYSRESET );

  \=37347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$37347\,
                  I0 =>  \37348\,
                  I1 =>  \37345\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=37348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37348\,
                  I0 =>  \GOJAM\,
                  I1 =>  \37346\,
                  I2 =>  \37347\,
                  I3 =>  '0' );

  -- Alias \T11\      
  \=37349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37349\,
                  I0 =>  \ODDSET/\,
                  I1 =>  \37347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RT/\      
  \=37350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37350\,
                  I0 =>  \RT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OVF\      
  \=37353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37353\,
                  I0 =>  \WL15/\,
                  I1 =>  \WL16\,
                  I2 =>  \OVFSTB/\,
                  I3 =>  '0' );

  -- Alias \UNF\      
  \=37354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37354\,
                  I0 =>  \OVFSTB/\,
                  I1 =>  \WL15\,
                  I2 =>  \WL16/\,
                  I3 =>  '0' );

  -- Alias \T12SET\   
  \=37355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37355\,
                  I0 =>  \EVNSET/\,
                  I1 =>  \37339\,
                  I2 =>  \37343\,
                  I3 => \&37356\ );

  -- Alias \37355\    
  \=37356\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37356\,
                  I0 =>  \37327\,
                  I1 =>  \37331\,
                  I2 =>  \37335\,
                  I3 => \&37357\ );

  -- Alias \37355\    
  \=37357\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37357\,
                  I0 =>  \37322\,
                  I1 =>  \37318\,
                  I2 =>  \37314\,
                  I3 => \&37358\ );

  -- Alias \37355\    
  \=37358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37358\,
                  I0 =>  \37310\,
                  I1 =>  \37306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CINORM\   
  \=37360\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37360\,
                  I0 =>  \MP3A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T01/\     
  \=37401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37401\,
                  I0 =>  \T01\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT01\     
  \=37404\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37404\,
                  I0 =>  \37401\,
                  I1 =>  \37401\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T02/\     
  \=37405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37405\,
                  I0 =>  \T02\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT02\     
  \=37407\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37407\,
                  I0 =>  \37405\,
                  I1 =>  \37405\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T03/\     
  \=37408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37408\,
                  I0 =>  \T03\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT03\     
  \=37411\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37411\,
                  I0 =>  \37408\,
                  I1 =>  \37408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T04/\     
  \=37412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37412\,
                  I0 =>  \T04\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT04\     
  \=37415\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37415\,
                  I0 =>  \37412\,
                  I1 =>  \37412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T05/\     
  \=37416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37416\,
                  I0 =>  \T05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT05\     
  \=37422\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37422\,
                  I0 =>  \37416\,
                  I1 =>  \37416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T06/\     
  \=37423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37423\,
                  I0 =>  \T06\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT06\     
  \=37427\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37427\,
                  I0 =>  \37423\,
                  I1 =>  \37423\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T07/\     
  \=37428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37428\,
                  I0 =>  \T07\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT07\     
  \=37432\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37432\,
                  I0 =>  \37428\,
                  I1 =>  \37428\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T08/\     
  \=37433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37433\,
                  I0 =>  \T08\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT08\     
  \=37437\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37437\,
                  I0 =>  \37433\,
                  I1 =>  \37433\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T09/\     
  \=37438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37438\,
                  I0 =>  \T09\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT09\     
  \=37442\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37442\,
                  I0 =>  \37438\,
                  I1 =>  \37438\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T10/\     
  \=37443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37443\,
                  I0 =>  \T10\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT10\     
  \=37447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37447\,
                  I0 =>  \37443\,
                  I1 =>  \37443\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T11/\     
  \=37448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37448\,
                  I0 =>  \T11\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT11\     
  \=37450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37450\,
                  I0 =>  \37448\,
                  I1 =>  \37448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T12/\     
  \=37451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37451\,
                  I0 =>  \T12\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MT12\     
  \=37454\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&37454\,
                  I0 =>  \37451\,
                  I1 =>  \37451\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OVF/\     
  \=37455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37455\,
                  I0 =>  \37353\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \UNF/\     
  \=37456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \37456\,
                  I0 =>  \37354\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *******************************************
  -- ***                                     ***
  -- ***  A3 /1 - SQ REGISTER AND DECODING.  ***
  -- ***                                     ***
  -- *******************************************

  \:30001\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30001\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30001\,
                   R => '0',
                   S => SYSRESET );

  \=30001\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30001\,
                  I0 =>  \NISQ\,
                  I1 =>  \30002\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30002\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30002\,
                  I0 =>  \30001\,
                  I1 =>  \INKBT1\,
                  I2 =>  \30107\,
                  I3 =>  '0' );

  \=30003\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30003\,
                  I0 =>  \T12/\,
                  I1 =>  \30001\,
                  I2 =>  \30127\,
                  I3 =>  '0' );

  -- Alias \NISQL/\   
  \=30004\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30004\,
                  I0 =>  \30002\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30005\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30005\,
                  I0 =>  \30107\,
                  I1 =>  \30003\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30006\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30006\,
                  I0 =>  \30003\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CSQG\     
  \=30007\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30007\,
                  I0 =>  \T12/\,
                  I1 =>  \30005\,
                  I2 =>  \CT/\,
                  I3 =>  '0' );

  -- Alias \RBSQ\     
  \=30009\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30009\,
                  I0 =>  \RT/\,
                  I1 =>  \30006\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30010\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30010\,
                  I0 =>  \30006\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WSQG/\    
  \=30011\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30011\,
                  I0 =>  \30010\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30013\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30013\,
                  I0 =>  \WL16/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30014\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30014\,
                  I0 =>  \WL14/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30015\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30015\,
                  I0 =>  \WL13/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30016\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30016\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30016\,
                   R => '0',
                   S => SYSRESET );

  \=30016\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30016\,
                  I0 =>  \30013\,
                  I1 =>  \30017\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR16\    
  \=30017\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30017\,
                  I0 =>  \30016\,
                  I1 =>  \30127\,
                  I2 =>  \30007\,
                  I3 =>  '0' );

  \:30018\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30018\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30018\,
                   R => '0',
                   S => SYSRESET );

  \=30018\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30018\,
                  I0 =>  \30014\,
                  I1 =>  \30019\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR14\    
  \=30019\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30019\,
                  I0 =>  \30018\,
                  I1 =>  \30127\,
                  I2 =>  \30007\,
                  I3 =>  '0' );

  \:30020\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30020\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30020\,
                   R => '0',
                   S => SYSRESET );

  \=30020\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30020\,
                  I0 =>  \30015\,
                  I1 =>  \30021\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR13\    
  \=30021\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30021\,
                  I0 =>  \30020\,
                  I1 =>  \30127\,
                  I2 =>  \30007\,
                  I3 =>  '0' );

  -- Alias \MSQ16\    
  \=30022\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30022\,
                  I0 =>  \30016\,
                  I1 =>  \30016\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30023\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30023\,
                  I0 =>  \30016\,
                  I1 =>  \INKL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30024\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30024\,
                  I0 =>  \30017\,
                  I1 =>  \INKL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSQ14\    
  \=30025\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30025\,
                  I0 =>  \30018\,
                  I1 =>  \30018\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSQ13\    
  \=30028\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30028\,
                  I0 =>  \30020\,
                  I1 =>  \30020\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30031\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30031\,
                  I0 =>  \30023\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30032\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30032\,
                  I0 =>  \30024\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30034\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30034\,
                  I0 =>  \30018\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30036\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30036\,
                  I0 =>  \30020\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30037\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30037\,
                  I0 =>  \30036\,
                  I1 =>  \30034\,
                  I2 =>  \30032\,
                  I3 =>  '0' );

  \=30038\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30038\,
                  I0 =>  \30020\,
                  I1 =>  \30034\,
                  I2 =>  \30032\,
                  I3 =>  '0' );

  -- Alias \SQ5\      
  \=30039\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30039\,
                  I0 =>  \30020\,
                  I1 =>  \30034\,
                  I2 =>  \30031\,
                  I3 =>  '0' );

  \=30040\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30040\,
                  I0 =>  \30036\,
                  I1 =>  \30018\,
                  I2 =>  \30032\,
                  I3 =>  '0' );

  \=30041\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30041\,
                  I0 =>  \30020\,
                  I1 =>  \30018\,
                  I2 =>  \30032\,
                  I3 =>  '0' );

  \=30042\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30042\,
                  I0 =>  \30036\,
                  I1 =>  \30034\,
                  I2 =>  \30031\,
                  I3 =>  '0' );

  \=30043\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30043\,
                  I0 =>  \30036\,
                  I1 =>  \30031\,
                  I2 =>  \30018\,
                  I3 =>  '0' );

  \=30044\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30044\,
                  I0 =>  \30020\,
                  I1 =>  \30018\,
                  I2 =>  \30031\,
                  I3 =>  '0' );

  -- Alias \SQ0/\     
  \=30045\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30045\,
                  I0 =>  \30037\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ1/\     
  \=30048\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30048\,
                  I0 =>  \30038\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ2/\     
  \=30049\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30049\,
                  I0 =>  \30040\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ3/\     
  \=30053\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30053\,
                  I0 =>  \30041\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ4/\     
  \=30054\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30054\,
                  I0 =>  \30042\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ6/\     
  \=30055\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30055\,
                  I0 =>  \30043\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ7/\     
  \=30056\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30056\,
                  I0 =>  \30044\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CON1\     
  \=30057\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30057\,
                  I0 =>  \DBLTST\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CON2\     
  \=30058\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30058\,
                  I0 =>  \CON1\,
                  I1 =>  \FS09\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SCAS10\   
  \=30059\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30059\,
                  I0 =>  \CON2\,
                  I1 =>  \FS10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INKBT1\   
  \=30061\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30061\,
                  I0 =>  \INKL\,
                  I1 =>  \T01/\,
                  I2 =>  '0',
                  I3 => \&32257\ );

  \=30101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30101\,
                  I0 =>  \GOJAM\,
                  I1 =>  \MTCSAI\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30103\,
                   R => '0',
                   S => SYSRESET );

  \=30103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30103\,
                  I0 =>  \INHPLS\,
                  I1 =>  \30104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INHINT\   
  \=30104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30104\,
                  I0 =>  \30103\,
                  I1 =>  \RELPLS\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \IIP/\     
  \:30105\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30105\,
                   R => '0',
                   S => SYSRESET );

  \=30105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30105\,
                  I0 =>  \KRPT\,
                  I1 =>  \30106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IIP\      
  \=30106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30106\,
                  I0 =>  \30105\,
                  I1 =>  \GOJAM\,
                  I2 =>  \5XP4\,
                  I3 =>  '0' );

  -- Alias \STRTFC\   
  \=30107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30107\,
                  I0 =>  \30101\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30108\,
                  I0 =>  \30004\,
                  I1 =>  \T12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30109\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30109\,
                   R => '0',
                   S => SYSRESET );

  \=30109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30109\,
                  I0 =>  \EXTPLS\,
                  I1 =>  \EXT\,
                  I2 =>  \30110\,
                  I3 =>  '0' );

  -- Alias \FUTEXT\   
  \=30110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30110\,
                  I0 =>  \30109\,
                  I1 =>  \INKBT1\,
                  I2 =>  \30107\,
                  I3 =>  '0' );

  -- Alias \MINHL\    
  \=30111\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30111\,
                  I0 =>  \30103\,
                  I1 =>  \30103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MIIP\     
  \=30112\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30112\,
                  I0 =>  \30105\,
                  I1 =>  \30105\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30113\,
                  I0 =>  \30107\,
                  I1 =>  \30108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30114\,
                  I0 =>  \30113\,
                  I1 =>  \30109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30115\,
                  I0 =>  \30113\,
                  I1 =>  \30110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \30117\    
  \=30116\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30116\,
                  I0 =>  \30110\,
                  I1 =>  \30004\,
                  I2 =>  \T12/\,
                  I3 => \&30118\ );

  -- Alias \RPTSET\   
  \=30117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30117\,
                  I0 =>  \PHS2/\,
                  I1 =>  \RUPTOR/\,
                  I2 =>  \MNHRPT\,
                  I3 => \&30116\ );

  -- Alias \30117\    
  \=30118\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30118\,
                  I0 =>  \OVNHRP\,
                  I1 =>  \30104\,
                  I2 =>  \30106\,
                  I3 => \&40441\ );

  \:30119\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30119\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30119\,
                   R => '0',
                   S => SYSRESET );

  \=30119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30119\,
                  I0 =>  \30127\,
                  I1 =>  \30114\,
                  I2 =>  \30120\,
                  I3 =>  '0' );

  \=30120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30120\,
                  I0 =>  \30119\,
                  I1 =>  \30115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30121\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30121\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30121\,
                   R => '0',
                   S => SYSRESET );

  \=30121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30121\,
                  I0 =>  \30117\,
                  I1 =>  \30122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30122\,
                  I0 =>  \30121\,
                  I1 =>  \30107\,
                  I2 =>  \T02\,
                  I3 =>  '0' );

  -- Alias \MSQEXT\   
  \=30123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30123\,
                  I0 =>  \30119\,
                  I1 =>  \30119\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQEXT/\   
  \=30124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30124\,
                  I0 =>  \30120\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RPTFRC\   
  \=30127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30127\,
                  I0 =>  \30121\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30129\,
                  I0 =>  \WL12/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30130\,
                  I0 =>  \WL11/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30131\,
                  I0 =>  \WL10/\,
                  I1 =>  \30011\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30132\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30132\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30132\,
                   R => '0',
                   S => SYSRESET );

  \=30132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30132\,
                  I0 =>  \30127\,
                  I1 =>  \30129\,
                  I2 =>  \30133\,
                  I3 =>  '0' );

  -- Alias \SQR12\    
  \=30133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30133\,
                  I0 =>  \30132\,
                  I1 =>  \30007\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30134\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30134\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30134\,
                   R => '0',
                   S => SYSRESET );

  \=30134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30134\,
                  I0 =>  \30127\,
                  I1 =>  \30130\,
                  I2 =>  \30135\,
                  I3 =>  '0' );

  -- Alias \SQR11\    
  \=30135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30135\,
                  I0 =>  \30134\,
                  I1 =>  \30007\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:30136\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \30136\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$30136\,
                   R => '0',
                   S => SYSRESET );

  \=30136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$30136\,
                  I0 =>  \30127\,
                  I1 =>  \30131\,
                  I2 =>  \30137\,
                  I3 =>  '0' );

  \=30137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30137\,
                  I0 =>  \30136\,
                  I1 =>  \30007\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSQ12\    
  \=30138\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30138\,
                  I0 =>  \30132\,
                  I1 =>  \30132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSQ11\    
  \=30139\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30139\,
                  I0 =>  \30134\,
                  I1 =>  \30134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSQ10\    
  \=30140\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30140\,
                  I0 =>  \30136\,
                  I1 =>  \30136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \QC0\      
  \=30141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30141\,
                  I0 =>  \30135\,
                  I1 =>  \30133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30142\,
                  I0 =>  \30134\,
                  I1 =>  \30133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30143\,
                  I0 =>  \30135\,
                  I1 =>  \30132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30144\,
                  I0 =>  \30132\,
                  I1 =>  \30134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \QC0/\     
  \=30145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30145\,
                  I0 =>  \30141\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \QC1/\     
  \=30148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30148\,
                  I0 =>  \30142\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \QC2/\     
  \=30151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30151\,
                  I0 =>  \30143\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \QC3/\     
  \=30152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30152\,
                  I0 =>  \30144\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR10\    
  \=30154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30154\,
                  I0 =>  \30136\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR10/\   
  \=30156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30156\,
                  I0 =>  \30137\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQR12/\   
  \=30157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30157\,
                  I0 =>  \30133\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQEXT\    
  \=30160\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30160\,
                  I0 =>  \30119\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *******************************************
  -- ***                                     ***
  -- ***  A3 /2 - SQ REGISTER AND DECODING.  ***
  -- ***                                     ***
  -- *******************************************

  \=30301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30301\,
                  I0 =>  \30310\,
                  I1 =>  \QC0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30302\,
                  I0 =>  \30310\,
                  I1 =>  \SQEXT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ5QC0/\  
  \=30303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30303\,
                  I0 =>  \30301\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30304\,
                  I0 =>  \30301\,
                  I1 =>  \30302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC1\      
  \=30305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30305\,
                  I0 =>  \30304\,
                  I1 =>  \ST0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC2\      
  \=30306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30306\,
                  I0 =>  \30304\,
                  I1 =>  \ST1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC2/\     
  \=30309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30309\,
                  I0 =>  \30306\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SQ5/\     
  \=30310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30310\,
                  I0 =>  \SQ5\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC11\     
  \=30313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30313\,
                  I0 =>  \SQ6/\,
                  I1 =>  \30360\,
                  I2 =>  \ST0/\,
                  I3 =>  '0' );

  \=30314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30314\,
                  I0 =>  \SQEXT/\,
                  I1 =>  \ST1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30315\,
                  I0 =>  \30314\,
                  I1 =>  \NEXST0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EXST1/\   
  \=30316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30316\,
                  I0 =>  \30314\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC6\      
  \=30317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30317\,
                  I0 =>  \30315\,
                  I1 =>  \SQ3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC7\      
  \=30318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30318\,
                  I0 =>  \30315\,
                  I1 =>  \SQ4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TC0\      
  \=30319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30319\,
                  I0 =>  \SQ0/\,
                  I1 =>  \NEXST0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TCF0\     
  \=30320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30320\,
                  I0 =>  \SQ1/\,
                  I1 =>  \NEXST0/\,
                  I2 =>  \QC0\,
                  I3 =>  '0' );

  -- Alias \NEXST0\   
  \=30321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30321\,
                  I0 =>  \SQEXT\,
                  I1 =>  \ST0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TC0/\     
  \=30322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30322\,
                  I0 =>  \30319\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC3/\     
  \=30323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30323\,
                  I0 =>  \30319\,
                  I1 =>  \STD2\,
                  I2 =>  \30320\,
                  I3 =>  '0' );

  -- Alias \NEXST0/\  
  \=30324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30324\,
                  I0 =>  \30321\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC3\      
  \=30326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30326\,
                  I0 =>  \30323\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DCS0\     
  \=30327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30327\,
                  I0 =>  \SQ4/\,
                  I1 =>  \30349\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DCA0\     
  \=30328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30328\,
                  I0 =>  \30349\,
                  I1 =>  \SQ3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC4/\     
  \=30329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30329\,
                  I0 =>  \30327\,
                  I1 =>  \30328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC4\      
  \=30330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30330\,
                  I0 =>  \30329\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC13/\    
  \=30331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30331\,
                  I0 =>  \30318\,
                  I1 =>  \30317\,
                  I2 =>  \30313\,
                  I3 => \&30332\ );

  -- Alias \30331\    
  \=30332\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30332\,
                  I0 =>  \30305\,
                  I1 =>  \30327\,
                  I2 =>  \30328\,
                  I3 =>  '0' );

  -- Alias \IC13\     
  \=30333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30333\,
                  I0 =>  \30331\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30335\,
                  I0 =>  \QC1/\,
                  I1 =>  \ST1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30336\,
                  I0 =>  \QC3/\,
                  I1 =>  \ST0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30337\,
                  I0 =>  \30335\,
                  I1 =>  \30336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC5\      
  \=30338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30338\,
                  I0 =>  \30337\,
                  I1 =>  \30310\,
                  I2 =>  \SQEXT\,
                  I3 =>  '0' );

  -- Alias \IC5/\     
  \=30339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30339\,
                  I0 =>  \30338\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC9/\     
  \=30340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30340\,
                  I0 =>  \30338\,
                  I1 =>  \TS0\,
                  I2 =>  '0',
                  I3 => \&30344\ );

  -- Alias \LXCH0\    
  \=30341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30341\,
                  I0 =>  \NEXST0/\,
                  I1 =>  \QC1/\,
                  I2 =>  \SQ2/\,
                  I3 =>  '0' );

  -- Alias \QXCH0\    
  \=30342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30342\,
                  I0 =>  \SQ2/\,
                  I1 =>  \QC1/\,
                  I2 =>  \30349\,
                  I3 =>  '0' );

  -- Alias \QXCH0/\   
  \=30343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30343\,
                  I0 =>  \30342\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \30340\    
  \=30344\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30344\,
                  I0 =>  \30342\,
                  I1 =>  \30341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC9\      
  \=30345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30345\,
                  I0 =>  \30340\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC8/\     
  \=30346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30346\,
                  I0 =>  \DXCH0\,
                  I1 =>  \LXCH0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30347\,
                  I0 =>  \ST0/\,
                  I1 =>  \SQEXT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TS0\      
  \=30348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30348\,
                  I0 =>  \30310\,
                  I1 =>  \QC2/\,
                  I2 =>  \NEXST0/\,
                  I3 =>  '0' );

  -- Alias \EXST0/\   
  \=30349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30349\,
                  I0 =>  \30347\,
                  I1 =>  \30347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TS0/\     
  \=30350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30350\,
                  I0 =>  \30348\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DXCH0\    
  \=30352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30352\,
                  I0 =>  \30310\,
                  I1 =>  \NEXST0/\,
                  I2 =>  \QC1/\,
                  I3 =>  '0' );

  -- Alias \DAS0\     
  \=30354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30354\,
                  I0 =>  \SQ2/\,
                  I1 =>  \NEXST0/\,
                  I2 =>  \QC0/\,
                  I3 =>  '0' );

  -- Alias \IC10/\    
  \=30356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30356\,
                  I0 =>  \30330\,
                  I1 =>  \30352\,
                  I2 =>  \30354\,
                  I3 =>  '0' );

  -- Alias \IC10\     
  \=30357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30357\,
                  I0 =>  \30356\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30360\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30360\,
                  I0 =>  \SQEXT/\,
                  I1 =>  \QC0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DAS0/\    
  \=30401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30401\,
                  I0 =>  \DAS0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BZF0\     
  \=30403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30403\,
                  I0 =>  \SQ1/\,
                  I1 =>  \QC0\,
                  I2 =>  \EXST0/\,
                  I3 =>  '0' );

  -- Alias \BZF0/\    
  \=30404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30404\,
                  I0 =>  \30403\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMF0\     
  \=30405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30405\,
                  I0 =>  \EXST0/\,
                  I1 =>  \QC0\,
                  I2 =>  \SQ6/\,
                  I3 =>  '0' );

  -- Alias \BMF0/\    
  \=30406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30406\,
                  I0 =>  \30405\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30407\,
                  I0 =>  \BZF0/\,
                  I1 =>  \BR2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30408\,
                  I0 =>  \BMF0/\,
                  I1 =>  \BR1B2B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC16/\    
  \=30409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30409\,
                  I0 =>  \30407\,
                  I1 =>  \30408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC15/\    
  \=30410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30410\,
                  I0 =>  \30405\,
                  I1 =>  \30403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC16\     
  \=30411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30411\,
                  I0 =>  \30409\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC17\     
  \=30412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30412\,
                  I0 =>  \30411\,
                  I1 =>  \30410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC15\     
  \=30413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30413\,
                  I0 =>  \30410\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCS0\     
  \=30415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30415\,
                  I0 =>  \SQ1/\,
                  I1 =>  \QC0/\,
                  I2 =>  \30324\,
                  I3 =>  '0' );

  -- Alias \CCS0/\    
  \=30416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30416\,
                  I0 =>  \30415\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30417\,
                  I0 =>  \SQ2/\,
                  I1 =>  \QC0/\,
                  I2 =>  '0',
                  I3 => \&30418\ );

  -- Alias \30417\    
  \=30418\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30418\,
                  I0 =>  \SQEXT\,
                  I1 =>  \ST1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DAS1/\    
  \=30419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30419\,
                  I0 =>  \30417\,
                  I1 =>  \30424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DAS1\     
  \=30421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30421\,
                  I0 =>  \30419\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC12/\    
  \=30422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30422\,
                  I0 =>  \30415\,
                  I1 =>  \30426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC12\     
  \=30423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30423\,
                  I0 =>  \30422\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ADS0\     
  \=30424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30424\,
                  I0 =>  \SQ2/\,
                  I1 =>  \QC3/\,
                  I2 =>  \30324\,
                  I3 =>  '0' );

  -- Alias \INCR0\    
  \=30425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30425\,
                  I0 =>  \QC2/\,
                  I1 =>  \SQ2/\,
                  I2 =>  \30324\,
                  I3 =>  '0' );

  -- Alias \MSU0\     
  \=30426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30426\,
                  I0 =>  \SQ2/\,
                  I1 =>  \EXST0/\,
                  I2 =>  \QC0/\,
                  I3 =>  '0' );

  -- Alias \MSU0/\    
  \=30427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30427\,
                  I0 =>  \30426\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \AUG0\     
  \=30428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30428\,
                  I0 =>  \SQ2/\,
                  I1 =>  \EXST0/\,
                  I2 =>  \QC2/\,
                  I3 =>  '0' );

  -- Alias \AUG0/\    
  \=30429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30429\,
                  I0 =>  \30428\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DIM0\     
  \=30430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30430\,
                  I0 =>  \SQ2/\,
                  I1 =>  \EXST0/\,
                  I2 =>  \QC3/\,
                  I3 =>  '0' );

  -- Alias \DIM0/\    
  \=30431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30431\,
                  I0 =>  \30430\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP3\      
  \=30432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30432\,
                  I0 =>  \ST3/\,
                  I1 =>  \SQ7/\,
                  I2 =>  \SQEXT/\,
                  I3 =>  '0' );

  -- Alias \MP3/\     
  \=30433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30433\,
                  I0 =>  \30432\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP1\      
  \=30435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30435\,
                  I0 =>  \ST1/\,
                  I1 =>  \SQEXT/\,
                  I2 =>  \SQ7/\,
                  I3 =>  '0' );

  -- Alias \MP1/\     
  \=30436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30436\,
                  I0 =>  \30435\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP0\      
  \=30437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30437\,
                  I0 =>  \ST0/\,
                  I1 =>  \SQEXT/\,
                  I2 =>  \SQ7/\,
                  I3 =>  '0' );

  -- Alias \MTCSA/\   
  \=30438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&30438\,
                  I0 =>  \TCSAJ3\,
                  I1 =>  \TCSAJ3\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP0/\     
  \=30439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30439\,
                  I0 =>  \30437\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TCSAJ3\   
  \=30441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30441\,
                  I0 =>  \SQ0/\,
                  I1 =>  \SQEXT\,
                  I2 =>  \ST3/\,
                  I3 =>  '0' );

  -- Alias \TCSAJ3/\  
  \=30442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30442\,
                  I0 =>  \30441\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSM3\     
  \=30443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30443\,
                  I0 =>  \ST3/\,
                  I1 =>  \30303\,
                  I2 =>  \SQEXT\,
                  I3 =>  '0' );

  -- Alias \RSM3/\    
  \=30444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30444\,
                  I0 =>  \30443\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SU0\      
  \=30445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30445\,
                  I0 =>  \SQ6/\,
                  I1 =>  \EXST0/\,
                  I2 =>  \QC0/\,
                  I3 =>  '0' );

  -- Alias \MASK0\    
  \=30446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30446\,
                  I0 =>  \SQ7/\,
                  I1 =>  \30324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MASK0/\   
  \=30447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30447\,
                  I0 =>  \30446\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \AD0\      
  \=30448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30448\,
                  I0 =>  \30324\,
                  I1 =>  \SQ6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NDX0\     
  \=30449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30449\,
                  I0 =>  \30324\,
                  I1 =>  \SQ5/\,
                  I2 =>  \QC0/\,
                  I3 =>  '0' );

  -- Alias \NDX0/\    
  \=30450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30450\,
                  I0 =>  \30449\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NDXX1\    
  \=30451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30451\,
                  I0 =>  \SQEXT/\,
                  I1 =>  \SQ5/\,
                  I2 =>  \ST1/\,
                  I3 =>  '0' );

  -- Alias \NDXX1/\   
  \=30452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30452\,
                  I0 =>  \30451\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GOJ1\     
  \=30453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30453\,
                  I0 =>  \SQEXT\,
                  I1 =>  \ST1/\,
                  I2 =>  \SQ0/\,
                  I3 =>  '0' );

  -- Alias \GOJ1/\    
  \=30454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30454\,
                  I0 =>  \30453\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=30455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30455\,
                  I0 =>  \30446\,
                  I1 =>  \30437\,
                  I2 =>  \RXOR0\,
                  I3 =>  '0' );

  -- Alias \IC14\     
  \=30456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \30456\,
                  I0 =>  \30455\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A4 /1 - STAGE BRANCH DECODING.  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \DIVSTG\   
  \=36101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36101\,
                  I0 =>  \36102\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T12USE/\  
  \:36102\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36102\,
                   R => '0',
                   S => SYSRESET );

  \=36102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36102\,
                  I0 =>  \DVST\,
                  I1 =>  \36109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36103\,
                  I0 =>  \T03/\,
                  I1 =>  \36102\,
                  I2 =>  \PHS3/\,
                  I3 =>  '0' );

  \=36104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36104\,
                  I0 =>  \36103\,
                  I1 =>  \36110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36105\,
                  I0 =>  \36120\,
                  I1 =>  \36151\,
                  I2 =>  \36137\,
                  I3 =>  '0' );

  -- Alias \ST0/\     
  \=36106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36106\,
                  I0 =>  \36105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP3A\     
  \=36108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36108\,
                  I0 =>  \MP3/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36109\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36109\,
                   R => SYSRESET,
                   S => '0' );

  \=36109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36109\,
                  I0 =>  \36102\,
                  I1 =>  \RSTSTG\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=36110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36110\,
                  I0 =>  \PHS3/\,
                  I1 =>  \36109\,
                  I2 =>  \T12/\,
                  I3 =>  '0' );

  -- Alias \36113\    
  \=36112\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36112\,
                  I0 =>  \GOJAM\,
                  I1 =>  \MTCSAI\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36113\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36113\,
                   R => '0',
                   S => SYSRESET );

  \=36113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36113\,
                  I0 =>  \ST1\,
                  I1 =>  \36124\,
                  I2 =>  \36118\,
                  I3 => \&36112\ );

  \=36114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36114\,
                  I0 =>  \36104\,
                  I1 =>  \36113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36115\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36115\,
                   R => '0',
                   S => SYSRESET );

  \=36115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36115\,
                  I0 =>  \36114\,
                  I1 =>  \36120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MST1\     
  \=36116\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36116\,
                  I0 =>  \36115\,
                  I1 =>  \36115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST1/\     
  \=36117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36117\,
                  I0 =>  \36121\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36118\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36118\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36118\,
                   R => SYSRESET,
                   S => '0' );

  \=36118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36118\,
                  I0 =>  \36113\,
                  I1 =>  \T01\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36119\,
                  I0 =>  \36104\,
                  I1 =>  \36118\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STG1\     
  \:36120\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36120\,
                   R => SYSRESET,
                   S => '0' );

  \=36120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36120\,
                  I0 =>  \36115\,
                  I1 =>  \36119\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST1D\     
  \=36121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36121\,
                  I0 =>  \36137\,
                  I1 =>  \36151\,
                  I2 =>  \36115\,
                  I3 =>  '0' );

  \=36124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36124\,
                  I0 =>  \36151\,
                  I1 =>  \DVST/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MST2\     
  \=36125\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36125\,
                  I0 =>  \36132\,
                  I1 =>  \36132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST1376/\  
  \=36126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36126\,
                  I0 =>  \36121\,
                  I1 =>  \36153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV1376\   
  \=36127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36127\,
                  I0 =>  \36126\,
                  I1 =>  \36202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV1376/\  
  \=36128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36128\,
                  I0 =>  \36127\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36130\    
  \=36129\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36129\,
                  I0 =>  \ST2\,
                  I1 =>  \36142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36130\,
                   R => '0',
                   S => SYSRESET );

  \=36130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36130\,
                  I0 =>  \36139\,
                  I1 =>  \MTCSAI\,
                  I2 =>  \36135\,
                  I3 => \&36129\ );

  \=36131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36131\,
                  I0 =>  \36104\,
                  I1 =>  \36130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36132\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36132\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36132\,
                   R => '0',
                   S => SYSRESET );

  \=36132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36132\,
                  I0 =>  \36131\,
                  I1 =>  \36137\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36138\    
  \=36134\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36134\,
                  I0 =>  \INKL\,
                  I1 =>  \36120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36135\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36135\,
                   R => SYSRESET,
                   S => '0' );

  \=36135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36135\,
                  I0 =>  \36130\,
                  I1 =>  \GOJAM\,
                  I2 =>  \T01\,
                  I3 =>  '0' );

  \=36136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36136\,
                  I0 =>  \36135\,
                  I1 =>  \36104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STG2\     
  \:36137\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36137\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36137\,
                   R => SYSRESET,
                   S => '0' );

  \=36137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36137\,
                  I0 =>  \36132\,
                  I1 =>  \36136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STD2\     
  \=36138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36138\,
                  I0 =>  \36151\,
                  I1 =>  \36132\,
                  I2 =>  '0',
                  I3 => \&36134\ );

  \=36139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36139\,
                  I0 =>  \DVST/\,
                  I1 =>  \36115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36140\,
                  I0 =>  \36151\,
                  I1 =>  \36132\,
                  I2 =>  \36115\,
                  I3 =>  '0' );

  -- Alias \ST3/\     
  \=36141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36141\,
                  I0 =>  \36140\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36142\,
                  I0 =>  \TRSM/\,
                  I1 =>  \XT1/\,
                  I2 =>  \XB7/\,
                  I3 => \&36161\ );

  -- Alias \MST3\     
  \=36143\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36143\,
                  I0 =>  \36148\,
                  I1 =>  \36148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36144\,
                  I0 =>  \36148\,
                  I1 =>  \36120\,
                  I2 =>  \36137\,
                  I3 =>  '0' );

  -- Alias \ST4/\     
  \=36145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36145\,
                  I0 =>  \36144\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36146\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36146\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36146\,
                   R => '0',
                   S => SYSRESET );

  \=36146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36146\,
                  I0 =>  '0',
                  I1 =>  \36155\,
                  I2 =>  \36149\,
                  I3 =>  '0' );

  \=36147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36147\,
                  I0 =>  \36104\,
                  I1 =>  \36146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36148\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36148\,
                   R => '0',
                   S => SYSRESET );

  \=36148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36148\,
                  I0 =>  \36147\,
                  I1 =>  \36151\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36149\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36149\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36149\,
                   R => SYSRESET,
                   S => '0' );

  \=36149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36149\,
                  I0 =>  \36146\,
                  I1 =>  \STRTFC\,
                  I2 =>  \T01\,
                  I3 => \&36159\ );

  \=36150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36150\,
                  I0 =>  \36149\,
                  I1 =>  \36104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STG3\     
  \=36151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36151\,
                  I0 =>  \36148\,
                  I1 =>  \36150\,
                  I2 =>  '0',
                  I3 => \&36158\ );

  \=36152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36152\,
                  I0 =>  \36120\,
                  I1 =>  \36151\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST376\    
  \=36153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36153\,
                  I0 =>  \36132\,
                  I1 =>  \36152\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST376/\   
  \=36154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36154\,
                  I0 =>  \36153\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36155\,
                  I0 =>  \DVST/\,
                  I1 =>  \36132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36156\,
                  I0 =>  \36144\,
                  I1 =>  \36153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV3764\   
  \=36157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36157\,
                  I0 =>  \36202\,
                  I1 =>  \36156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36151\    
  \=36158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36158\,
                  I0 =>  \36150\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36149\    
  \=36159\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36159\,
                  I0 =>  \RSTSTG\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36142\    
  \=36161\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36161\,
                  I0 =>  \NDR100/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36201\,
                  I0 =>  \QC0/\,
                  I1 =>  \SQEXT/\,
                  I2 =>  \SQ1/\,
                  I3 =>  '0' );

  -- Alias \DIV/\     
  \=36202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36202\,
                  I0 =>  \36201\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV0\      
  \=36204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36204\,
                  I0 =>  \36202\,
                  I1 =>  \36106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV0/\     
  \=36205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36205\,
                  I0 =>  \36204\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV376\    
  \=36206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36206\,
                  I0 =>  \36202\,
                  I1 =>  \36154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV376/\   
  \=36207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36207\,
                  I0 =>  \36206\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV4\      
  \=36208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36208\,
                  I0 =>  \36202\,
                  I1 =>  \36145\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV1\      
  \=36209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36209\,
                  I0 =>  \36202\,
                  I1 =>  \36117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV1/\     
  \=36210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36210\,
                  I0 =>  \36209\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36213\,
                  I0 =>  \SUMB16/\,
                  I1 =>  \SUMA16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SGUM\     
  \=36214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36214\,
                  I0 =>  \SUMA16/\,
                  I1 =>  \SUMB16/\,
                  I2 =>  \TSGU/\,
                  I3 => \&36215\ );

  -- Alias \36214\    
  \=36215\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36215\,
                  I0 =>  \PHS4\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36216\,
                  I0 =>  \UNF/\,
                  I1 =>  \TOV/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36217\,
                  I0 =>  \TL15\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36218\,
                  I0 =>  \L15/\,
                  I1 =>  \36217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36222\    
  \=36219\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36219\,
                  I0 =>  \36214\,
                  I1 =>  \36216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR1\      
  \=36220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36220\,
                  I0 =>  \36222\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36221\,
                  I0 =>  \PHS4/\,
                  I1 =>  \WL16/\,
                  I2 =>  \TSGN/\,
                  I3 =>  '0' );

  \:36222\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36222\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36222\,
                   R => '0',
                   S => SYSRESET );

  \=36222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36222\,
                  I0 =>  \36218\,
                  I1 =>  \36221\,
                  I2 =>  \36228\,
                  I3 => \&36219\ );

  \=36224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36224\,
                  I0 =>  \TSGN/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36228\    
  \=36225\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36225\,
                  I0 =>  \36222\,
                  I1 =>  \36224\,
                  I2 =>  \36227\,
                  I3 =>  '0' );

  -- Alias \BR1/\     
  \=36226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36226\,
                  I0 =>  \36228\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36227\,
                  I0 =>  \36217\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:36228\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36228\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36228\,
                   R => SYSRESET,
                   S => '0' );

  \=36228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36228\,
                  I0 =>  \36230\,
                  I1 =>  \36231\,
                  I2 =>  '0',
                  I3 => \&36225\ );

  \=36230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36230\,
                  I0 =>  \TOV/\,
                  I1 =>  \PHS2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36231\,
                  I0 =>  \36213\,
                  I1 =>  \PHS3/\,
                  I2 =>  \TSGU/\,
                  I3 => \&36232\ );

  -- Alias \36231\    
  \=36232\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36232\,
                  I0 =>  \PHS4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36233\,
                  I0 =>  \GEQZRO/\,
                  I1 =>  \PHS4/\,
                  I2 =>  \TPZG/\,
                  I3 =>  '0' );

  \=36236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36236\,
                  I0 =>  \TOV/\,
                  I1 =>  \OVF/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36241\    
  \=36237\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36237\,
                  I0 =>  \36233\,
                  I1 =>  \36236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR2\      
  \=36238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36238\,
                  I0 =>  \36241\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36239\,
                  I0 =>  \TSGN2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36240\,
                  I0 =>  \WL16/\,
                  I1 =>  \PHS4/\,
                  I2 =>  \36239\,
                  I3 =>  '0' );

  \:36241\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \36241\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36241\,
                   R => '0',
                   S => SYSRESET );

  \=36241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36241\,
                  I0 =>  \36240\,
                  I1 =>  \36243\,
                  I2 =>  \36249\,
                  I3 => \&36237\ );

  \=36243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36243\,
                  I0 =>  \WL16/\,
                  I1 =>  \WL15/\,
                  I2 =>  \WL14/\,
                  I3 => \&36247\ );

  \=36244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36244\,
                  I0 =>  \36239\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36249\    
  \=36245\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36245\,
                  I0 =>  \36241\,
                  I1 =>  \36244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR2/\     
  \=36246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36246\,
                  I0 =>  \36249\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36243\    
  \=36247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36247\,
                  I0 =>  \WL13/\,
                  I1 =>  \WL12/\,
                  I2 =>  \WL11/\,
                  I3 => \&36251\ );

  \:36249\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \36249\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$36249\,
                   R => SYSRESET,
                   S => '0' );

  \=36249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$36249\,
                  I0 =>  \36230\,
                  I1 =>  \36252\,
                  I2 =>  '0',
                  I3 => \&36245\ );

  -- Alias \36243\    
  \=36251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36251\,
                  I0 =>  \WL10/\,
                  I1 =>  \WL09/\,
                  I2 =>  \WL08/\,
                  I3 => \&36253\ );

  \=36252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36252\,
                  I0 =>  \PHS3/\,
                  I1 =>  \TMZ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36243\    
  \=36253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36253\,
                  I0 =>  \WL07/\,
                  I1 =>  \WL06/\,
                  I2 =>  \WL05/\,
                  I3 => \&36254\ );

  -- Alias \36243\    
  \=36254\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36254\,
                  I0 =>  \WL04/\,
                  I1 =>  \WL03/\,
                  I2 =>  \WL02/\,
                  I3 => \&36255\ );

  -- Alias \36243\    
  \=36255\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36255\,
                  I0 =>  \WL01/\,
                  I1 =>  \TMZ/\,
                  I2 =>  \PHS4/\,
                  I3 =>  '0' );

  -- Alias \MBR1\     
  \=36260\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36260\,
                  I0 =>  \36222\,
                  I1 =>  \36222\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MBR2\     
  \=36262\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36262\,
                  I0 =>  \36241\,
                  I1 =>  \36241\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TRSM/\    
  \=36263\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36263\,
                  I0 =>  \TRSM\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DVST/\    
  \=36264\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36264\,
                  I0 =>  \DVST\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A4 /2 - STAGE BRANCH DECODING.  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \DV4/\     
  \=36301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36301\,
                  I0 =>  \DV4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36303\,
                  I0 =>  \SQ0/\,
                  I1 =>  \EXST0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36304\,
                  I0 =>  \36303\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \READ0\    
  \=36305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36305\,
                  I0 =>  \36304\,
                  I1 =>  \SQR10\,
                  I2 =>  \QC0/\,
                  I3 =>  '0' );

  -- Alias \READ0/\   
  \=36306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36306\,
                  I0 =>  \36305\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WRITE0\   
  \=36308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36308\,
                  I0 =>  \QC0/\,
                  I1 =>  \36304\,
                  I2 =>  \SQR10/\,
                  I3 =>  '0' );

  -- Alias \WRITE0/\  
  \=36309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36309\,
                  I0 =>  \36308\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RAND0\    
  \=36310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36310\,
                  I0 =>  \SQR10\,
                  I1 =>  \36304\,
                  I2 =>  \QC1/\,
                  I3 =>  '0' );

  -- Alias \WAND0\    
  \=36312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36312\,
                  I0 =>  \QC1/\,
                  I1 =>  \SQR10/\,
                  I2 =>  \36304\,
                  I3 =>  '0' );

  -- Alias \INOUT/\   
  \=36313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36313\,
                  I0 =>  \36314\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INOUT\    
  \=36314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36314\,
                  I0 =>  \EXST0/\,
                  I1 =>  \SQ0/\,
                  I2 =>  \36320\,
                  I3 =>  '0' );

  -- Alias \ROR0\     
  \=36315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36315\,
                  I0 =>  \SQR10\,
                  I1 =>  \36304\,
                  I2 =>  \QC2/\,
                  I3 =>  '0' );

  -- Alias \WOR0\     
  \=36316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36316\,
                  I0 =>  \QC2/\,
                  I1 =>  \36304\,
                  I2 =>  \SQR10/\,
                  I3 =>  '0' );

  -- Alias \WOR0/\    
  \=36317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36317\,
                  I0 =>  \36316\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RXOR0\    
  \=36318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36318\,
                  I0 =>  \SQR10\,
                  I1 =>  \36304\,
                  I2 =>  \QC3/\,
                  I3 =>  '0' );

  -- Alias \RXOR0/\   
  \=36319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36319\,
                  I0 =>  \36318\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RUPT0\    
  \=36320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36320\,
                  I0 =>  \QC3/\,
                  I1 =>  \36304\,
                  I2 =>  \SQR10/\,
                  I3 =>  '0' );

  -- Alias \RUPT0/\   
  \=36321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36321\,
                  I0 =>  \36320\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8PP4\     
  \=36322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36322\,
                  I0 =>  \36314\,
                  I1 =>  \DV4\,
                  I2 =>  \36327\,
                  I3 => \&40348\ );

  -- Alias \RUPT1\    
  \=36323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36323\,
                  I0 =>  \SQ0/\,
                  I1 =>  \EXST1/\,
                  I2 =>  \QC3/\,
                  I3 => \&36325\ );

  -- Alias \RUPT1/\   
  \=36324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36324\,
                  I0 =>  \36323\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \36323\    
  \=36325\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36325\,
                  I0 =>  \SQR10/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36326\,
                  I0 =>  \QC3/\,
                  I1 =>  \SQEXT\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PRINC\    
  \=36327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36327\,
                  I0 =>  \36326\,
                  I1 =>  \36329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36328\,
                  I0 =>  \ST0/\,
                  I1 =>  \SQR12/\,
                  I2 =>  \SQ2/\,
                  I3 =>  '0' );

  \=36329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36329\,
                  I0 =>  \36328\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RRPA\     
  \=36331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36331\,
                  I0 =>  \T03/\,
                  I1 =>  \RUPT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3XP7\     
  \=36332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36332\,
                  I0 =>  \T03/\,
                  I1 =>  \RXOR0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36333\,
                  I0 =>  \ROR0\,
                  I1 =>  \WOR0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36334\,
                  I0 =>  \36333\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=36335\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36335\,
                  I0 =>  \36334\,
                  I1 =>  \36348\,
                  I2 =>  \36343\,
                  I3 => \&36430\ );

  -- Alias \9XP1\     
  \=36336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36336\,
                  I0 =>  \T09/\,
                  I1 =>  \RUPT0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36337\,
                  I0 =>  \RAND0\,
                  I1 =>  \WAND0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36338\,
                  I0 =>  \T03/\,
                  I1 =>  \36337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=36339\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36339\,
                  I0 =>  \36338\,
                  I1 =>  \36354\,
                  I2 =>  \36340\,
                  I3 => \&36428\ );

  \=36340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36340\,
                  I0 =>  \T09/\,
                  I1 =>  \RXOR0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP28\    
  \=36341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36341\,
                  I0 =>  \DV4/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36342\,
                  I0 =>  \RUPT1\,
                  I1 =>  \IC13\,
                  I2 =>  \IC12\,
                  I3 =>  '0' );

  \=36343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36343\,
                  I0 =>  \T09/\,
                  I1 =>  \36342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP11\    
  \=36344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36344\,
                  I0 =>  \T05/\,
                  I1 =>  \INOUT/\,
                  I2 =>  \READ0\,
                  I3 => \&36346\ );

  -- Alias \WG/\      
  \=36345\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36345\,
                  I0 =>  \36336\,
                  I1 =>  \36340\,
                  I2 =>  \36354\,
                  I3 => \&36347\ );

  -- Alias \36344\    
  \=36346\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36346\,
                  I0 =>  \WRITE0\,
                  I1 =>  \RXOR0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WG/\      
  \=36347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36347\,
                  I0 =>  \36343\,
                  I1 =>  \36351\,
                  I2 =>  '0',
                  I3 => \&36411\ );

  \=36348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36348\,
                  I0 =>  \READ0/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36349\,
                  I0 =>  \WRITE0/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WCH/\     
  \=36350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36350\,
                  I0 =>  \36349\,
                  I1 =>  \7XP14\,
                  I2 =>  \36353\,
                  I3 =>  '0' );

  \=36351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36351\,
                  I0 =>  \T02/\,
                  I1 =>  \WRITE0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \2XP3\     
  \=36352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36352\,
                  I0 =>  \T02/\,
                  I1 =>  \INOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36353\,
                  I0 =>  \T05/\,
                  I1 =>  \WOR0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36354\,
                  I0 =>  \T05/\,
                  I1 =>  \RXOR0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RA/\      
  \=36355\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36355\,
                  I0 =>  \36349\,
                  I1 =>  \36354\,
                  I2 =>  \36352\,
                  I3 => \&36409\ );

  \=36360\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36360\,
                  I0 =>  \STORE1/\,
                  I1 =>  \T09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36401\,
                  I0 =>  \RUPT0\,
                  I1 =>  \RUPT1\,
                  I2 =>  \RSM3\,
                  I3 =>  '0' );

  -- Alias \R15\      
  \=36402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36402\,
                  I0 =>  \36401\,
                  I1 =>  \T01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB2\      
  \=36403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36403\,
                  I0 =>  \T01/\,
                  I1 =>  \RUPT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \1XP10\    
  \=36404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36404\,
                  I0 =>  \T01/\,
                  I1 =>  \DV0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \2PP1\     
  \=36405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36405\,
                  I0 =>  \INOUT\,
                  I1 =>  \MP1\,
                  I2 =>  \MP3A\,
                  I3 => \&40428\ );

  \=36406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36406\,
                  I0 =>  \36405\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36407\,
                  I0 =>  \T02/\,
                  I1 =>  \36406\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \2XP5\     
  \=36408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36408\,
                  I0 =>  \T02/\,
                  I1 =>  \DV0/\,
                  I2 =>  \BR1\,
                  I3 =>  '0' );

  -- Alias \RA/\      
  \=36409\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36409\,
                  I0 =>  \36404\,
                  I1 =>  \36432\,
                  I2 =>  \36446\,
                  I3 => \&39123\ );

  -- Alias \RSC/\     
  \=36410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36410\,
                  I0 =>  \36407\,
                  I1 =>  \36435\,
                  I2 =>  \36456\,
                  I3 => \&34158\ );

  -- Alias \WG/\      
  \=36411\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36411\,
                  I0 =>  \36407\,
                  I1 =>  \36360\,
                  I2 =>  \36435\,
                  I3 => \&39139\ );

  -- Alias \TMZ/\     
  \=36412\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36412\,
                  I0 =>  \36404\,
                  I1 =>  \36408\,
                  I2 =>  '0',
                  I3 => \&39135\ );

  \=36413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36413\,
                  I0 =>  \MP0/\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36414\,
                  I0 =>  \INOUT/\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY/\      
  \=36415\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36415\,
                  I0 =>  \36414\,
                  I1 =>  \36443\,
                  I2 =>  \36457\,
                  I3 => \&36441\ );

  -- Alias \3XP2\     
  \=36416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36416\,
                  I0 =>  \T03/\,
                  I1 =>  \TS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR1B2\    
  \=36417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36417\,
                  I0 =>  \BR1\,
                  I1 =>  \BR2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR1B2/\   
  \=36418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36418\,
                  I0 =>  \36417\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR12B\    
  \=36419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36419\,
                  I0 =>  \BR1/\,
                  I1 =>  \BR2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR12B/\   
  \=36420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36420\,
                  I0 =>  \36419\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BRDIF/\   
  \=36421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36421\,
                  I0 =>  \36417\,
                  I1 =>  \36419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR1B2B\   
  \=36422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36422\,
                  I0 =>  \BR2\,
                  I1 =>  \BR1\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BR1B2B/\  
  \=36423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36423\,
                  I0 =>  \36422\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36424\,
                  I0 =>  \36421\,
                  I1 =>  \TS0/\,
                  I2 =>  \T04/\,
                  I3 =>  '0' );

  \=36425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36425\,
                  I0 =>  \T04/\,
                  I1 =>  \BR1\,
                  I2 =>  \MP0/\,
                  I3 =>  '0' );

  -- Alias \WL/\      
  \=36426\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36426\,
                  I0 =>  \36425\,
                  I1 =>  \36427\,
                  I2 =>  \36447\,
                  I3 => \&39437\ );

  \=36427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36427\,
                  I0 =>  \MP0/\,
                  I1 =>  \BR1/\,
                  I2 =>  \T04/\,
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=36428\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36428\,
                  I0 =>  \36427\,
                  I1 =>  \36408\,
                  I2 =>  \36439\,
                  I3 => \&39144\ );

  -- Alias \4XP5\     
  \=36429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36429\,
                  I0 =>  \TS0/\,
                  I1 =>  \T04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=36430\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36430\,
                  I0 =>  \36425\,
                  I1 =>  \36457\,
                  I2 =>  \36437\,
                  I3 => \&39110\ );

  \=36431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36431\,
                  I0 =>  \DV1/\,
                  I1 =>  \T04/\,
                  I2 =>  \BR2/\,
                  I3 =>  '0' );

  -- Alias \8XP5\     
  \=36432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36432\,
                  I0 =>  \T08/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \4XP11\    
  \=36433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36433\,
                  I0 =>  \T04/\,
                  I1 =>  \INOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8XP6\     
  \=36434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36434\,
                  I0 =>  \T08/\,
                  I1 =>  \DV1/\,
                  I2 =>  \BR2\,
                  I3 =>  '0' );

  \=36435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36435\,
                  I0 =>  \T04/\,
                  I1 =>  \MP3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36436\,
                  I0 =>  \TS0/\,
                  I1 =>  \T05/\,
                  I2 =>  \BR1B2/\,
                  I3 =>  '0' );

  \=36437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36437\,
                  I0 =>  \T09/\,
                  I1 =>  \BR1\,
                  I2 =>  \MP0/\,
                  I3 =>  '0' );

  \=36438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36438\,
                  I0 =>  \T05/\,
                  I1 =>  \TS0/\,
                  I2 =>  \BR12B/\,
                  I3 =>  '0' );

  \=36439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36439\,
                  I0 =>  \T09/\,
                  I1 =>  \MP0/\,
                  I2 =>  \BR1/\,
                  I3 =>  '0' );

  -- Alias \CI/\      
  \=36440\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36440\,
                  I0 =>  \36424\,
                  I1 =>  \36444\,
                  I2 =>  '0',
                  I3 => \&39154\ );

  -- Alias \WY/\      
  \=36441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36441\,
                  I0 =>  \36439\,
                  I1 =>  \36432\,
                  I2 =>  \36437\,
                  I3 => \&39153\ );

  -- Alias \TSGN/\    
  \=36442\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36442\,
                  I0 =>  \36404\,
                  I1 =>  \36450\,
                  I2 =>  '0',
                  I3 => \&36454\ );

  -- Alias \B15X\     
  \=36443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36443\,
                  I0 =>  \T05/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36444\,
                  I0 =>  \MP0/\,
                  I1 =>  \T09/\,
                  I2 =>  \36421\,
                  I3 =>  '0' );

  -- Alias \5XP4\     
  \=36445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36445\,
                  I0 =>  \T05/\,
                  I1 =>  \RSM3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36446\,
                  I0 =>  \T09/\,
                  I1 =>  \MP3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \6XP5\     
  \=36447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36447\,
                  I0 =>  \T06/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \KRPT\     
  \=36448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36448\,
                  I0 =>  \T09/\,
                  I1 =>  \RUPT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TL15\     
  \=36449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36449\,
                  I0 =>  \T06/\,
                  I1 =>  \MP3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MP0T10\   
  \=36450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36450\,
                  I0 =>  \T10/\,
                  I1 =>  \MP0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36451\,
                  I0 =>  \BR1/\,
                  I1 =>  \MP0/\,
                  I2 =>  \T11/\,
                  I3 =>  '0' );

  -- Alias \RB1/\     
  \=36452\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36452\,
                  I0 =>  \36436\,
                  I1 =>  \36451\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \R1C/\     
  \=36453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36453\,
                  I0 =>  \36451\,
                  I1 =>  \36438\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TSGN/\    
  \=36454\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36454\,
                  I0 =>  \36431\,
                  I1 =>  \36413\,
                  I2 =>  \36456\,
                  I3 => \&39443\ );

  -- Alias \TSGN2\    
  \=36455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36455\,
                  I0 =>  \T07/\,
                  I1 =>  \MP0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=36456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36456\,
                  I0 =>  \T07/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \7XP19\    
  \=36457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \36457\,
                  I0 =>  \T07/\,
                  I1 =>  \BR1/\,
                  I2 =>  \MP3/\,
                  I3 =>  '0' );

  -- Alias \MRSC\     
  \=36459\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36459\,
                  I0 =>  \36410\,
                  I1 =>  \36410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L16/\     
  \=36460\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&36460\,
                  I0 =>  \36451\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ********************************************
  -- ***                                      ***
  -- ***  A5 /1 - CROSS POINT GENERATOR NQI.  ***
  -- ***                                      ***
  -- ********************************************

  \=39101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39101\,
                  I0 =>  \IC10\,
                  I1 =>  \IC3\,
                  I2 =>  \IC2\,
                  I3 =>  '0' );

  \=39102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39102\,
                  I0 =>  \T01/\,
                  I1 =>  \39101\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39103\,
                  I0 =>  \T01/\,
                  I1 =>  \IC10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MONEX/\   
  \=39104\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39104\,
                  I0 =>  \10XP6\,
                  I1 =>  \10XP7\,
                  I2 =>  \39103\,
                  I3 =>  '0' );

  \=39105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39105\,
                  I0 =>  \STD2\,
                  I1 =>  \IC2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39106\,
                  I0 =>  \T01/\,
                  I1 =>  \39105\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RZ/\      
  \=39107\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39107\,
                  I0 =>  \39106\,
                  I1 =>  \39122\,
                  I2 =>  \39131\,
                  I3 => \&39155\ );

  \=39108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39108\,
                  I0 =>  \TC0\,
                  I1 =>  \TCF0\,
                  I2 =>  \IC4\,
                  I3 =>  '0' );

  \=39109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39109\,
                  I0 =>  \T01/\,
                  I1 =>  \39108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=39110\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39110\,
                  I0 =>  \39109\,
                  I1 =>  \39120\,
                  I2 =>  '0',
                  I3 => \&39146\ );

  \=39111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39111\,
                  I0 =>  \IC2\,
                  I1 =>  \IC3\,
                  I2 =>  \RSM3\,
                  I3 =>  '0' );

  \=39112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39112\,
                  I0 =>  \T02/\,
                  I1 =>  \39111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NISQ/\    
  \=39113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39113\,
                  I0 =>  \39112\,
                  I1 =>  \39117\,
                  I2 =>  \8XP15\,
                  I3 =>  '0' );

  -- Alias \DVST\     
  \=39115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39115\,
                  I0 =>  \T02/\,
                  I1 =>  \STD2\,
                  I2 =>  \DIV/\,
                  I3 =>  '0' );

  \=39116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39116\,
                  I0 =>  \MP3/\,
                  I1 =>  \T10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \2XP7\     
  \=39117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39117\,
                  I0 =>  \T02/\,
                  I1 =>  \MP3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39120\,
                  I0 =>  \T03/\,
                  I1 =>  \IC2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39121\,
                  I0 =>  \T01/\,
                  I1 =>  \IC15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3XP6\     
  \=39122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39122\,
                  I0 =>  \T03/\,
                  I1 =>  \TC0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RA/\      
  \=39123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39123\,
                  I0 =>  \39121\,
                  I1 =>  \39124\,
                  I2 =>  '0',
                  I3 => \&39226\ );

  \=39124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39124\,
                  I0 =>  \T04/\,
                  I1 =>  \IC2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39125\,
                  I0 =>  \T02/\,
                  I1 =>  \IC15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TPZG/\    
  \=39126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39126\,
                  I0 =>  \39125\,
                  I1 =>  \39134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39127\,
                  I0 =>  \T04/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WA/\      
  \=39128\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39128\,
                  I0 =>  \39127\,
                  I1 =>  \39129\,
                  I2 =>  '0',
                  I3 => \&39244\ );

  \=39129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39129\,
                  I0 =>  \T04/\,
                  I1 =>  \MASK0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL/\      
  \=39130\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39130\,
                  I0 =>  \39127\,
                  I1 =>  \39116\,
                  I2 =>  \8XP12\,
                  I3 =>  '0' );

  \=39131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39131\,
                  I0 =>  \T05/\,
                  I1 =>  \IC2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PARTC\    
  \=39132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39132\,
                  I0 =>  \INKL/\,
                  I1 =>  \SHIFT\,
                  I2 =>  \MON+CH\,
                  I3 =>  '0' );

  \=39133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39133\,
                  I0 =>  \39132\,
                  I1 =>  \PRINC\,
                  I2 =>  \CCS0\,
                  I3 =>  '0' );

  \=39134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39134\,
                  I0 =>  \T05/\,
                  I1 =>  \39133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TMZ/\     
  \=39135\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39135\,
                  I0 =>  \39121\,
                  I1 =>  \39134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP12\    
  \=39136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39136\,
                  I0 =>  \T05/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TSGN/\    
  \=39137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39137\,
                  I0 =>  \39134\,
                  I1 =>  \39121\,
                  I2 =>  \39147\,
                  I3 => \&36442\ );

  \=39138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39138\,
                  I0 =>  \T06/\,
                  I1 =>  \RSM3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WG/\      
  \=39139\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39139\,
                  I0 =>  \9XP5\,
                  I1 =>  \39121\,
                  I2 =>  \39138\,
                  I3 => \&40342\ );

  \=39140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39140\,
                  I0 =>  \T06/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RG/\      
  \=39141\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39141\,
                  I0 =>  \39134\,
                  I1 =>  \39149\,
                  I2 =>  \39140\,
                  I3 => \&39325\ );

  \=39143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39143\,
                  I0 =>  \MSU0/\,
                  I1 =>  \T06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=39144\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39144\,
                  I0 =>  \39129\,
                  I1 =>  \39143\,
                  I2 =>  '0',
                  I3 => \&39242\ );

  \=39145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39145\,
                  I0 =>  \T07/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=39146\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39146\,
                  I0 =>  \39138\,
                  I1 =>  \39145\,
                  I2 =>  '0',
                  I3 => \&39204\ );

  -- Alias \7XP9\     
  \=39147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39147\,
                  I0 =>  \T07/\,
                  I1 =>  \MSU0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A2X/\     
  \=39148\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39148\,
                  I0 =>  \39149\,
                  I1 =>  \39143\,
                  I2 =>  \39140\,
                  I3 => \&39334\ );

  \=39149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39149\,
                  I0 =>  \T07/\,
                  I1 =>  \IC2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \7XP4\     
  \=39150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39150\,
                  I0 =>  \CCS0/\,
                  I1 =>  \T07/\,
                  I2 =>  \BR2/\,
                  I3 =>  '0' );

  -- Alias \PTWOX\    
  \=39151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39151\,
                  I0 =>  \BR1/\,
                  I1 =>  \CCS0/\,
                  I2 =>  \T07/\,
                  I3 =>  '0' );

  \=39152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39152\,
                  I0 =>  \T07/\,
                  I1 =>  \CCS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY/\      
  \=39153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39153\,
                  I0 =>  \39149\,
                  I1 =>  \39143\,
                  I2 =>  \39140\,
                  I3 => \&39234\ );

  -- Alias \CI/\      
  \=39154\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39154\,
                  I0 =>  \39143\,
                  I1 =>  \39102\,
                  I2 =>  \10XP6\,
                  I3 => \&39328\ );

  -- Alias \RZ/\      
  \=39155\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39155\,
                  I0 =>  \8XP3\,
                  I1 =>  \39152\,
                  I2 =>  \4XP5\,
                  I3 => \&39338\ );

  -- Alias \WY12/\    
  \=39156\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39156\,
                  I0 =>  \4XP5\,
                  I1 =>  \39152\,
                  I2 =>  \39102\,
                  I3 =>  '0' );

  \=39201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39201\,
                  I0 =>  \T08/\,
                  I1 =>  \CCS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WZ/\      
  \=39202\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39202\,
                  I0 =>  \39120\,
                  I1 =>  \39221\,
                  I2 =>  \39201\,
                  I3 => \&39417\ );

  \=39203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39203\,
                  I0 =>  \INKL/\,
                  I1 =>  \FETCH0\,
                  I2 =>  \T08/\,
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=39204\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39204\,
                  I0 =>  \39203\,
                  I1 =>  \39223\,
                  I2 =>  '0',
                  I3 => \&39336\ );

  -- Alias \TSUDO/\   
  \=39205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39205\,
                  I0 =>  \IC3\,
                  I1 =>  \RSM3\,
                  I2 =>  \MP3\,
                  I3 => \&39206\ );

  -- Alias \39205\    
  \=39206\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39206\,
                  I0 =>  \IC16\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RAD\      
  \=39207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39207\,
                  I0 =>  \39205\,
                  I1 =>  \T08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WB/\      
  \=39208\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39208\,
                  I0 =>  \39207\,
                  I1 =>  \39217\,
                  I2 =>  '0',
                  I3 => \&39315\ );

  \=39209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39209\,
                  I0 =>  \IC16\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8XP15\    
  \=39210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39210\,
                  I0 =>  \T08/\,
                  I1 =>  \39209\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39211\,
                  I0 =>  \MP0\,
                  I1 =>  \IC1\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8XP3\     
  \=39212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39212\,
                  I0 =>  \T08/\,
                  I1 =>  \39211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39213\,
                  I0 =>  \IC2\,
                  I1 =>  \IC4\,
                  I2 =>  \DXCH0\,
                  I3 =>  '0' );

  \=39214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39214\,
                  I0 =>  \T08/\,
                  I1 =>  \39213\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RU/\      
  \=39215\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39215\,
                  I0 =>  \39201\,
                  I1 =>  \39214\,
                  I2 =>  \39224\,
                  I3 => \&39429\ );

  \=39216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39216\,
                  I0 =>  \DXCH0\,
                  I1 =>  \GOJ1\,
                  I2 =>  \DAS0\,
                  I3 =>  '0' );

  \=39217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39217\,
                  I0 =>  \T08/\,
                  I1 =>  \39216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSTRT\    
  \=39219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39219\,
                  I0 =>  \T08/\,
                  I1 =>  \GOJ1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8XP12\    
  \=39220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39220\,
                  I0 =>  \T08/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39221\,
                  I0 =>  \T08/\,
                  I1 =>  \TCSAJ3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39222\,
                  I0 =>  \IC2\,
                  I1 =>  \DV1B1B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39223\,
                  I0 =>  \T09/\,
                  I1 =>  \39222\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \9XP5\     
  \=39224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39224\,
                  I0 =>  \T09/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39225\,
                  I0 =>  \T09/\,
                  I1 =>  \MASK0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RA/\      
  \=39226\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39226\,
                  I0 =>  \39225\,
                  I1 =>  \39233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39227\,
                  I0 =>  \T10/\,
                  I1 =>  \CCS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST2/\     
  \=39228\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39228\,
                  I0 =>  \39221\,
                  I1 =>  \39227\,
                  I2 =>  '0',
                  I3 => \&40416\ );

  -- Alias \10XP6\    
  \=39229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39229\,
                  I0 =>  \CCS0/\,
                  I1 =>  \BR2\,
                  I2 =>  \T10/\,
                  I3 =>  '0' );

  \=39230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39230\,
                  I0 =>  \IC1\,
                  I1 =>  \IC10\,
                  I2 =>  \RUPT0\,
                  I3 =>  '0' );

  -- Alias \10XP1\    
  \=39231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39231\,
                  I0 =>  \39230\,
                  I1 =>  \T10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39232\,
                  I0 =>  \DAS0\,
                  I1 =>  \39239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39233\,
                  I0 =>  \T10/\,
                  I1 =>  \39232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY/\      
  \=39234\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39234\,
                  I0 =>  \39227\,
                  I1 =>  \39225\,
                  I2 =>  \39233\,
                  I3 => \&40119\ );

  \=39235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39235\,
                  I0 =>  \39239\,
                  I1 =>  \39237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \10XP7\    
  \=39236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39236\,
                  I0 =>  \T10/\,
                  I1 =>  \39235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39237\,
                  I0 =>  \BR12B/\,
                  I1 =>  \DAS0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \10XP8\    
  \=39238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39238\,
                  I0 =>  \T10/\,
                  I1 =>  \DAS0/\,
                  I2 =>  \BR1B2/\,
                  I3 =>  '0' );

  \=39239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39239\,
                  I0 =>  \MSU0/\,
                  I1 =>  \BR1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \11XP2\    
  \=39240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39240\,
                  I0 =>  \T11/\,
                  I1 =>  \MSU0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39241\,
                  I0 =>  \T11/\,
                  I1 =>  \MASK0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=39242\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39242\,
                  I0 =>  \39225\,
                  I1 =>  \39241\,
                  I2 =>  '0',
                  I3 => \&39418\ );

  \=39243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39243\,
                  I0 =>  \T11/\,
                  I1 =>  \39245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WA/\      
  \=39244\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39244\,
                  I0 =>  \39223\,
                  I1 =>  \39243\,
                  I2 =>  \5XP11\,
                  I3 => \&39422\ );

  \=39245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39245\,
                  I0 =>  \MSU0\,
                  I1 =>  \IC14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39248\,
                  I0 =>  \GOJAM\,
                  I1 =>  \39249\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GNHNC\    
  \:39249\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \39249\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$39249\,
                   R => '0',
                   S => SYSRESET );

  \=39249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$39249\,
                  I0 =>  \39248\,
                  I1 =>  \T01\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39250\,
                  I0 =>  \C24A\,
                  I1 =>  \C25A\,
                  I2 =>  \C26A\,
                  I3 => \&39251\ );

  -- Alias \39250\    
  \=39251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39251\,
                  I0 =>  \C27A\,
                  I1 =>  \C30A\,
                  I2 =>  '0',
                  I3 => \&39252\ );

  -- Alias \39250\    
  \=39252\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39252\,
                  I0 =>  \C37P\,
                  I1 =>  \C40P\,
                  I2 =>  \C41P\,
                  I3 => \&39253\ );

  -- Alias \39250\    
  \=39253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39253\,
                  I0 =>  \C42P\,
                  I1 =>  \C43P\,
                  I2 =>  \C44P\,
                  I3 =>  '0' );

  \=39254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39254\,
                  I0 =>  \INCSET/\,
                  I1 =>  \39250\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PINC/\    
  \:39255\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \39255\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$39255\,
                   R => '0',
                   S => SYSRESET );

  \=39255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$39255\,
                  I0 =>  \39254\,
                  I1 =>  \39256\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PINC\     
  \=39256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39256\,
                  I0 =>  \39255\,
                  I1 =>  \T12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P03\      
  \=39261\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39261\,
                  I0 =>  '0',
                  I1 =>  \EDSET\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ********************************************
  -- ***                                      ***
  -- ***  A5 /2 - CROSS POINT GENERATOR NQI.  ***
  -- ***                                      ***
  -- ********************************************

  \=39301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39301\,
                  I0 =>  \IC12\,
                  I1 =>  \DAS0\,
                  I2 =>  \DAS1\,
                  I3 => \&39302\ );

  -- Alias \39301\    
  \=39302\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39302\,
                  I0 =>  \IC9\,
                  I1 =>  \DXCH0\,
                  I2 =>  '0',
                  I3 => \&39303\ );

  -- Alias \39301\    
  \=39303\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39303\,
                  I0 =>  \PRINC\,
                  I1 =>  \INOUT\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL10BB\   
  \=39304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39304\,
                  I0 =>  \T01/\,
                  I1 =>  \39301\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WS/\      
  \=39305\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39305\,
                  I0 =>  \39304\,
                  I1 =>  \39307\,
                  I2 =>  \39309\,
                  I3 =>  '0' );

  -- Alias \R6\       
  \=39306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39306\,
                  I0 =>  \T01/\,
                  I1 =>  \FETCH0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39307\,
                  I0 =>  \T01/\,
                  I1 =>  \CHINC/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \2XP8\     
  \=39308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39308\,
                  I0 =>  \FETCH0/\,
                  I1 =>  \T02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSCT\     
  \=39309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39309\,
                  I0 =>  \MON+CH\,
                  I1 =>  \T01/\,
                  I2 =>  \INKL/\,
                  I3 =>  '0' );

  \=39310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39310\,
                  I0 =>  \TS0\,
                  I1 =>  \DAS0\,
                  I2 =>  \MASK0\,
                  I3 => \&39311\ );

  -- Alias \39310\    
  \=39311\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39311\,
                  I0 =>  \IC5\,
                  I1 =>  \MP0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39312\,
                  I0 =>  \T03/\,
                  I1 =>  \39310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39313\,
                  I0 =>  \T03/\,
                  I1 =>  \IC8/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RQ\       
  \=39314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39314\,
                  I0 =>  \T03/\,
                  I1 =>  \QXCH0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WB/\      
  \=39315\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39315\,
                  I0 =>  \39312\,
                  I1 =>  \39314\,
                  I2 =>  \39313\,
                  I3 => \&39316\ );

  -- Alias \WB/\      
  \=39316\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39316\,
                  I0 =>  \39320\,
                  I1 =>  \39324\,
                  I2 =>  \6XP2\,
                  I3 => \&39434\ );

  \=39318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39318\,
                  I0 =>  \DV1\,
                  I1 =>  \INOUT\,
                  I2 =>  \IC2\,
                  I3 =>  '0' );

  \=39319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39319\,
                  I0 =>  \T04/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39320\,
                  I0 =>  \T04/\,
                  I1 =>  \39318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL/\      
  \=39321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39321\,
                  I0 =>  \39313\,
                  I1 =>  \39319\,
                  I2 =>  \11XP6\,
                  I3 => \&39130\ );

  -- Alias \RA/\      
  \=39322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39322\,
                  I0 =>  \39312\,
                  I1 =>  \6XP2\,
                  I2 =>  '0',
                  I3 => \&36355\ );

  -- Alias \TRSM\     
  \=39323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39323\,
                  I0 =>  \T05/\,
                  I1 =>  \NDX0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39324\,
                  I0 =>  \IC12/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RG/\      
  \=39325\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39325\,
                  I0 =>  \39324\,
                  I1 =>  \39327\,
                  I2 =>  \39332\,
                  I3 => \&39326\ );

  -- Alias \RG/\      
  \=39326\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39326\,
                  I0 =>  \39337\,
                  I1 =>  \39339\,
                  I2 =>  \39344\,
                  I3 => \&39435\ );

  \=39327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39327\,
                  I0 =>  \DAS1/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI/\      
  \=39328\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39328\,
                  I0 =>  \39335\,
                  I1 =>  \39341\,
                  I2 =>  \39343\,
                  I3 =>  '0' );

  \=39329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39329\,
                  I0 =>  \PRINC\,
                  I1 =>  \DAS1\,
                  I2 =>  \PARTC\,
                  I3 =>  '0' );

  \=39330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39330\,
                  I0 =>  \39329\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY12/\    
  \=39331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39331\,
                  I0 =>  \39341\,
                  I1 =>  \39343\,
                  I2 =>  '0',
                  I3 => \&39156\ );

  -- Alias \5XP9\     
  \=39332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39332\,
                  I0 =>  \SHIFT/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY/\      
  \=39333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39333\,
                  I0 =>  \39330\,
                  I1 =>  \39308\,
                  I2 =>  \10XP10\,
                  I3 => \&36415\ );

  -- Alias \A2X/\     
  \=39334\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39334\,
                  I0 =>  \39327\,
                  I1 =>  \10XP10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39335\,
                  I0 =>  \SHANC/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=39336\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39336\,
                  I0 =>  \5XP19\,
                  I1 =>  \39341\,
                  I2 =>  '0',
                  I3 => \&40347\ );

  -- Alias \5XP13\    
  \=39337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39337\,
                  I0 =>  \IC8/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RZ/\      
  \=39338\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39338\,
                  I0 =>  \39343\,
                  I1 =>  \6XP7\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP15\    
  \=39339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39339\,
                  I0 =>  \QXCH0/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP21\    
  \=39340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39340\,
                  I0 =>  \CHINC/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39341\,
                  I0 =>  \IC16/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39342\,
                  I0 =>  \MP3\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39343\,
                  I0 =>  \39342\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39344\,
                  I0 =>  \IC5/\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \39346\    
  \=39345\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39345\,
                  I0 =>  \S11\,
                  I1 =>  \S12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SCAD\     
  \=39346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39346\,
                  I0 =>  \YT0/\,
                  I1 =>  \YB0/\,
                  I2 =>  \XT0/\,
                  I3 => \&39345\ );

  -- Alias \SCAD/\    
  \=39347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39347\,
                  I0 =>  \39346\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39348\,
                  I0 =>  \YB0/\,
                  I1 =>  \YT0/\,
                  I2 =>  '0',
                  I3 => \&39349\ );

  -- Alias \39348\    
  \=39349\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39349\,
                  I0 =>  \S12\,
                  I1 =>  \S11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NDR100/\  
  \=39350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39350\,
                  I0 =>  \39348\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OCTAD2\   
  \=39352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39352\,
                  I0 =>  \XT2/\,
                  I1 =>  \39350\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OCTAD3\   
  \=39353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39353\,
                  I0 =>  \39350\,
                  I1 =>  \XT3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OCTAD4\   
  \=39354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39354\,
                  I0 =>  \39350\,
                  I1 =>  \XT4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OCTAD5\   
  \=39355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39355\,
                  I0 =>  \39350\,
                  I1 =>  \XT5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OCTAD6\   
  \=39356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39356\,
                  I0 =>  \39350\,
                  I1 =>  \XT6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39401\,
                  I0 =>  \BR1/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DV1B1B\   
  \=39402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39402\,
                  I0 =>  \DV1/\,
                  I1 =>  \BR1\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39403\,
                  I0 =>  \39401\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39404\,
                  I0 =>  \RAND0\,
                  I1 =>  \WAND0\,
                  I2 =>  \39401\,
                  I3 =>  '0' );

  \=39405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39405\,
                  I0 =>  \ROR0\,
                  I1 =>  \39402\,
                  I2 =>  \WOR0\,
                  I3 =>  '0' );

  \=39406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39406\,
                  I0 =>  \39404\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \5XP19\    
  \=39407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39407\,
                  I0 =>  \T05/\,
                  I1 =>  \39405\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39408\,
                  I0 =>  \TS0/\,
                  I1 =>  \BRDIF/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39409\,
                  I0 =>  \IC2\,
                  I1 =>  \IC5\,
                  I2 =>  \READ0\,
                  I3 => \&39410\ );

  -- Alias \39409\    
  \=39410\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39410\,
                  I0 =>  \39408\,
                  I1 =>  \DV4\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39411\,
                  I0 =>  \39403\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39412\,
                  I0 =>  \39409\,
                  I1 =>  \T05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z16/\     
  \=39413\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39413\,
                  I0 =>  \39411\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \39415\    
  \=39414\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39414\,
                  I0 =>  \IC2\,
                  I1 =>  \IC3\,
                  I2 =>  \TS0\,
                  I3 =>  '0' );

  \=39415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39415\,
                  I0 =>  \IC16\,
                  I1 =>  \MP3\,
                  I2 =>  '0',
                  I3 => \&39414\ );

  \=39416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39416\,
                  I0 =>  \T06/\,
                  I1 =>  \39415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WZ/\      
  \=39417\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39417\,
                  I0 =>  \39416\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=39418\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39418\,
                  I0 =>  \39406\,
                  I1 =>  \39432\,
                  I2 =>  '0',
                  I3 => \&39423\ );

  -- Alias \6XP8\     
  \=39419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39419\,
                  I0 =>  \T06/\,
                  I1 =>  \DAS1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \6XP7\     
  \=39420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39420\,
                  I0 =>  \DV4/\,
                  I1 =>  \T06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \6XP2\     
  \=39421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39421\,
                  I0 =>  \T06/\,
                  I1 =>  \RXOR0\,
                  I2 =>  \INOUT/\,
                  I3 =>  '0' );

  -- Alias \WA/\      
  \=39422\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39422\,
                  I0 =>  \39412\,
                  I1 =>  \39432\,
                  I2 =>  '0',
                  I3 => \&40328\ );

  -- Alias \RC/\      
  \=39423\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39423\,
                  I0 =>  \39439\,
                  I1 =>  \39451\,
                  I2 =>  '0',
                  I3 => \&40415\ );

  -- Alias \TOV/\     
  \=39424\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39424\,
                  I0 =>  \39420\,
                  I1 =>  \39419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39425\,
                  I0 =>  \STFET1/\,
                  I1 =>  \T07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \U2BBK\    
  \=39426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39426\,
                  I0 =>  \STFET1/\,
                  I1 =>  \MONWBK\,
                  I2 =>  \T08/\,
                  I3 =>  '0' );

  \=39427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39427\,
                  I0 =>  \IC13\,
                  I1 =>  \IC14\,
                  I2 =>  \DV1\,
                  I3 =>  '0' );

  \=39428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39428\,
                  I0 =>  \T07/\,
                  I1 =>  \39427\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RU/\      
  \=39429\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39429\,
                  I0 =>  \39416\,
                  I1 =>  \39419\,
                  I2 =>  \5XP11\,
                  I3 => \&39430\ );

  -- Alias \RU/\      
  \=39430\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39430\,
                  I0 =>  \39441\,
                  I1 =>  \39436\,
                  I2 =>  \39452\,
                  I3 => \&40157\ );

  -- Alias \RSTSTG\   
  \=39431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39431\,
                  I0 =>  \T08/\,
                  I1 =>  \DV4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39432\,
                  I0 =>  \T09/\,
                  I1 =>  \39403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z15/\     
  \=39433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39433\,
                  I0 =>  \39432\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WB/\      
  \=39434\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39434\,
                  I0 =>  \39428\,
                  I1 =>  \39436\,
                  I2 =>  \39441\,
                  I3 => \&40153\ );

  -- Alias \RG/\      
  \=39435\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39435\,
                  I0 =>  \39428\,
                  I1 =>  \39425\,
                  I2 =>  \39451\,
                  I3 => \&40141\ );

  \=39436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39436\,
                  I0 =>  \T09/\,
                  I1 =>  \DV4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL/\      
  \=39437\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39437\,
                  I0 =>  \5XP13\,
                  I1 =>  \39452\,
                  I2 =>  '0',
                  I3 => \&39438\ );

  -- Alias \WL/\      
  \=39438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39438\,
                  I0 =>  \39436\,
                  I1 =>  \39449\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39439\,
                  I0 =>  \T09/\,
                  I1 =>  \DAS1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TMZ/\     
  \=39440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39440\,
                  I0 =>  \39439\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36412\ );

  \=39441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39441\,
                  I0 =>  \T10/\,
                  I1 =>  \39445\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \10XP10\   
  \=39442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39442\,
                  I0 =>  \T10/\,
                  I1 =>  \IC11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TSGN/\    
  \=39443\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39443\,
                  I0 =>  \39431\,
                  I1 =>  \5XP9\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WYD/\     
  \=39444\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&39444\,
                  I0 =>  \5XP9\,
                  I1 =>  \39450\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39445\,
                  I0 =>  \IC14\,
                  I1 =>  \IC2\,
                  I2 =>  \DV1\,
                  I3 =>  '0' );

  -- Alias \DV4B1B\   
  \=39446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39446\,
                  I0 =>  \DV4/\,
                  I1 =>  \BR1\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39447\,
                  I0 =>  \DAS1/\,
                  I1 =>  \ADS0\,
                  I2 =>  \BR2\,
                  I3 =>  '0' );

  \=39448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39448\,
                  I0 =>  \39446\,
                  I1 =>  \IC4\,
                  I2 =>  \39447\,
                  I3 =>  '0' );

  \=39449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39449\,
                  I0 =>  \T10/\,
                  I1 =>  \39448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \11XP6\    
  \=39450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39450\,
                  I0 =>  \T11/\,
                  I1 =>  \DV1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39451\,
                  I0 =>  \T11/\,
                  I1 =>  \RXOR0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=39452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \39452\,
                  I0 =>  \T12/\,
                  I1 =>  \T12USE/\,
                  I2 =>  \DV1/\,
                  I3 =>  '0' );

  -- *******************************************
  -- ***                                     ***
  -- ***  A6 /1 - CROSS POINT GENERATOR II.  ***
  -- ***                                     ***
  -- *******************************************

  \=40101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40101\,
                  I0 =>  \T04\,
                  I1 =>  \T07\,
                  I2 =>  \T10\,
                  I3 =>  '0' );

  \=40102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40102\,
                  I0 =>  \40101\,
                  I1 =>  \DV376/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40103\,
                  I0 =>  \T01/\,
                  I1 =>  \DV1376/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40104\,
                  I0 =>  \T04/\,
                  I1 =>  \DV4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40105\,
                  I0 =>  \40102\,
                  I1 =>  \40103\,
                  I2 =>  \40104\,
                  I3 =>  '0' );

  -- Alias \DVXP1\    
  \=40106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40106\,
                  I0 =>  \40105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A2X/\     
  \=40107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40107\,
                  I0 =>  \7XP19\,
                  I1 =>  \40117\,
                  I2 =>  \40106\,
                  I3 => \&39148\ );

  -- Alias \L2GD/\    
  \=40108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40108\,
                  I0 =>  \40106\,
                  I1 =>  \40117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=40109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40109\,
                  I0 =>  \40106\,
                  I1 =>  \40128\,
                  I2 =>  \RBSQ\,
                  I3 => \&36335\ );

  -- Alias \WYD/\     
  \=40110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40110\,
                  I0 =>  \40106\,
                  I1 =>  \40118\,
                  I2 =>  '0',
                  I3 => \&39444\ );

  \=40111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40111\,
                  I0 =>  \T01\,
                  I1 =>  \T03\,
                  I2 =>  \T05\,
                  I3 => \&40112\ );

  -- Alias \40111\    
  \=40112\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40112\,
                  I0 =>  \T07\,
                  I1 =>  \T09\,
                  I2 =>  \T11\,
                  I3 =>  '0' );

  \=40113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40113\,
                  I0 =>  \MP1/\,
                  I1 =>  \40111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40114\,
                  I0 =>  \40113\,
                  I1 =>  \2XP7\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40115\,
                  I0 =>  \40114\,
                  I1 =>  \40125\,
                  I2 =>  \40126\,
                  I3 =>  '0' );

  \=40116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40116\,
                  I0 =>  \40126\,
                  I1 =>  \40125\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZIP\      
  \=40117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40117\,
                  I0 =>  \40114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40118\,
                  I0 =>  \40114\,
                  I1 =>  \40116\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WY/\      
  \=40119\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40119\,
                  I0 =>  \40115\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40120\,
                  I0 =>  \L01/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40121\,
                  I0 =>  \L02A/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40122\,
                  I0 =>  \L15A/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40123\,
                  I0 =>  \40126\,
                  I1 =>  \40125\,
                  I2 =>  \L02A/\,
                  I3 =>  '0' );

  \=40124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40124\,
                  I0 =>  \40120\,
                  I1 =>  \40121\,
                  I2 =>  \40122\,
                  I3 =>  '0' );

  \=40125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40125\,
                  I0 =>  \40122\,
                  I1 =>  \40120\,
                  I2 =>  \L02A/\,
                  I3 =>  '0' );

  \=40126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40126\,
                  I0 =>  \40121\,
                  I1 =>  \L15A/\,
                  I2 =>  \L01/\,
                  I3 =>  '0' );

  \=40127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40127\,
                  I0 =>  \40123\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40128\,
                  I0 =>  \40123\,
                  I1 =>  \40124\,
                  I2 =>  \40114\,
                  I3 =>  '0' );

  \=40129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40129\,
                  I0 =>  \40114\,
                  I1 =>  \40127\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZIPCI\    
  \=40130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40130\,
                  I0 =>  \40114\,
                  I1 =>  \40127\,
                  I2 =>  \40133\,
                  I3 =>  '0' );

  -- Alias \RC/\      
  \=40131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40131\,
                  I0 =>  \40130\,
                  I1 =>  \3XP7\,
                  I2 =>  '0',
                  I3 => \&36339\ );

  -- Alias \RCH/\     
  \=40132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40132\,
                  I0 =>  \3XP7\,
                  I1 =>  \5XP21\,
                  I2 =>  \4XP11\,
                  I3 =>  '0' );

  \=40133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40133\,
                  I0 =>  \L15A/\,
                  I1 =>  \L02A/\,
                  I2 =>  \L01/\,
                  I3 =>  '0' );

  \=40134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40134\,
                  I0 =>  \T05\,
                  I1 =>  \T08\,
                  I2 =>  \T11\,
                  I3 =>  '0' );

  \=40135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40135\,
                  I0 =>  \40134\,
                  I1 =>  \DV376/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40136\,
                  I0 =>  \DV1376/\,
                  I1 =>  \T02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40137\,
                  I0 =>  \40135\,
                  I1 =>  \40136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40138\,
                  I0 =>  \40137\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TSGU/\    
  \=40139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40139\,
                  I0 =>  \5XP28\,
                  I1 =>  \40138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL/\      
  \=40140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40140\,
                  I0 =>  \40138\,
                  I1 =>  \5XP12\,
                  I2 =>  '0',
                  I3 => \&36426\ );

  -- Alias \40146\    
  \=40141\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40141\,
                  I0 =>  \5XP4\,
                  I1 =>  \RADRG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40142\,
                  I0 =>  \T06\,
                  I1 =>  \T09\,
                  I2 =>  \T12\,
                  I3 =>  '0' );

  \=40143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40143\,
                  I0 =>  \DV376/\,
                  I1 =>  \40142\,
                  I2 =>  \T12USE/\,
                  I3 =>  '0' );

  \=40144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40144\,
                  I0 =>  \40143\,
                  I1 =>  \DIVSTG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40145\,
                  I0 =>  \40144\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RG/\      
  \=40146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40146\,
                  I0 =>  \40138\,
                  I1 =>  \5XP28\,
                  I2 =>  '0',
                  I3 => \&39141\ );

  \=40147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40147\,
                  I0 =>  \T02\,
                  I1 =>  \T04\,
                  I2 =>  \T06\,
                  I3 => \&40148\ );

  -- Alias \40147\    
  \=40148\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40148\,
                  I0 =>  \T08\,
                  I1 =>  \T10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40149\,
                  I0 =>  \T01\,
                  I1 =>  \T03\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40150\,
                  I0 =>  \MP1/\,
                  I1 =>  \40147\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40151\,
                  I0 =>  \40149\,
                  I1 =>  \MP3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZAP/\     
  \=40152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40152\,
                  I0 =>  \40150\,
                  I1 =>  \40151\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40155\    
  \=40153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40153\,
                  I0 =>  \2XP3\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZAP\      
  \=40154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40154\,
                  I0 =>  \40152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WB/\      
  \=40155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40155\,
                  I0 =>  \5XP28\,
                  I1 =>  \1XP10\,
                  I2 =>  \40145\,
                  I3 => \&39208\ );

  -- Alias \RU/\      
  \=40156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40156\,
                  I0 =>  \40145\,
                  I1 =>  \40154\,
                  I2 =>  '0',
                  I3 => \&39215\ );

  -- Alias \40156\    
  \=40157\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40157\,
                  I0 =>  \5XP12\,
                  I1 =>  \6XP5\,
                  I2 =>  '0',
                  I3 => \&40344\ );

  -- Alias \WZ/\      
  \=40158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40158\,
                  I0 =>  \RRPA\,
                  I1 =>  \5XP4\,
                  I2 =>  '0',
                  I3 => \&39202\ );

  -- Alias \MCRO/\    
  \=40160\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40160\,
                  I0 =>  \40129\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB1F\     
  \=40201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40201\,
                  I0 =>  \BR1/\,
                  I1 =>  \PHS4/\,
                  I2 =>  \40139\,
                  I3 =>  '0' );

  -- Alias \CLXC\     
  \=40202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40202\,
                  I0 =>  \40139\,
                  I1 =>  \40139\,
                  I2 =>  \40139\,
                  I3 => \&40203\ );

  -- Alias \40202\    
  \=40203\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40203\,
                  I0 =>  \BR1\,
                  I1 =>  \BR1\,
                  I2 =>  \BR1\,
                  I3 => \&40204\ );

  -- Alias \40202\    
  \=40204\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40204\,
                  I0 =>  \PHS4/\,
                  I1 =>  \PHS4/\,
                  I2 =>  \PHS4/\,
                  I3 =>  '0' );

  -- Alias \WQ/\      
  \=40206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40206\,
                  I0 =>  \5XP15\,
                  I1 =>  \3XP6\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TOV/\     
  \=40207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40207\,
                  I0 =>  \6XP5\,
                  I1 =>  \3XP2\,
                  I2 =>  \9XP5\,
                  I3 => \&39424\ );

  -- Alias \WSC/\     
  \=40208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40208\,
                  I0 =>  \9XP5\,
                  I1 =>  \6XP8\,
                  I2 =>  '0',
                  I3 => \&40343\ );

  -- Alias \WG/\      
  \=40209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40209\,
                  I0 =>  \6XP8\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36345\ );

  -- Alias \MONEX\    
  \=40210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40210\,
                  I0 =>  \MONEX/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40213\,
                  I0 =>  \PTWOX\,
                  I1 =>  \40210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TWOX\     
  \=40214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40214\,
                  I0 =>  \40213\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40215\,
                  I0 =>  \40210\,
                  I1 =>  \B15X\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BXVX\     
  \=40216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40216\,
                  I0 =>  \40215\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40217\,
                  I0 =>  \40134\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIFL/\    
  \:40220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40220\,
                   R => '0',
                   S => SYSRESET );

  \=40220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40220\,
                  I0 =>  \40106\,
                  I1 =>  \40221\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40221\,
                  I0 =>  \40220\,
                  I1 =>  \40217\,
                  I2 =>  \T02\,
                  I3 =>  '0' );

  \=40222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40222\,
                  I0 =>  \RSTK/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSTKX/\   
  \=40224\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40224\,
                  I0 =>  \40222\,
                  I1 =>  \40222\,
                  I2 =>  \40222\,
                  I3 =>  '0' );

  -- Alias \RSTKY/\   
  \=40225\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40225\,
                  I0 =>  \40222\,
                  I1 =>  \40222\,
                  I2 =>  \40222\,
                  I3 =>  '0' );

  -- Alias \IL01\     
  \=40226\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40226\,
                  I0 =>  \S01\,
                  I1 =>  \S01\,
                  I2 =>  \S01\,
                  I3 =>  '0' );

  -- Alias \IL01/\    
  \=40227\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40227\,
                  I0 =>  \S01/\,
                  I1 =>  \S01/\,
                  I2 =>  \S01/\,
                  I3 =>  '0' );

  -- Alias \IL02\     
  \=40228\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40228\,
                  I0 =>  \S02\,
                  I1 =>  \S02\,
                  I2 =>  \S02\,
                  I3 =>  '0' );

  -- Alias \IL02/\    
  \=40229\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40229\,
                  I0 =>  \S02/\,
                  I1 =>  \S02/\,
                  I2 =>  \S02/\,
                  I3 =>  '0' );

  -- Alias \IL03\     
  \=40230\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40230\,
                  I0 =>  \S03\,
                  I1 =>  \S03\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- Alias \IL03/\    
  \=40231\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40231\,
                  I0 =>  \S03/\,
                  I1 =>  \S03/\,
                  I2 =>  \S03/\,
                  I3 =>  '0' );

  -- Alias \IL04\     
  \=40232\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40232\,
                  I0 =>  \S04\,
                  I1 =>  \S04\,
                  I2 =>  \S04\,
                  I3 =>  '0' );

  -- Alias \IL04/\    
  \=40233\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40233\,
                  I0 =>  \S04/\,
                  I1 =>  \S04/\,
                  I2 =>  \S04/\,
                  I3 =>  '0' );

  -- Alias \IL05\     
  \=40234\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40234\,
                  I0 =>  \S05\,
                  I1 =>  \S05\,
                  I2 =>  \S05\,
                  I3 =>  '0' );

  -- Alias \IL05/\    
  \=40235\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40235\,
                  I0 =>  \S05/\,
                  I1 =>  \S05/\,
                  I2 =>  \S05/\,
                  I3 =>  '0' );

  -- Alias \IL06\     
  \=40236\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40236\,
                  I0 =>  \S06\,
                  I1 =>  \S06\,
                  I2 =>  \S06\,
                  I3 =>  '0' );

  -- Alias \IL06/\    
  \=40237\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40237\,
                  I0 =>  \S06/\,
                  I1 =>  \S06/\,
                  I2 =>  \S06/\,
                  I3 =>  '0' );

  -- Alias \IL07\     
  \=40238\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40238\,
                  I0 =>  \S07\,
                  I1 =>  \S07\,
                  I2 =>  \S07\,
                  I3 =>  '0' );

  -- Alias \IL07/\    
  \=40239\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40239\,
                  I0 =>  \S07/\,
                  I1 =>  \S07/\,
                  I2 =>  \S07/\,
                  I3 =>  '0' );

  \=40240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40240\,
                  I0 =>  \STBE\,
                  I1 =>  \1XP10\,
                  I2 =>  \STBF\,
                  I3 =>  '0' );

  -- Alias \CGMC\     
  \=40241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40241\,
                  I0 =>  \40240\,
                  I1 =>  \40258\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40242\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40242\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40242\,
                   R => '0',
                   S => SYSRESET );

  \=40242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40242\,
                  I0 =>  \40241\,
                  I1 =>  \40243\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40243\,
                  I0 =>  \40242\,
                  I1 =>  \40240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40244\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40244\,
                   R => '0',
                   S => SYSRESET );

  \=40244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40244\,
                  I0 =>  \40243\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40245\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \40245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40245\,
                   R => SYSRESET,
                   S => '0' );

  \=40245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40245\,
                  I0 =>  \40244\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40246\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40246\,
                   R => '0',
                   S => SYSRESET );

  \=40246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40246\,
                  I0 =>  \P01\,
                  I1 =>  \40247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40247\,
                  I0 =>  \40246\,
                  I1 =>  \STOP/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40248\,
                  I0 =>  \P04\,
                  I1 =>  \P05/\,
                  I2 =>  '0',
                  I3 => \&40249\ );

  -- Alias \40248\    
  \=40249\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40249\,
                  I0 =>  \40246\,
                  I1 =>  \STOP/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40250\,
                  I0 =>  \STRT2\,
                  I1 =>  \40248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TIMR\     
  \=40251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40251\,
                  I0 =>  \40250\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40253\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40253\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40253\,
                   R => '0',
                   S => SYSRESET );

  \=40253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40253\,
                  I0 =>  \40245\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40254\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \40254\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40254\,
                   R => SYSRESET,
                   S => '0' );

  \=40254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40254\,
                  I0 =>  \40253\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40255\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40255\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40255\,
                   R => '0',
                   S => SYSRESET );

  \=40255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40255\,
                  I0 =>  \40254\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40256\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \40256\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40256\,
                   R => SYSRESET,
                   S => '0' );

  \=40256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40256\,
                  I0 =>  \40255\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40257\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40257\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40257\,
                   R => '0',
                   S => SYSRESET );

  \=40257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40257\,
                  I0 =>  \40256\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40258\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \40258\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40258\,
                   R => SYSRESET,
                   S => '0' );

  \=40258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40258\,
                  I0 =>  \40257\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *******************************************
  -- ***                                     ***
  -- ***  A6 /2 - CROSS POINT GENERATOR II.  ***
  -- ***                                     ***
  -- *******************************************

  \=40302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40302\,
                  I0 =>  \BR1\,
                  I1 =>  \AUG0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40303\,
                  I0 =>  \DIM0/\,
                  I1 =>  \BR12B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40304\,
                  I0 =>  \40302\,
                  I1 =>  \40303\,
                  I2 =>  \INCR0\,
                  I3 => \&40306\ );

  -- Alias \6XP10\    
  \=40305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40305\,
                  I0 =>  \T06/\,
                  I1 =>  \40304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40304\    
  \=40306\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40306\,
                  I0 =>  \PINC\,
                  I1 =>  \40307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40307\,
                  I0 =>  \BR12B/\,
                  I1 =>  \DINC/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40309\,
                  I0 =>  \MINC\,
                  I1 =>  \MCDU\,
                  I2 =>  '0',
                  I3 => \&40315\ );

  \=40310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40310\,
                  I0 =>  \T06/\,
                  I1 =>  \40309\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MONEX/\   
  \=40311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40311\,
                  I0 =>  \40310\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&39104\ );

  \=40312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40312\,
                  I0 =>  \AUG0/\,
                  I1 =>  \BR1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40313\,
                  I0 =>  \DIM0/\,
                  I1 =>  \BR1B2B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40314\,
                  I0 =>  \BR1B2B/\,
                  I1 =>  \DINC/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40309\    
  \=40315\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40315\,
                  I0 =>  \40312\,
                  I1 =>  \40313\,
                  I2 =>  \40314\,
                  I3 =>  '0' );

  \=40317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40317\,
                  I0 =>  \T06/\,
                  I1 =>  \40318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40318\,
                  I0 =>  \PCDU\,
                  I1 =>  \MCDU\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \POUT\     
  \=40320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40320\,
                  I0 =>  \BR1B2B/\,
                  I1 =>  \CDUSTB/\,
                  I2 =>  \DINC/\,
                  I3 =>  '0' );

  -- Alias \MOUT\     
  \=40321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40321\,
                  I0 =>  \BR12B/\,
                  I1 =>  \CDUSTB/\,
                  I2 =>  \DINC/\,
                  I3 =>  '0' );

  -- Alias \ZOUT\     
  \=40322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40322\,
                  I0 =>  \BR2/\,
                  I1 =>  \DINC/\,
                  I2 =>  \CDUSTB/\,
                  I3 =>  '0' );

  \=40323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40323\,
                  I0 =>  \DAS0\,
                  I1 =>  \DAS1\,
                  I2 =>  \MSU0\,
                  I3 =>  '0' );

  \=40324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40324\,
                  I0 =>  \DV4/\,
                  I1 =>  \BR1B2B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40325\,
                  I0 =>  \40324\,
                  I1 =>  \WAND0\,
                  I2 =>  \RAND0\,
                  I3 =>  '0' );

  \=40326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40326\,
                  I0 =>  \40323\,
                  I1 =>  \T07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \7XP7\     
  \=40327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40327\,
                  I0 =>  \T07/\,
                  I1 =>  \40325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WA/\      
  \=40328\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40328\,
                  I0 =>  \40326\,
                  I1 =>  \40327\,
                  I2 =>  \40354\,
                  I3 =>  '0' );

  \=40329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40329\,
                  I0 =>  \WAND0\,
                  I1 =>  \INOTLD\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40330\,
                  I0 =>  \T04/\,
                  I1 =>  \MON/\,
                  I2 =>  \FETCH1\,
                  I3 =>  '0' );

  -- Alias \7XP14\    
  \=40331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40331\,
                  I0 =>  \T07/\,
                  I1 =>  \40329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40333\,
                  I0 =>  \DAS1/\,
                  I1 =>  \T07/\,
                  I2 =>  \BR1B2/\,
                  I3 =>  '0' );

  \=40334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40334\,
                  I0 =>  \DAS1/\,
                  I1 =>  \T07/\,
                  I2 =>  \BR12B/\,
                  I3 =>  '0' );

  \=40335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40335\,
                  I0 =>  \PCDU\,
                  I1 =>  \MCDU\,
                  I2 =>  \SHIFT\,
                  I3 =>  '0' );

  \=40336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40336\,
                  I0 =>  \PRINC\,
                  I1 =>  \PINC\,
                  I2 =>  \MINC\,
                  I3 => \&40339\ );

  \=40337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40337\,
                  I0 =>  \40335\,
                  I1 =>  \T07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40338\,
                  I0 =>  \40336\,
                  I1 =>  \T07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40336\    
  \=40339\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40339\,
                  I0 =>  \DINC\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40340\,
                  I0 =>  \PRINC\,
                  I1 =>  \INKL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WOVR\     
  \=40341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40341\,
                  I0 =>  \40340\,
                  I1 =>  \T07/\,
                  I2 =>  \MON+CH\,
                  I3 =>  '0' );

  -- Alias \WG/\      
  \=40342\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40342\,
                  I0 =>  \40341\,
                  I1 =>  \40346\,
                  I2 =>  '0',
                  I3 => \&34159\ );

  -- Alias \WSC/\     
  \=40343\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40343\,
                  I0 =>  \40341\,
                  I1 =>  \40330\,
                  I2 =>  \40346\,
                  I3 =>  '0' );

  -- Alias \RU/\      
  \=40344\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40344\,
                  I0 =>  \40338\,
                  I1 =>  \40438\,
                  I2 =>  \40354\,
                  I3 => \&40358\ );

  \=40345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40345\,
                  I0 =>  \IC9\,
                  I1 =>  \DXCH0\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40346\,
                  I0 =>  \T07/\,
                  I1 =>  \40345\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RB/\      
  \=40347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40347\,
                  I0 =>  \40346\,
                  I1 =>  \10XP9\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8PP4\     
  \=40348\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40348\,
                  I0 =>  \RUPT1\,
                  I1 =>  \DAS1\,
                  I2 =>  \MSU0\,
                  I3 => \&40417\ );

  -- Alias \8XP4\     
  \=40349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40349\,
                  I0 =>  \T08/\,
                  I1 =>  \8PP4\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8XP10\    
  \=40350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40350\,
                  I0 =>  \T08/\,
                  I1 =>  \RUPT0\,
                  I2 =>  \DAS0\,
                  I3 => \&40351\ );

  -- Alias \40350\    
  \=40351\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40351\,
                  I0 =>  \MP1\,
                  I1 =>  \DV1376\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40352\,
                  I0 =>  \MP3/\,
                  I1 =>  \BR1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40353\,
                  I0 =>  \40352\,
                  I1 =>  \CCS0\,
                  I2 =>  '0',
                  I3 => \&40356\ );

  \=40354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40354\,
                  I0 =>  \T11/\,
                  I1 =>  \40353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40355\,
                  I0 =>  \DAS1/\,
                  I1 =>  \BR2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40353\    
  \=40356\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40356\,
                  I0 =>  \ADS0\,
                  I1 =>  \IC11\,
                  I2 =>  \40355\,
                  I3 =>  '0' );

  -- Alias \RD_BANK\  
  \=40357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40357\,
                  I0 =>  \T06/\,
                  I1 =>  \STFET1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RU/\      
  \=40358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40358\,
                  I0 =>  \RD_BANK\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40401\,
                  I0 =>  \IC6\,
                  I1 =>  \DCA0\,
                  I2 =>  \AD0\,
                  I3 => \&40406\ );

  -- Alias \EXT\      
  \=40402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40402\,
                  I0 =>  \T10/\,
                  I1 =>  \NDXX1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \10XP9\    
  \=40403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40403\,
                  I0 =>  \T10/\,
                  I1 =>  \40401\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40405\,
                  I0 =>  \CCS0/\,
                  I1 =>  \BR1B2B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40401\    
  \=40406\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40406\,
                  I0 =>  \40405\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40407\,
                  I0 =>  \IC6\,
                  I1 =>  \IC7\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40408\,
                  I0 =>  \T10/\,
                  I1 =>  \40407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40409\,
                  I0 =>  \IC7\,
                  I1 =>  \DCS0\,
                  I2 =>  \SU0\,
                  I3 => \&40412\ );

  \=40410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40410\,
                  I0 =>  \T10/\,
                  I1 =>  \40409\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40411\,
                  I0 =>  \CCS0/\,
                  I1 =>  \BR12B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40409\    
  \=40412\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40412\,
                  I0 =>  \40411\,
                  I1 =>  \DV4B1B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=40413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40413\,
                  I0 =>  \T10/\,
                  I1 =>  \MP1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WA/\      
  \=40414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40414\,
                  I0 =>  \40408\,
                  I1 =>  \40438\,
                  I2 =>  \2XP5\,
                  I3 => \&39128\ );

  -- Alias \RC/\      
  \=40415\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40415\,
                  I0 =>  \40410\,
                  I1 =>  \7XP7\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \40424\    
  \=40416\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40416\,
                  I0 =>  \8XP4\,
                  I1 =>  \40413\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \8PP4\     
  \=40417\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40417\,
                  I0 =>  \IC17\,
                  I1 =>  \MASK0\,
                  I2 =>  \IC11\,
                  I3 => \&40418\ );

  -- Alias \8PP4\     
  \=40418\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40418\,
                  I0 =>  \IC6\,
                  I1 =>  \IC7\,
                  I2 =>  \IC9\,
                  I3 =>  '0' );

  -- Alias \RUS/\     
  \=40419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40419\,
                  I0 =>  \7XP9\,
                  I1 =>  \11XP2\,
                  I2 =>  \40337\,
                  I3 =>  '0' );

  -- Alias \RZ/\      
  \=40420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40420\,
                  I0 =>  \8XP4\,
                  I1 =>  \RADRZ\,
                  I2 =>  \9XP1\,
                  I3 => \&39107\ );

  -- Alias \40422\    
  \=40421\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40421\,
                  I0 =>  \2XP8\,
                  I1 =>  \10XP1\,
                  I2 =>  \MP0T10\,
                  I3 =>  '0' );

  \=40422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40422\,
                  I0 =>  \40413\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40421\ );

  -- Alias \ST1\      
  \=40423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40423\,
                  I0 =>  \40422\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ST2/\     
  \=40424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40424\,
                  I0 =>  \RADRZ\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&39228\ );

  -- Alias \ST2\      
  \=40425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40425\,
                  I0 =>  \40424\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:40426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40426\,
                   R => '0',
                   S => SYSRESET );

  \=40426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40426\,
                  I0 =>  \MP0T10\,
                  I1 =>  \40427\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NEAC\     
  \=40427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40427\,
                  I0 =>  \TL15\,
                  I1 =>  \40426\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \2PP1\     
  \=40428\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40428\,
                  I0 =>  \DV0\,
                  I1 =>  \IC15\,
                  I2 =>  \DV1376\,
                  I3 =>  '0' );

  -- Alias \WS/\      
  \=40430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40430\,
                  I0 =>  \8XP10\,
                  I1 =>  \R6\,
                  I2 =>  \R15\,
                  I3 => \&39305\ );

  -- Alias \CI/\      
  \=40431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40431\,
                  I0 =>  \ZIPCI\,
                  I1 =>  \40317\,
                  I2 =>  '0',
                  I3 => \&36440\ );

  \=40432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40432\,
                  I0 =>  \8XP6\,
                  I1 =>  \7XP4\,
                  I2 =>  \10XP8\,
                  I3 => \&40433\ );

  -- Alias \40432\    
  \=40433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40433\,
                  I0 =>  \6XP10\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PONEX\    
  \=40434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40434\,
                  I0 =>  \40432\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \R1C/\     
  \=40435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40435\,
                  I0 =>  \40334\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36453\ );

  -- Alias \RB1/\     
  \=40436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40436\,
                  I0 =>  \40333\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36452\ );

  \=40438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40438\,
                  I0 =>  \DAS1/\,
                  I1 =>  \ADS0\,
                  I2 =>  \T03/\,
                  I3 =>  '0' );

  \:40439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \40439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$40439\,
                   R => '0',
                   S => SYSRESET );

  \=40439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$40439\,
                  I0 =>  \RADRZ\,
                  I1 =>  \40440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PSEUDO\   
  \=40440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \40440\,
                  I0 =>  \40439\,
                  I1 =>  \GOJAM\,
                  I2 =>  \RADRG\,
                  I3 =>  '0' );

  -- Alias \RPTSET\   
  \=40441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&40441\,
                  I0 =>  \40440\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ********************************
  -- ***                          ***
  -- ***  A7 /1 - SERVICE GATES.  ***
  -- ***                          ***
  -- ********************************

  -- Alias \WALSG/\   
  \=33101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33101\,
                  I0 =>  \33102\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WALSG\    
  \=33102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33102\,
                  I0 =>  \ZAP/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33105\,
                  I0 =>  \WY12/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33106\,
                  I0 =>  \WY/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33107\,
                  I0 =>  \33105\,
                  I1 =>  \33106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33108\,
                  I0 =>  \33107\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WYLOG/\   
  \=33109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33109\,
                  I0 =>  \33108\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33111\,
                  I0 =>  \WY/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WYHIG/\   
  \=33112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33112\,
                  I0 =>  \33111\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33113\,
                  I0 =>  \33108\,
                  I1 =>  \33108\,
                  I2 =>  '0',
                  I3 => \&33114\ );

  -- Alias \33113\    
  \=33114\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33114\,
                  I0 =>  \33122\,
                  I1 =>  \33122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWYG\     
  \=33115\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33115\,
                  I0 =>  \33113\,
                  I1 =>  \33113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CUG\      
  \=33116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33116\,
                  I0 =>  \33113\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33122\,
                  I0 =>  \WYD/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \33124\    
  \=33123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33123\,
                  I0 =>  \WYD/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33124\,
                  I0 =>  \SHIFT\,
                  I1 =>  \NEAC\,
                  I2 =>  \33125\,
                  I3 => \&33123\ );

  \=33125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33125\,
                  I0 =>  \L15/\,
                  I1 =>  \PIFL/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WYDG/\    
  \=33126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33126\,
                  I0 =>  \33122\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WYDLOG/\  
  \=33129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33129\,
                  I0 =>  \33124\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33130\,
                  I0 =>  \WB/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WBG/\     
  \=33131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33131\,
                  I0 =>  \33130\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWBG\     
  \=33135\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33135\,
                  I0 =>  \33131\,
                  I1 =>  \33131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CBG\      
  \=33136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33136\,
                  I0 =>  \33131\,
                  I1 =>  \33131\,
                  I2 =>  \33131\,
                  I3 => \&33138\ );

  -- Alias \33136\    
  \=33138\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33138\,
                  I0 =>  \CT/\,
                  I1 =>  \CT/\,
                  I2 =>  \CT/\,
                  I3 =>  '0' );

  -- Alias \MWG\      
  \=33139\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33139\,
                  I0 =>  \WGA/\,
                  I1 =>  \WGA/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WGNORM\   
  \=33140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33140\,
                  I0 =>  \WGA/\,
                  I1 =>  \WT/\,
                  I2 =>  \GINH\,
                  I3 =>  '0' );

  -- Alias \WG1G/\    
  \=33141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33141\,
                  I0 =>  \33140\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33144\,
                  I0 =>  \WGA/\,
                  I1 =>  \WT/\,
                  I2 =>  \SR/\,
                  I3 =>  '0' );

  -- Alias \WG2G/\    
  \=33145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33145\,
                  I0 =>  \33140\,
                  I1 =>  \33144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WG4G/\    
  \=33146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33146\,
                  I0 =>  \33144\,
                  I1 =>  \33149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33149\,
                  I0 =>  \WGA/\,
                  I1 =>  \WT/\,
                  I2 =>  \CYR/\,
                  I3 =>  '0' );

  -- Alias \WG5G/\    
  \=33150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33150\,
                  I0 =>  \33149\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33151\,
                  I0 =>  \WGA/\,
                  I1 =>  \WT/\,
                  I2 =>  \CYL/\,
                  I3 =>  '0' );

  -- Alias \WG3G/\    
  \=33152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33152\,
                  I0 =>  \33151\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33155\,
                  I0 =>  \WGA/\,
                  I1 =>  \WT/\,
                  I2 =>  \EDOP/\,
                  I3 =>  '0' );

  -- Alias \WEDOPG/\  
  \=33156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33156\,
                  I0 =>  \33155\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPSAM\   
  \=33160\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33160\,
                  I0 =>  \PIPPLS/\,
                  I1 =>  \SB2/\,
                  I2 =>  \P04A\,
                  I3 =>  '0' );

  \=33201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33201\,
                  I0 =>  \WT/\,
                  I1 =>  \WZ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WZG/\     
  \=33202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33202\,
                  I0 =>  \33201\,
                  I1 =>  \33204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33204\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWZG\     
  \=33207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33207\,
                  I0 =>  \33202\,
                  I1 =>  \33202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CZG\      
  \=33208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33208\,
                  I0 =>  \33202\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33211\,
                  I0 =>  \WL/\,
                  I1 =>  \WT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33212\,
                  I0 =>  \XB1/\,
                  I1 =>  \XT0/\,
                  I2 =>  \WCHG/\,
                  I3 =>  '0' );

  \=33213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33213\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WLG/\     
  \=33214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33214\,
                  I0 =>  \33211\,
                  I1 =>  \33212\,
                  I2 =>  \33213\,
                  I3 =>  '0' );

  \=33217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33217\,
                  I0 =>  \33213\,
                  I1 =>  \33211\,
                  I2 =>  \33212\,
                  I3 =>  '0' );

  -- Alias \MWLG\     
  \=33218\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33218\,
                  I0 =>  \33217\,
                  I1 =>  \33217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33219\,
                  I0 =>  \33213\,
                  I1 =>  \33211\,
                  I2 =>  \33212\,
                  I3 => \&33220\ );

  -- Alias \33219\    
  \=33220\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33220\,
                  I0 =>  \WALSG\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CLG2G\    
  \=33221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33221\,
                  I0 =>  \33219\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33222\,
                  I0 =>  \33212\,
                  I1 =>  \33211\,
                  I2 =>  \33213\,
                  I3 => \&33223\ );

  -- Alias \33222\    
  \=33223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33223\,
                  I0 =>  \G2LSG\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CLG1G\    
  \=33224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33224\,
                  I0 =>  \CT/\,
                  I1 =>  \33222\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33227\,
                  I0 =>  \WT/\,
                  I1 =>  \WA/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33228\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WAG/\     
  \=33229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33229\,
                  I0 =>  \33227\,
                  I1 =>  \33228\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33232\,
                  I0 =>  \33227\,
                  I1 =>  \33228\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33233\,
                  I0 =>  \33227\,
                  I1 =>  \33228\,
                  I2 =>  \WALSG\,
                  I3 =>  '0' );

  -- Alias \CAG\      
  \=33234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33234\,
                  I0 =>  \33233\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33237\,
                  I0 =>  \WT/\,
                  I1 =>  \WS/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WSG/\     
  \=33238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33238\,
                  I0 =>  \33237\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWSG\     
  \=33241\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33241\,
                  I0 =>  \33238\,
                  I1 =>  \33238\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CSG\      
  \=33242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33242\,
                  I0 =>  \33238\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33244\,
                  I0 =>  \WT/\,
                  I1 =>  \WQ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33245\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33246\,
                  I0 =>  \XB2/\,
                  I1 =>  \XT0/\,
                  I2 =>  \WCHG/\,
                  I3 =>  '0' );

  -- Alias \WQG/\     
  \=33247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33247\,
                  I0 =>  \33245\,
                  I1 =>  \33244\,
                  I2 =>  \33246\,
                  I3 =>  '0' );

  -- Alias \MWQG\     
  \=33251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33251\,
                  I0 =>  \33247\,
                  I1 =>  \33247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CQG\      
  \=33252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33252\,
                  I0 =>  \33247\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWAG\     
  \=33255\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33255\,
                  I0 =>  \33232\,
                  I1 =>  \33232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \P04A\     
  \=33257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33257\,
                  I0 =>  '0',
                  I1 =>  \P04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ********************************
  -- ***                          ***
  -- ***  A7 /2 - SERVICE GATES.  ***
  -- ***                          ***
  -- ********************************

  \=33301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33301\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WEBG/\    
  \=33302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33302\,
                  I0 =>  \33301\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWEBG\    
  \=33303\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33303\,
                  I0 =>  \33302\,
                  I1 =>  \33302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33305\,
                  I0 =>  \33301\,
                  I1 =>  \U2BBK\,
                  I2 =>  \33312\,
                  I3 =>  '0' );

  -- Alias \CEBG\     
  \=33306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33306\,
                  I0 =>  \33305\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33307\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WFBG/\    
  \=33308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33308\,
                  I0 =>  \33312\,
                  I1 =>  \33307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CFBG\     
  \=33310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33310\,
                  I0 =>  \CT/\,
                  I1 =>  \33359\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWFBG\    
  \=33311\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33311\,
                  I0 =>  \33308\,
                  I1 =>  \33308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33312\,
                  I0 =>  \WSCG/\,
                  I1 =>  \XB6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WBBEG/\   
  \=33313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33313\,
                  I0 =>  \33312\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWBBEG\   
  \=33315\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33315\,
                  I0 =>  \33313\,
                  I1 =>  \33313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RGG1\     
  \=33316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33316\,
                  I0 =>  \RT/\,
                  I1 =>  \RG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RGG/\     
  \=33317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33317\,
                  I0 =>  \33316\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRGG\     
  \=33320\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33320\,
                  I0 =>  \33317\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33321\,
                  I0 =>  \RT/\,
                  I1 =>  \RA/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33322\,
                  I0 =>  \XB0/\,
                  I1 =>  \RSCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RAG/\     
  \=33323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33323\,
                  I0 =>  \33321\,
                  I1 =>  \33322\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRAG\     
  \=33326\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33326\,
                  I0 =>  \33323\,
                  I1 =>  \33323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33327\,
                  I0 =>  \RSCG/\,
                  I1 =>  \XB3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \REBG/\    
  \=33328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33328\,
                  I0 =>  \33327\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLG2\     
  \=33329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33329\,
                  I0 =>  \RT/\,
                  I1 =>  \RL/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLG/\     
  \=33330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33330\,
                  I0 =>  \33331\,
                  I1 =>  \33329\,
                  I2 =>  \33333\,
                  I3 =>  '0' );

  -- Alias \RLG1\     
  \=33331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33331\,
                  I0 =>  \RSCG/\,
                  I1 =>  \XB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLG3\     
  \=33333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33333\,
                  I0 =>  \XB1/\,
                  I1 =>  \XT0/\,
                  I2 =>  \RCHG/\,
                  I3 =>  '0' );

  -- Alias \MRLG\     
  \=33335\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33335\,
                  I0 =>  \33330\,
                  I1 =>  \33330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33336\,
                  I0 =>  \RT/\,
                  I1 =>  \RZ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33337\,
                  I0 =>  \XB5/\,
                  I1 =>  \RSCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RZG/\     
  \=33338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33338\,
                  I0 =>  \33337\,
                  I1 =>  \33336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33341\,
                  I0 =>  \RT/\,
                  I1 =>  \RU/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RULOG/\   
  \=33342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33342\,
                  I0 =>  \33345\,
                  I1 =>  \33341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33345\,
                  I0 =>  \RT/\,
                  I1 =>  \RUS/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33346\,
                  I0 =>  \33345\,
                  I1 =>  \33341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRULOG\   
  \=33347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33347\,
                  I0 =>  \33346\,
                  I1 =>  \33346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RUG/\     
  \=33348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33348\,
                  I0 =>  \33341\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RUSG/\    
  \=33349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33349\,
                  I0 =>  \33345\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33350\,
                  I0 =>  \RT/\,
                  I1 =>  \RB/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RBHG/\    
  \=33351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33351\,
                  I0 =>  \33350\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33352\,
                  I0 =>  \RT/\,
                  I1 =>  \33355\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RBLG/\    
  \=33353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33353\,
                  I0 =>  \33350\,
                  I1 =>  \33352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33355\,
                  I0 =>  \RL10BB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI01/\    
  \:33356\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \33356\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$33356\,
                   R => '0',
                   S => SYSRESET );

  \=33356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$33356\,
                  I0 =>  \CIFF\,
                  I1 =>  \CINORM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33359\,
                  I0 =>  \33312\,
                  I1 =>  \U2BBK\,
                  I2 =>  \33307\,
                  I3 =>  '0' );

  \=33401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33401\,
                  I0 =>  \RT/\,
                  I1 =>  \RC/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCG/\     
  \=33402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33402\,
                  I0 =>  \33401\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33405\,
                  I0 =>  \RT/\,
                  I1 =>  \RQ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RQG/\     
  \=33406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33406\,
                  I0 =>  \33405\,
                  I1 =>  \33409\,
                  I2 =>  \33407\,
                  I3 =>  '0' );

  \=33407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33407\,
                  I0 =>  \RSCG/\,
                  I1 =>  \XB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33409\,
                  I0 =>  \XB2/\,
                  I1 =>  \XT0/\,
                  I2 =>  \RCHG/\,
                  I3 =>  '0' );

  \=33411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33411\,
                  I0 =>  \RSCG/\,
                  I1 =>  \XB4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RFBG/\    
  \=33412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33412\,
                  I0 =>  \33411\,
                  I1 =>  \RBBK\,
                  I2 =>  \33413\,
                  I3 =>  '0' );

  \=33413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33413\,
                  I0 =>  \RSCG/\,
                  I1 =>  \XB6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RBBEG/\   
  \=33414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33414\,
                  I0 =>  \33413\,
                  I1 =>  \RBBK\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G2LSG\    
  \=33415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33415\,
                  I0 =>  \TT/\,
                  I1 =>  \ZAP/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G2LSG/\   
  \=33416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33416\,
                  I0 =>  \33415\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33419\,
                  I0 =>  \TT/\,
                  I1 =>  \L2GD/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L2GDG/\   
  \=33420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33420\,
                  I0 =>  \33419\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33423\,
                  I0 =>  \TT/\,
                  I1 =>  \A2X/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A2XG/\    
  \=33424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33424\,
                  I0 =>  \33423\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33427\,
                  I0 =>  \L2GD/\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33428\,
                  I0 =>  \CT/\,
                  I1 =>  \WG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=33429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33429\,
                  I0 =>  \33427\,
                  I1 =>  \33428\,
                  I2 =>  \CGMC\,
                  I3 =>  '0' );

  -- Alias \CGG\      
  \=33430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33430\,
                  I0 =>  \33429\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT0\      
  \=33433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33433\,
                  I0 =>  \EAD11\,
                  I1 =>  \EAD10\,
                  I2 =>  \EAD09\,
                  I3 =>  '0' );

  -- Alias \YT0/\     
  \=33434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33434\,
                  I0 =>  \33433\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT0E\     
  \=33435\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33435\,
                  I0 =>  \33434\,
                  I1 =>  \33434\,
                  I2 =>  \33434\,
                  I3 =>  '0' );

  -- Alias \YT1\      
  \=33436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33436\,
                  I0 =>  \EAD11\,
                  I1 =>  \EAD10\,
                  I2 =>  \EAD09/\,
                  I3 =>  '0' );

  -- Alias \YT1/\     
  \=33437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33437\,
                  I0 =>  \33436\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT1E\     
  \=33438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33438\,
                  I0 =>  \33437\,
                  I1 =>  \33437\,
                  I2 =>  \33437\,
                  I3 =>  '0' );

  -- Alias \YT2\      
  \=33439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33439\,
                  I0 =>  \EAD11\,
                  I1 =>  \EAD10/\,
                  I2 =>  \EAD09\,
                  I3 =>  '0' );

  -- Alias \YT2/\     
  \=33440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33440\,
                  I0 =>  \33439\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT2E\     
  \=33441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33441\,
                  I0 =>  \33440\,
                  I1 =>  \33440\,
                  I2 =>  \33440\,
                  I3 =>  '0' );

  -- Alias \YT3\      
  \=33442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33442\,
                  I0 =>  \EAD11\,
                  I1 =>  \EAD10/\,
                  I2 =>  \EAD09/\,
                  I3 =>  '0' );

  -- Alias \YT3/\     
  \=33443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33443\,
                  I0 =>  \33442\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT3E\     
  \=33444\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33444\,
                  I0 =>  \33443\,
                  I1 =>  \33443\,
                  I2 =>  \33443\,
                  I3 =>  '0' );

  -- Alias \YT4\      
  \=33445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33445\,
                  I0 =>  \EAD11/\,
                  I1 =>  \EAD10\,
                  I2 =>  \EAD09\,
                  I3 =>  '0' );

  -- Alias \YT4/\     
  \=33446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33446\,
                  I0 =>  \33445\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT4E\     
  \=33447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33447\,
                  I0 =>  \33446\,
                  I1 =>  \33446\,
                  I2 =>  \33446\,
                  I3 =>  '0' );

  -- Alias \YT5\      
  \=33448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33448\,
                  I0 =>  \EAD11/\,
                  I1 =>  \EAD10\,
                  I2 =>  \EAD09/\,
                  I3 =>  '0' );

  -- Alias \YT5/\     
  \=33449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33449\,
                  I0 =>  \33448\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT5E\     
  \=33450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33450\,
                  I0 =>  \33449\,
                  I1 =>  \33449\,
                  I2 =>  \33449\,
                  I3 =>  '0' );

  -- Alias \YT6\      
  \=33451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33451\,
                  I0 =>  \EAD11/\,
                  I1 =>  \EAD10/\,
                  I2 =>  \EAD09\,
                  I3 =>  '0' );

  -- Alias \YT6/\     
  \=33452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33452\,
                  I0 =>  \33451\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT6E\     
  \=33453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33453\,
                  I0 =>  \33452\,
                  I1 =>  \33452\,
                  I2 =>  \33452\,
                  I3 =>  '0' );

  -- Alias \YT7\      
  \=33454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33454\,
                  I0 =>  \EAD11/\,
                  I1 =>  \EAD09/\,
                  I2 =>  \EAD10/\,
                  I3 =>  '0' );

  -- Alias \YT7/\     
  \=33455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33455\,
                  I0 =>  \33454\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YT7E\     
  \=33456\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&33456\,
                  I0 =>  \33455\,
                  I1 =>  \33455\,
                  I2 =>  \33455\,
                  I3 =>  '0' );

  -- Alias \CINORM\   
  \=33457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33457\,
                  I0 =>  \NEAC\,
                  I1 =>  \EAC/\,
                  I2 =>  '0',
                  I3 => \&37360\ );

  \:33458\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \33458\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$33458\,
                   R => '0',
                   S => SYSRESET );

  \=33458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$33458\,
                  I0 =>  \CI\,
                  I1 =>  \33459\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CIFF\     
  \=33459\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33459\,
                  I0 =>  \33458\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RBBK\     
  \=33460\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \33460\,
                  I0 =>  \T10/\,
                  I1 =>  \STFET1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A8 /1 - 4 BIT MODULE (1 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO04\     
  \=51101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51101\,
                  I0 =>  \XUY03/\,
                  I1 =>  \51110\,
                  I2 =>  \CI01/\,
                  I3 => \&51201\ );

  \=51102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51102\,
                  I0 =>  \A2XG/\,
                  I1 =>  \51120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51103\,
                   R => '0',
                   S => SYSRESET );

  \=51103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51103\,
                  I0 =>  \PONEX\,
                  I1 =>  \51102\,
                  I2 =>  \51104\,
                  I3 =>  '0' );

  \=51104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51104\,
                  I0 =>  \51103\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=51105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51105\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51106\,
                  I0 =>  \WL16/\,
                  I1 =>  \WYDLOG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51107\,
                   R => '0',
                   S => SYSRESET );

  \=51107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51107\,
                  I0 =>  \51105\,
                  I1 =>  \51106\,
                  I2 =>  \51108\,
                  I3 =>  '0' );

  \=51108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51108\,
                  I0 =>  \51107\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51109\,
                  I0 =>  \51103\,
                  I1 =>  \51107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY01/\   
  \=51110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51110\,
                  I0 =>  \51104\,
                  I1 =>  \51108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51111\,
                  I0 =>  \CI01/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA01/\  
  \=51112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51112\,
                  I0 =>  \51109\,
                  I1 =>  \CI01/\,
                  I2 =>  \51110\,
                  I3 =>  '0' );

  \=51113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51113\,
                  I0 =>  \51109\,
                  I1 =>  \51110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI02/\    
  \=51114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51114\,
                  I0 =>  \51109\,
                  I1 =>  \51112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB01/\  
  \=51115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51115\,
                  I0 =>  \51113\,
                  I1 =>  \51111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51117\,
                  I0 =>  \51112\,
                  I1 =>  \51115\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=51118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51118\,
                  I0 =>  \WAG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51119\,
                  I0 =>  \WL03/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A01/\     
  \:51120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51120\,
                   R => '0',
                   S => SYSRESET );

  \=51120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51120\,
                  I0 =>  \51118\,
                  I1 =>  \51119\,
                  I2 =>  \51121\,
                  I3 =>  '0' );

  \=51121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51121\,
                  I0 =>  \51120\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51122\,
                  I0 =>  \RAG/\,
                  I1 =>  \51120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51157\    
  \=51123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51123\,
                  I0 =>  \51117\,
                  I1 =>  \51122\,
                  I2 =>  \CH01\,
                  I3 => \&51133\ );

  \=51124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51124\,
                  I0 =>  \WLG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51125\,
                  I0 =>  \G04/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L01/\     
  \:51126\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51126\,
                   R => '0',
                   S => SYSRESET );

  \=51126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51126\,
                  I0 =>  \51124\,
                  I1 =>  \51125\,
                  I2 =>  \51127\,
                  I3 =>  '0' );

  \=51127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51127\,
                  I0 =>  \51126\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51128\,
                  I0 =>  \RLG/\,
                  I1 =>  \51126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51129\,
                  I0 =>  \WQG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51130\,
                   R => '0',
                   S => SYSRESET );

  \=51130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51130\,
                  I0 =>  \51129\,
                  I1 =>  \51131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51131\,
                  I0 =>  \51130\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51132\,
                  I0 =>  \RQG/\,
                  I1 =>  \51130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51157\    
  \=51133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51133\,
                  I0 =>  \51128\,
                  I1 =>  \51132\,
                  I2 =>  \51137\,
                  I3 => \&51158\ );

  \=51134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51134\,
                  I0 =>  \WZG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z01/\     
  \:51135\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51135\,
                   R => '0',
                   S => SYSRESET );

  \=51135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51135\,
                  I0 =>  \51134\,
                  I1 =>  \51136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51136\,
                  I0 =>  \51135\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51137\,
                  I0 =>  \RZG/\,
                  I1 =>  \51135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51138\,
                  I0 =>  \WBG/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51139\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51139\,
                   R => '0',
                   S => SYSRESET );

  \=51139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51139\,
                  I0 =>  \51138\,
                  I1 =>  \51140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51140\,
                  I0 =>  \51139\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51141\,
                  I0 =>  \RBLG/\,
                  I1 =>  \51139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51142\,
                  I0 =>  \51140\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51143\,
                  I0 =>  \WL16/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51144\,
                  I0 =>  \WL02/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51145\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \MCRO/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51146\,
                  I0 =>  \WG1G/\,
                  I1 =>  \51154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51148\    
  \=51147\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51147\,
                  I0 =>  \SA01\,
                  I1 =>  \51143\,
                  I2 =>  \51144\,
                  I3 => \&51162\ );

  -- Alias \G01/\     
  \:51148\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51148\,
                   R => '0',
                   S => SYSRESET );

  \=51148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51148\,
                  I0 =>  \51145\,
                  I1 =>  \51146\,
                  I2 =>  \51149\,
                  I3 => \&51147\ );

  -- Alias \G01\      
  \=51149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51149\,
                  I0 =>  \51148\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM01\    
  \=51150\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51150\,
                  I0 =>  \51148\,
                  I1 =>  \51148\,
                  I2 =>  \51148\,
                  I3 =>  '0' );

  \=51151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51151\,
                  I0 =>  \RGG/\,
                  I1 =>  \51148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL01\     
  \=51152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51152\,
                  I0 =>  \51157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL01\    
  \=51153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51153\,
                  I0 =>  \51157\,
                  I1 =>  \51157\,
                  I2 =>  \51157\,
                  I3 =>  '0' );

  -- Alias \WL01/\    
  \=51154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51154\,
                  I0 =>  \51152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL01/\    
  \=51157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51157\,
                  I0 =>  \51141\,
                  I1 =>  \51142\,
                  I2 =>  \51151\,
                  I3 => \&51123\ );

  -- Alias \51157\    
  \=51158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51158\,
                  I0 =>  \MDT01\,
                  I1 =>  \RB1\,
                  I2 =>  \R15\,
                  I3 => \&35460\ );

  -- Alias \CLEARA\   
  \=51161\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51161\,
                  I0 =>  \SETAB/\,
                  I1 =>  \S08A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G01/\     
  \=51162\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51162\,
                  I0 =>  \G01ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G02/\     
  \=51163\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51163\,
                  I0 =>  \G02ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51247\ );

  -- Alias \CO04\     
  \=51201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51201\,
                  I0 =>  \XUY04/\,
                  I1 =>  \51210\,
                  I2 =>  '0',
                  I3 => \&53462\ );

  \=51202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51202\,
                  I0 =>  \A2XG/\,
                  I1 =>  \51220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51203\,
                   R => '0',
                   S => SYSRESET );

  \=51203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51203\,
                  I0 =>  \TWOX\,
                  I1 =>  \51202\,
                  I2 =>  \51204\,
                  I3 =>  '0' );

  \=51204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51204\,
                  I0 =>  \51203\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=51205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51205\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51206\,
                  I0 =>  \WL01/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51207\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51207\,
                   R => '0',
                   S => SYSRESET );

  \=51207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51207\,
                  I0 =>  \51205\,
                  I1 =>  \51206\,
                  I2 =>  \51208\,
                  I3 =>  '0' );

  \=51208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51208\,
                  I0 =>  \51207\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51209\,
                  I0 =>  \51203\,
                  I1 =>  \51207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY02/\   
  \=51210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51210\,
                  I0 =>  \51204\,
                  I1 =>  \51208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51211\,
                  I0 =>  \CI02/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA02/\  
  \=51212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51212\,
                  I0 =>  \51209\,
                  I1 =>  \51210\,
                  I2 =>  \CI02/\,
                  I3 => \&54162\ );

  \=51213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51213\,
                  I0 =>  \51209\,
                  I1 =>  \51210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI03/\    
  \=51214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51214\,
                  I0 =>  \51209\,
                  I1 =>  \51212\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB02/\  
  \=51215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51215\,
                  I0 =>  \51213\,
                  I1 =>  \51211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51217\,
                  I0 =>  \51212\,
                  I1 =>  \51215\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=51218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51218\,
                  I0 =>  \WAG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51219\,
                  I0 =>  \WL04/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A02/\     
  \:51220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51220\,
                   R => '0',
                   S => SYSRESET );

  \=51220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51220\,
                  I0 =>  \51218\,
                  I1 =>  \51219\,
                  I2 =>  \51221\,
                  I3 =>  '0' );

  \=51221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51221\,
                  I0 =>  \51220\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51222\,
                  I0 =>  \RAG/\,
                  I1 =>  \51220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51257\    
  \=51223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51223\,
                  I0 =>  \51217\,
                  I1 =>  \51222\,
                  I2 =>  \CH02\,
                  I3 => \&51233\ );

  \=51224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51224\,
                  I0 =>  \WLG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51225\,
                  I0 =>  \G05/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L02/\     
  \:51226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51226\,
                   R => '0',
                   S => SYSRESET );

  \=51226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51226\,
                  I0 =>  \51224\,
                  I1 =>  \51225\,
                  I2 =>  \51227\,
                  I3 =>  '0' );

  \=51227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51227\,
                  I0 =>  \51226\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51228\,
                  I0 =>  \RLG/\,
                  I1 =>  \51226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51229\,
                  I0 =>  \WQG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51230\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51230\,
                   R => '0',
                   S => SYSRESET );

  \=51230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51230\,
                  I0 =>  \51229\,
                  I1 =>  \51231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51231\,
                  I0 =>  \51230\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51232\,
                  I0 =>  \RQG/\,
                  I1 =>  \51230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51257\    
  \=51233\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51233\,
                  I0 =>  \51228\,
                  I1 =>  \51232\,
                  I2 =>  \51237\,
                  I3 => \&51258\ );

  \=51234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51234\,
                  I0 =>  \WZG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z02/\     
  \:51235\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51235\,
                   R => '0',
                   S => SYSRESET );

  \=51235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51235\,
                  I0 =>  \51234\,
                  I1 =>  \51236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51236\,
                  I0 =>  \51235\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51237\,
                  I0 =>  \RZG/\,
                  I1 =>  \51235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51238\,
                  I0 =>  \WBG/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51239\,
                   R => '0',
                   S => SYSRESET );

  \=51239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51239\,
                  I0 =>  \51238\,
                  I1 =>  \51240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51240\,
                  I0 =>  \51239\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51241\,
                  I0 =>  \RBLG/\,
                  I1 =>  \51239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51242\,
                  I0 =>  \51240\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51243\,
                  I0 =>  \WL01/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51244\,
                  I0 =>  \WL03/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51245\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51246\,
                  I0 =>  \WG1G/\,
                  I1 =>  \51254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51248\    
  \=51247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51247\,
                  I0 =>  \SA02\,
                  I1 =>  \51243\,
                  I2 =>  \51244\,
                  I3 =>  '0' );

  -- Alias \G02/\     
  \:51248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51248\,
                   R => '0',
                   S => SYSRESET );

  \=51248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51248\,
                  I0 =>  \51245\,
                  I1 =>  \51246\,
                  I2 =>  \51249\,
                  I3 => \&51163\ );

  -- Alias \G02\      
  \=51249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51249\,
                  I0 =>  \51248\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM02\    
  \=51250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51250\,
                  I0 =>  \51248\,
                  I1 =>  \51248\,
                  I2 =>  \51248\,
                  I3 =>  '0' );

  \=51251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51251\,
                  I0 =>  \RGG/\,
                  I1 =>  \51248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL02\     
  \=51252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51252\,
                  I0 =>  \51257\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL02\    
  \=51253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51253\,
                  I0 =>  \51257\,
                  I1 =>  \51257\,
                  I2 =>  \51257\,
                  I3 =>  '0' );

  -- Alias \WL02/\    
  \=51254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51254\,
                  I0 =>  \51252\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL02/\    
  \=51257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51257\,
                  I0 =>  \51241\,
                  I1 =>  \51242\,
                  I2 =>  \51251\,
                  I3 => \&51223\ );

  -- Alias \51257\    
  \=51258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51258\,
                  I0 =>  \MDT02\,
                  I1 =>  \R1C\,
                  I2 =>  \RB2\,
                  I3 => \&35360\ );

  -- Alias \S08A/\    
  \=51261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51261\,
                  I0 =>  \S08\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S08A\     
  \=51262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51262\,
                  I0 =>  \S08/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G03/\     
  \=51263\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51263\,
                  I0 =>  \G03ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51447\ );

  -- ****************************************
  -- ***                                  ***
  -- ***  A8 /2 - 4 BIT MODULE (1 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO06\     
  \=51301\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51301\,
                  I0 =>  \XUY06/\,
                  I1 =>  \51310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51302\,
                  I0 =>  \A2XG/\,
                  I1 =>  \51320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51303\,
                   R => '0',
                   S => SYSRESET );

  \=51303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51303\,
                  I0 =>  \MONEX\,
                  I1 =>  \51302\,
                  I2 =>  \51304\,
                  I3 =>  '0' );

  \=51304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51304\,
                  I0 =>  \51303\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=51305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51305\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51306\,
                  I0 =>  \WL03/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51307\,
                   R => '0',
                   S => SYSRESET );

  \=51307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51307\,
                  I0 =>  \51305\,
                  I1 =>  \51306\,
                  I2 =>  \51308\,
                  I3 =>  '0' );

  \=51308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51308\,
                  I0 =>  \51307\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51309\,
                  I0 =>  \51303\,
                  I1 =>  \51307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY04/\   
  \=51310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51310\,
                  I0 =>  \51304\,
                  I1 =>  \51308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51311\,
                  I0 =>  \CI04/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA04/\  
  \=51312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51312\,
                  I0 =>  \51309\,
                  I1 =>  \51310\,
                  I2 =>  \CI04/\,
                  I3 => \&54163\ );

  \=51313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51313\,
                  I0 =>  \51309\,
                  I1 =>  \51310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI05/\    
  \=51314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51314\,
                  I0 =>  \51309\,
                  I1 =>  \51312\,
                  I2 =>  \CO04\,
                  I3 =>  '0' );

  -- Alias \SUMB04/\  
  \=51315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51315\,
                  I0 =>  \51313\,
                  I1 =>  \51311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51317\,
                  I0 =>  \51312\,
                  I1 =>  \51315\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=51318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51318\,
                  I0 =>  \WAG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51319\,
                  I0 =>  \WL06/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A04/\     
  \:51320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51320\,
                   R => '0',
                   S => SYSRESET );

  \=51320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51320\,
                  I0 =>  \51318\,
                  I1 =>  \51319\,
                  I2 =>  \51321\,
                  I3 =>  '0' );

  \=51321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51321\,
                  I0 =>  \51320\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51322\,
                  I0 =>  \RAG/\,
                  I1 =>  \51320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51357\    
  \=51323\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51323\,
                  I0 =>  \51317\,
                  I1 =>  \51322\,
                  I2 =>  \CH04\,
                  I3 => \&51333\ );

  \=51324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51324\,
                  I0 =>  \WLG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51325\,
                  I0 =>  \G07/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L04/\     
  \:51326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51326\,
                   R => '0',
                   S => SYSRESET );

  \=51326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51326\,
                  I0 =>  \51324\,
                  I1 =>  \51325\,
                  I2 =>  \51327\,
                  I3 =>  '0' );

  \=51327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51327\,
                  I0 =>  \51326\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51328\,
                  I0 =>  \RLG/\,
                  I1 =>  \51326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51329\,
                  I0 =>  \WQG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51330\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51330\,
                   R => '0',
                   S => SYSRESET );

  \=51330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51330\,
                  I0 =>  \51329\,
                  I1 =>  \51331\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51331\,
                  I0 =>  \51330\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51332\,
                  I0 =>  \RQG/\,
                  I1 =>  \51330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51357\    
  \=51333\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51333\,
                  I0 =>  \51328\,
                  I1 =>  \51332\,
                  I2 =>  \51337\,
                  I3 => \&51358\ );

  \=51334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51334\,
                  I0 =>  \WZG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z04/\     
  \:51335\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51335\,
                   R => '0',
                   S => SYSRESET );

  \=51335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51335\,
                  I0 =>  \51334\,
                  I1 =>  \51336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51336\,
                  I0 =>  \51335\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51337\,
                  I0 =>  \RZG/\,
                  I1 =>  \51335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51338\,
                  I0 =>  \WBG/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51339\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51339\,
                   R => '0',
                   S => SYSRESET );

  \=51339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51339\,
                  I0 =>  \51338\,
                  I1 =>  \51340\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51340\,
                  I0 =>  \51339\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51341\,
                  I0 =>  \RBLG/\,
                  I1 =>  \51339\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51342\,
                  I0 =>  \51340\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51343\,
                  I0 =>  \WL03/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51344\,
                  I0 =>  \WL05/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51345\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51346\,
                  I0 =>  \WG1G/\,
                  I1 =>  \51354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51348\    
  \=51347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51347\,
                  I0 =>  \SA04\,
                  I1 =>  \51343\,
                  I2 =>  \51344\,
                  I3 => \&51462\ );

  -- Alias \G04/\     
  \:51348\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51348\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51348\,
                   R => '0',
                   S => SYSRESET );

  \=51348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51348\,
                  I0 =>  \51345\,
                  I1 =>  \51346\,
                  I2 =>  \51349\,
                  I3 => \&51347\ );

  -- Alias \G04\      
  \=51349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51349\,
                  I0 =>  \51348\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM04\    
  \=51350\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51350\,
                  I0 =>  \51348\,
                  I1 =>  \51348\,
                  I2 =>  \51348\,
                  I3 =>  '0' );

  \=51351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51351\,
                  I0 =>  \RGG/\,
                  I1 =>  \51348\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL04\     
  \=51352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51352\,
                  I0 =>  \51357\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL04\    
  \=51353\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51353\,
                  I0 =>  \51357\,
                  I1 =>  \51357\,
                  I2 =>  \51357\,
                  I3 =>  '0' );

  -- Alias \WL04/\    
  \=51354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51354\,
                  I0 =>  \51352\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL04/\    
  \=51357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51357\,
                  I0 =>  \51341\,
                  I1 =>  \51342\,
                  I2 =>  \51351\,
                  I3 => \&51323\ );

  -- Alias \51357\    
  \=51358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51358\,
                  I0 =>  \MDT04\,
                  I1 =>  \R1C\,
                  I2 =>  \R15\,
                  I3 => \&34451\ );

  -- Alias \CLEARC\   
  \=51361\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51361\,
                  I0 =>  \SETCD/\,
                  I1 =>  \S08A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CLEARD\   
  \=51362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51362\,
                  I0 =>  \SETCD/\,
                  I1 =>  \S08A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G06/\     
  \=51363\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51363\,
                  I0 =>  \G06ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52247\ );

  -- Alias \CO06\     
  \=51401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51401\,
                  I0 =>  \XUY05/\,
                  I1 =>  \51410\,
                  I2 =>  \CI03/\,
                  I3 => \&51301\ );

  \=51402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51402\,
                  I0 =>  \A2XG/\,
                  I1 =>  \51420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51403\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51403\,
                   R => '0',
                   S => SYSRESET );

  \=51403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51403\,
                  I0 =>  \MONEX\,
                  I1 =>  \51402\,
                  I2 =>  \51404\,
                  I3 =>  '0' );

  \=51404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51404\,
                  I0 =>  \51403\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=51405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51405\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51406\,
                  I0 =>  \WL02/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51407\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51407\,
                   R => '0',
                   S => SYSRESET );

  \=51407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51407\,
                  I0 =>  \51405\,
                  I1 =>  \51406\,
                  I2 =>  \51408\,
                  I3 =>  '0' );

  \=51408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51408\,
                  I0 =>  \51407\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51409\,
                  I0 =>  \51403\,
                  I1 =>  \51407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY03/\   
  \=51410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51410\,
                  I0 =>  \51404\,
                  I1 =>  \51408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51411\,
                  I0 =>  \CI03/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA03/\  
  \=51412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51412\,
                  I0 =>  \51409\,
                  I1 =>  \CI03/\,
                  I2 =>  \51410\,
                  I3 =>  '0' );

  \=51413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51413\,
                  I0 =>  \51409\,
                  I1 =>  \51410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI04/\    
  \=51414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51414\,
                  I0 =>  \51409\,
                  I1 =>  \51412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB03/\  
  \=51415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51415\,
                  I0 =>  \51413\,
                  I1 =>  \51411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51417\,
                  I0 =>  \51412\,
                  I1 =>  \51415\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=51418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51418\,
                  I0 =>  \WAG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51419\,
                  I0 =>  \WL05/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A03/\     
  \:51420\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51420\,
                   R => '0',
                   S => SYSRESET );

  \=51420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51420\,
                  I0 =>  \51418\,
                  I1 =>  \51419\,
                  I2 =>  \51421\,
                  I3 =>  '0' );

  \=51421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51421\,
                  I0 =>  \51420\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51422\,
                  I0 =>  \RAG/\,
                  I1 =>  \51420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51457\    
  \=51423\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51423\,
                  I0 =>  \51417\,
                  I1 =>  \51422\,
                  I2 =>  \CH03\,
                  I3 => \&51433\ );

  \=51424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51424\,
                  I0 =>  \WLG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51425\,
                  I0 =>  \G06/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L03/\     
  \:51426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51426\,
                   R => '0',
                   S => SYSRESET );

  \=51426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51426\,
                  I0 =>  \51424\,
                  I1 =>  \51425\,
                  I2 =>  \51427\,
                  I3 =>  '0' );

  \=51427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51427\,
                  I0 =>  \51426\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51428\,
                  I0 =>  \RLG/\,
                  I1 =>  \51426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51429\,
                  I0 =>  \WQG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51430\,
                   R => '0',
                   S => SYSRESET );

  \=51430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51430\,
                  I0 =>  \51429\,
                  I1 =>  \51431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51431\,
                  I0 =>  \51430\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51432\,
                  I0 =>  \RQG/\,
                  I1 =>  \51430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51457\    
  \=51433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51433\,
                  I0 =>  \51428\,
                  I1 =>  \51432\,
                  I2 =>  \51437\,
                  I3 => \&51458\ );

  \=51434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51434\,
                  I0 =>  \WZG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z03/\     
  \:51435\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51435\,
                   R => '0',
                   S => SYSRESET );

  \=51435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51435\,
                  I0 =>  \51434\,
                  I1 =>  \51436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51436\,
                  I0 =>  \51435\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51437\,
                  I0 =>  \RZG/\,
                  I1 =>  \51435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51438\,
                  I0 =>  \WBG/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:51439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51439\,
                   R => '0',
                   S => SYSRESET );

  \=51439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51439\,
                  I0 =>  \51438\,
                  I1 =>  \51440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51440\,
                  I0 =>  \51439\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51441\,
                  I0 =>  \RBLG/\,
                  I1 =>  \51439\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51442\,
                  I0 =>  \51440\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51443\,
                  I0 =>  \WL02/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51444\,
                  I0 =>  \WL04/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51445\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=51446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51446\,
                  I0 =>  \WG1G/\,
                  I1 =>  \51454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \51448\    
  \=51447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51447\,
                  I0 =>  \SA03\,
                  I1 =>  \51443\,
                  I2 =>  \51444\,
                  I3 =>  '0' );

  -- Alias \G03/\     
  \:51448\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \51448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$51448\,
                   R => '0',
                   S => SYSRESET );

  \=51448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$51448\,
                  I0 =>  \51445\,
                  I1 =>  \51446\,
                  I2 =>  \51449\,
                  I3 => \&51263\ );

  -- Alias \G03\      
  \=51449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51449\,
                  I0 =>  \51448\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM03\    
  \=51450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51450\,
                  I0 =>  \51448\,
                  I1 =>  \51448\,
                  I2 =>  \51448\,
                  I3 =>  '0' );

  \=51451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51451\,
                  I0 =>  \RGG/\,
                  I1 =>  \51448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL03\     
  \=51452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51452\,
                  I0 =>  \51457\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL03\    
  \=51453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51453\,
                  I0 =>  \51457\,
                  I1 =>  \51457\,
                  I2 =>  \51457\,
                  I3 =>  '0' );

  -- Alias \WL03/\    
  \=51454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51454\,
                  I0 =>  \51452\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL03/\    
  \=51457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51457\,
                  I0 =>  \51441\,
                  I1 =>  \51442\,
                  I2 =>  \51451\,
                  I3 => \&51423\ );

  -- Alias \51457\    
  \=51458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51458\,
                  I0 =>  \MDT03\,
                  I1 =>  \R1C\,
                  I2 =>  \R15\,
                  I3 => \&34450\ );

  -- Alias \CLEARB\   
  \=51461\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \51461\,
                  I0 =>  \SETAB/\,
                  I1 =>  \S08A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G04/\     
  \=51462\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51462\,
                  I0 =>  \G04ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G05/\     
  \=51463\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&51463\,
                  I0 =>  \G05ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52147\ );

  -- ****************************************
  -- ***                                  ***
  -- ***  A9 /1 - 4 BIT MODULE (2 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO08\     
  \=52101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52101\,
                  I0 =>  \XUY07/\,
                  I1 =>  \52110\,
                  I2 =>  \CI05/\,
                  I3 => \&52201\ );

  \=52102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52102\,
                  I0 =>  \A2XG/\,
                  I1 =>  \52120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52103\,
                   R => '0',
                   S => SYSRESET );

  \=52103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52103\,
                  I0 =>  \MONEX\,
                  I1 =>  \52102\,
                  I2 =>  \52104\,
                  I3 =>  '0' );

  \=52104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52104\,
                  I0 =>  \52103\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=52105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52105\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52106\,
                  I0 =>  \WL04/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52107\,
                   R => '0',
                   S => SYSRESET );

  \=52107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52107\,
                  I0 =>  \52105\,
                  I1 =>  \52106\,
                  I2 =>  \52108\,
                  I3 =>  '0' );

  \=52108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52108\,
                  I0 =>  \52107\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52109\,
                  I0 =>  \52103\,
                  I1 =>  \52107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY05/\   
  \=52110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52110\,
                  I0 =>  \52104\,
                  I1 =>  \52108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52111\,
                  I0 =>  \CI05/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA05/\  
  \=52112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52112\,
                  I0 =>  \52109\,
                  I1 =>  \CI05/\,
                  I2 =>  \52110\,
                  I3 =>  '0' );

  \=52113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52113\,
                  I0 =>  \52109\,
                  I1 =>  \52110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI06/\    
  \=52114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52114\,
                  I0 =>  \52109\,
                  I1 =>  \52112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB05/\  
  \=52115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52115\,
                  I0 =>  \52113\,
                  I1 =>  \52111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52117\,
                  I0 =>  \52112\,
                  I1 =>  \52115\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=52118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52118\,
                  I0 =>  \WAG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52119\,
                  I0 =>  \WL07/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A05/\     
  \:52120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52120\,
                   R => '0',
                   S => SYSRESET );

  \=52120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52120\,
                  I0 =>  \52118\,
                  I1 =>  \52119\,
                  I2 =>  \52121\,
                  I3 =>  '0' );

  \=52121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52121\,
                  I0 =>  \52120\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52122\,
                  I0 =>  \RAG/\,
                  I1 =>  \52120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52157\    
  \=52123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52123\,
                  I0 =>  \52117\,
                  I1 =>  \52122\,
                  I2 =>  \CH05\,
                  I3 => \&52133\ );

  \=52124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52124\,
                  I0 =>  \WLG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52125\,
                  I0 =>  \G08/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L05/\     
  \:52126\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52126\,
                   R => '0',
                   S => SYSRESET );

  \=52126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52126\,
                  I0 =>  \52124\,
                  I1 =>  \52125\,
                  I2 =>  \52127\,
                  I3 =>  '0' );

  \=52127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52127\,
                  I0 =>  \52126\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52128\,
                  I0 =>  \RLG/\,
                  I1 =>  \52126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52129\,
                  I0 =>  \WQG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52130\,
                   R => '0',
                   S => SYSRESET );

  \=52130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52130\,
                  I0 =>  \52129\,
                  I1 =>  \52131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52131\,
                  I0 =>  \52130\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52132\,
                  I0 =>  \RQG/\,
                  I1 =>  \52130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52157\    
  \=52133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52133\,
                  I0 =>  \52128\,
                  I1 =>  \52132\,
                  I2 =>  \52137\,
                  I3 => \&52158\ );

  \=52134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52134\,
                  I0 =>  \WZG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z05/\     
  \:52135\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52135\,
                   R => '0',
                   S => SYSRESET );

  \=52135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52135\,
                  I0 =>  \52134\,
                  I1 =>  \52136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52136\,
                  I0 =>  \52135\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52137\,
                  I0 =>  \RZG/\,
                  I1 =>  \52135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52138\,
                  I0 =>  \WBG/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52139\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52139\,
                   R => '0',
                   S => SYSRESET );

  \=52139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52139\,
                  I0 =>  \52138\,
                  I1 =>  \52140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52140\,
                  I0 =>  \52139\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52141\,
                  I0 =>  \RBLG/\,
                  I1 =>  \52139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52142\,
                  I0 =>  \52140\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52143\,
                  I0 =>  \WL04/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52144\,
                  I0 =>  \WL06/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52145\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52146\,
                  I0 =>  \WG1G/\,
                  I1 =>  \52154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52148\    
  \=52147\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52147\,
                  I0 =>  \SA05\,
                  I1 =>  \52143\,
                  I2 =>  \52144\,
                  I3 =>  '0' );

  -- Alias \G05/\     
  \:52148\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52148\,
                   R => '0',
                   S => SYSRESET );

  \=52148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52148\,
                  I0 =>  \52145\,
                  I1 =>  \52146\,
                  I2 =>  \52149\,
                  I3 => \&51463\ );

  -- Alias \G05\      
  \=52149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52149\,
                  I0 =>  \52148\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM05\    
  \=52150\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52150\,
                  I0 =>  \52148\,
                  I1 =>  \52148\,
                  I2 =>  \52148\,
                  I3 =>  '0' );

  \=52151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52151\,
                  I0 =>  \RGG/\,
                  I1 =>  \52148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL05\     
  \=52152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52152\,
                  I0 =>  \52157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL05\    
  \=52153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52153\,
                  I0 =>  \52157\,
                  I1 =>  \52157\,
                  I2 =>  \52157\,
                  I3 =>  '0' );

  -- Alias \WL05/\    
  \=52154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52154\,
                  I0 =>  \52152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL05/\    
  \=52157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52157\,
                  I0 =>  \52141\,
                  I1 =>  \52142\,
                  I2 =>  \52151\,
                  I3 => \&52123\ );

  -- Alias \52157\    
  \=52158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52158\,
                  I0 =>  \MDT05\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&34452\ );

  -- Alias \CLROPE\   
  \=52162\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52162\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 => \&42152\ );

  -- Alias \G07/\     
  \=52163\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52163\,
                  I0 =>  \G07ED\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52447\ );

  -- Alias \CO08\     
  \=52201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52201\,
                  I0 =>  \XUY08/\,
                  I1 =>  \52210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52202\,
                  I0 =>  \A2XG/\,
                  I1 =>  \52220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52203\,
                   R => '0',
                   S => SYSRESET );

  \=52203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52203\,
                  I0 =>  \MONEX\,
                  I1 =>  \52202\,
                  I2 =>  \52204\,
                  I3 =>  '0' );

  \=52204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52204\,
                  I0 =>  \52203\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=52205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52205\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52206\,
                  I0 =>  \WL05/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52207\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52207\,
                   R => '0',
                   S => SYSRESET );

  \=52207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52207\,
                  I0 =>  \52205\,
                  I1 =>  \52206\,
                  I2 =>  \52208\,
                  I3 =>  '0' );

  \=52208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52208\,
                  I0 =>  \52207\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52209\,
                  I0 =>  \52203\,
                  I1 =>  \52207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY06/\   
  \=52210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52210\,
                  I0 =>  \52204\,
                  I1 =>  \52208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52211\,
                  I0 =>  \CI06/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA06/\  
  \=52212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52212\,
                  I0 =>  \52209\,
                  I1 =>  \52210\,
                  I2 =>  \CI06/\,
                  I3 =>  '0' );

  \=52213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52213\,
                  I0 =>  \52209\,
                  I1 =>  \52210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI07/\    
  \=52214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52214\,
                  I0 =>  \52209\,
                  I1 =>  \52212\,
                  I2 =>  \CO06\,
                  I3 =>  '0' );

  -- Alias \SUMB06/\  
  \=52215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52215\,
                  I0 =>  \52213\,
                  I1 =>  \52211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52217\,
                  I0 =>  \52212\,
                  I1 =>  \52215\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=52218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52218\,
                  I0 =>  \WAG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52219\,
                  I0 =>  \WL08/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A06/\     
  \:52220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52220\,
                   R => '0',
                   S => SYSRESET );

  \=52220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52220\,
                  I0 =>  \52218\,
                  I1 =>  \52219\,
                  I2 =>  \52221\,
                  I3 =>  '0' );

  \=52221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52221\,
                  I0 =>  \52220\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52222\,
                  I0 =>  \RAG/\,
                  I1 =>  \52220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52257\    
  \=52223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52223\,
                  I0 =>  \52217\,
                  I1 =>  \52222\,
                  I2 =>  \CH06\,
                  I3 => \&52233\ );

  \=52224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52224\,
                  I0 =>  \WLG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52225\,
                  I0 =>  \G09/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L06/\     
  \:52226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52226\,
                   R => '0',
                   S => SYSRESET );

  \=52226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52226\,
                  I0 =>  \52224\,
                  I1 =>  \52225\,
                  I2 =>  \52227\,
                  I3 =>  '0' );

  \=52227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52227\,
                  I0 =>  \52226\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52228\,
                  I0 =>  \RLG/\,
                  I1 =>  \52226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52229\,
                  I0 =>  \WQG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52230\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52230\,
                   R => '0',
                   S => SYSRESET );

  \=52230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52230\,
                  I0 =>  \52229\,
                  I1 =>  \52231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52231\,
                  I0 =>  \52230\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52232\,
                  I0 =>  \RQG/\,
                  I1 =>  \52230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52257\    
  \=52233\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52233\,
                  I0 =>  \52228\,
                  I1 =>  \52232\,
                  I2 =>  \52237\,
                  I3 => \&52258\ );

  \=52234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52234\,
                  I0 =>  \WZG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z06/\     
  \:52235\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52235\,
                   R => '0',
                   S => SYSRESET );

  \=52235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52235\,
                  I0 =>  \52234\,
                  I1 =>  \52236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52236\,
                  I0 =>  \52235\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52237\,
                  I0 =>  \RZG/\,
                  I1 =>  \52235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52238\,
                  I0 =>  \WBG/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52239\,
                   R => '0',
                   S => SYSRESET );

  \=52239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52239\,
                  I0 =>  \52238\,
                  I1 =>  \52240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52240\,
                  I0 =>  \52239\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52241\,
                  I0 =>  \RBLG/\,
                  I1 =>  \52239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52242\,
                  I0 =>  \52240\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52243\,
                  I0 =>  \WL05/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52244\,
                  I0 =>  \WL07/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52245\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52246\,
                  I0 =>  \WG1G/\,
                  I1 =>  \52254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52248\    
  \=52247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52247\,
                  I0 =>  \SA06\,
                  I1 =>  \52243\,
                  I2 =>  \52244\,
                  I3 =>  '0' );

  -- Alias \G06/\     
  \:52248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52248\,
                   R => '0',
                   S => SYSRESET );

  \=52248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52248\,
                  I0 =>  \52245\,
                  I1 =>  \52246\,
                  I2 =>  \52249\,
                  I3 => \&51363\ );

  -- Alias \G06\      
  \=52249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52249\,
                  I0 =>  \52248\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM06\    
  \=52250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52250\,
                  I0 =>  \52248\,
                  I1 =>  \52248\,
                  I2 =>  \52248\,
                  I3 =>  '0' );

  \=52251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52251\,
                  I0 =>  \RGG/\,
                  I1 =>  \52248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL06\     
  \=52252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52252\,
                  I0 =>  \52257\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL06\    
  \=52253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52253\,
                  I0 =>  \52257\,
                  I1 =>  \52257\,
                  I2 =>  \52257\,
                  I3 =>  '0' );

  -- Alias \WL06/\    
  \=52254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52254\,
                  I0 =>  \52252\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL06/\    
  \=52257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52257\,
                  I0 =>  \52241\,
                  I1 =>  \52242\,
                  I2 =>  \52251\,
                  I3 => \&52223\ );

  -- Alias \52257\    
  \=52258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52258\,
                  I0 =>  \MDT06\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&34453\ );

  -- Alias \PIPSAM/\  
  \=52261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52261\,
                  I0 =>  \PIPSAM\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A9 /2 - 4 BIT MODULE (2 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO10\     
  \=52301\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52301\,
                  I0 =>  \XUY10/\,
                  I1 =>  \52310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52302\,
                  I0 =>  \A2XG/\,
                  I1 =>  \52320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52303\,
                   R => '0',
                   S => SYSRESET );

  \=52303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52303\,
                  I0 =>  \MONEX\,
                  I1 =>  \52302\,
                  I2 =>  \52304\,
                  I3 =>  '0' );

  \=52304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52304\,
                  I0 =>  \52303\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=52305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52305\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52306\,
                  I0 =>  \WL07/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52307\,
                   R => '0',
                   S => SYSRESET );

  \=52307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52307\,
                  I0 =>  \52305\,
                  I1 =>  \52306\,
                  I2 =>  \52308\,
                  I3 =>  '0' );

  \=52308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52308\,
                  I0 =>  \52307\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52309\,
                  I0 =>  \52303\,
                  I1 =>  \52307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY08/\   
  \=52310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52310\,
                  I0 =>  \52304\,
                  I1 =>  \52308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52311\,
                  I0 =>  \CI08/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA08/\  
  \=52312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52312\,
                  I0 =>  \52309\,
                  I1 =>  \52310\,
                  I2 =>  \CI08/\,
                  I3 =>  '0' );

  \=52313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52313\,
                  I0 =>  \52309\,
                  I1 =>  \52310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI09/\    
  \=52314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52314\,
                  I0 =>  \52309\,
                  I1 =>  \52312\,
                  I2 =>  \CO08\,
                  I3 =>  '0' );

  -- Alias \SUMB08/\  
  \=52315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52315\,
                  I0 =>  \52313\,
                  I1 =>  \52311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52317\,
                  I0 =>  \52312\,
                  I1 =>  \52315\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=52318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52318\,
                  I0 =>  \WAG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52319\,
                  I0 =>  \WL10/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A08/\     
  \:52320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52320\,
                   R => '0',
                   S => SYSRESET );

  \=52320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52320\,
                  I0 =>  \52318\,
                  I1 =>  \52319\,
                  I2 =>  \52321\,
                  I3 =>  '0' );

  \=52321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52321\,
                  I0 =>  \52320\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52322\,
                  I0 =>  \RAG/\,
                  I1 =>  \52320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52357\    
  \=52323\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52323\,
                  I0 =>  \52317\,
                  I1 =>  \52322\,
                  I2 =>  \CH08\,
                  I3 => \&52333\ );

  \=52324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52324\,
                  I0 =>  \WLG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52325\,
                  I0 =>  \G11/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L08/\     
  \:52326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52326\,
                   R => '0',
                   S => SYSRESET );

  \=52326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52326\,
                  I0 =>  \52324\,
                  I1 =>  \52325\,
                  I2 =>  \52327\,
                  I3 =>  '0' );

  \=52327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52327\,
                  I0 =>  \52326\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52328\,
                  I0 =>  \RLG/\,
                  I1 =>  \52326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52329\,
                  I0 =>  \WQG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52330\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52330\,
                   R => '0',
                   S => SYSRESET );

  \=52330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52330\,
                  I0 =>  \52329\,
                  I1 =>  \52331\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52331\,
                  I0 =>  \52330\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52332\,
                  I0 =>  \RQG/\,
                  I1 =>  \52330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52357\    
  \=52333\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52333\,
                  I0 =>  \52328\,
                  I1 =>  \52332\,
                  I2 =>  \52337\,
                  I3 => \&52358\ );

  \=52334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52334\,
                  I0 =>  \WZG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z08/\     
  \:52335\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52335\,
                   R => '0',
                   S => SYSRESET );

  \=52335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52335\,
                  I0 =>  \52334\,
                  I1 =>  \52336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52336\,
                  I0 =>  \52335\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52337\,
                  I0 =>  \RZG/\,
                  I1 =>  \52335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52338\,
                  I0 =>  \WBG/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52339\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52339\,
                   R => '0',
                   S => SYSRESET );

  \=52339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52339\,
                  I0 =>  \52338\,
                  I1 =>  \52340\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52340\,
                  I0 =>  \52339\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52341\,
                  I0 =>  \RBLG/\,
                  I1 =>  \52339\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52342\,
                  I0 =>  \52340\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52343\,
                  I0 =>  \WL07/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52344\,
                  I0 =>  \WL09/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52345\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52346\,
                  I0 =>  \WG1G/\,
                  I1 =>  \52354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52348\    
  \=52347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52347\,
                  I0 =>  \SA08\,
                  I1 =>  \52343\,
                  I2 =>  \52344\,
                  I3 =>  '0' );

  -- Alias \G08/\     
  \:52348\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52348\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52348\,
                   R => '0',
                   S => SYSRESET );

  \=52348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52348\,
                  I0 =>  \52345\,
                  I1 =>  \52346\,
                  I2 =>  \52349\,
                  I3 => \&52347\ );

  -- Alias \G08\      
  \=52349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52349\,
                  I0 =>  \52348\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM08\    
  \=52350\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52350\,
                  I0 =>  \52348\,
                  I1 =>  \52348\,
                  I2 =>  \52348\,
                  I3 =>  '0' );

  \=52351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52351\,
                  I0 =>  \RGG/\,
                  I1 =>  \52348\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL08\     
  \=52352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52352\,
                  I0 =>  \52357\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL08\    
  \=52353\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52353\,
                  I0 =>  \52357\,
                  I1 =>  \52357\,
                  I2 =>  \52357\,
                  I3 =>  '0' );

  -- Alias \WL08/\    
  \=52354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52354\,
                  I0 =>  \52352\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL08/\    
  \=52357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52357\,
                  I0 =>  \52341\,
                  I1 =>  \52342\,
                  I2 =>  \52351\,
                  I3 => \&52323\ );

  -- Alias \52357\    
  \=52358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52358\,
                  I0 =>  \MDT08\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPGX-\   
  \=52361\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52361\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAX-/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPGY+\   
  \=52362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52362\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAY+/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ROPET\    
  \=52363\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52363\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 => \&35458\ );

  -- Alias \CO10\     
  \=52401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52401\,
                  I0 =>  \XUY09/\,
                  I1 =>  \52410\,
                  I2 =>  \CI07/\,
                  I3 => \&52301\ );

  \=52402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52402\,
                  I0 =>  \A2XG/\,
                  I1 =>  \52420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52403\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52403\,
                   R => '0',
                   S => SYSRESET );

  \=52403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52403\,
                  I0 =>  \MONEX\,
                  I1 =>  \52402\,
                  I2 =>  \52404\,
                  I3 =>  '0' );

  \=52404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52404\,
                  I0 =>  \52403\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=52405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52405\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52406\,
                  I0 =>  \WL06/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52407\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52407\,
                   R => '0',
                   S => SYSRESET );

  \=52407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52407\,
                  I0 =>  \52405\,
                  I1 =>  \52406\,
                  I2 =>  \52408\,
                  I3 =>  '0' );

  \=52408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52408\,
                  I0 =>  \52407\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52409\,
                  I0 =>  \52403\,
                  I1 =>  \52407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY07/\   
  \=52410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52410\,
                  I0 =>  \52404\,
                  I1 =>  \52408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52411\,
                  I0 =>  \CI07/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA07/\  
  \=52412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52412\,
                  I0 =>  \52409\,
                  I1 =>  \CI07/\,
                  I2 =>  \52410\,
                  I3 => \&54462\ );

  \=52413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52413\,
                  I0 =>  \52409\,
                  I1 =>  \52410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI08/\    
  \=52414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52414\,
                  I0 =>  \52409\,
                  I1 =>  \52412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB07/\  
  \=52415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52415\,
                  I0 =>  \52413\,
                  I1 =>  \52411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52417\,
                  I0 =>  \52412\,
                  I1 =>  \52415\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=52418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52418\,
                  I0 =>  \WAG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52419\,
                  I0 =>  \WL09/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A07/\     
  \:52420\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52420\,
                   R => '0',
                   S => SYSRESET );

  \=52420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52420\,
                  I0 =>  \52418\,
                  I1 =>  \52419\,
                  I2 =>  \52421\,
                  I3 =>  '0' );

  \=52421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52421\,
                  I0 =>  \52420\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52422\,
                  I0 =>  \RAG/\,
                  I1 =>  \52420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52457\    
  \=52423\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52423\,
                  I0 =>  \52417\,
                  I1 =>  \52422\,
                  I2 =>  \CH07\,
                  I3 => \&52433\ );

  \=52424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52424\,
                  I0 =>  \WLG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52425\,
                  I0 =>  \G10/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L07/\     
  \:52426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52426\,
                   R => '0',
                   S => SYSRESET );

  \=52426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52426\,
                  I0 =>  \52424\,
                  I1 =>  \52425\,
                  I2 =>  \52427\,
                  I3 =>  '0' );

  \=52427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52427\,
                  I0 =>  \52426\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52428\,
                  I0 =>  \RLG/\,
                  I1 =>  \52426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52429\,
                  I0 =>  \WQG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52430\,
                   R => '0',
                   S => SYSRESET );

  \=52430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52430\,
                  I0 =>  \52429\,
                  I1 =>  \52431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52431\,
                  I0 =>  \52430\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52432\,
                  I0 =>  \RQG/\,
                  I1 =>  \52430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52457\    
  \=52433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52433\,
                  I0 =>  \52428\,
                  I1 =>  \52432\,
                  I2 =>  \52437\,
                  I3 => \&52458\ );

  \=52434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52434\,
                  I0 =>  \WZG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z07/\     
  \:52435\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52435\,
                   R => '0',
                   S => SYSRESET );

  \=52435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52435\,
                  I0 =>  \52434\,
                  I1 =>  \52436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52436\,
                  I0 =>  \52435\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52437\,
                  I0 =>  \RZG/\,
                  I1 =>  \52435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52438\,
                  I0 =>  \WBG/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:52439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52439\,
                   R => '0',
                   S => SYSRESET );

  \=52439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52439\,
                  I0 =>  \52438\,
                  I1 =>  \52440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52440\,
                  I0 =>  \52439\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52441\,
                  I0 =>  \RBLG/\,
                  I1 =>  \52439\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52442\,
                  I0 =>  \52440\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52443\,
                  I0 =>  \WL06/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52444\,
                  I0 =>  \WL08/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52445\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=52446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52446\,
                  I0 =>  \WG1G/\,
                  I1 =>  \52454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \52448\    
  \=52447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52447\,
                  I0 =>  \SA07\,
                  I1 =>  \52443\,
                  I2 =>  \52444\,
                  I3 =>  '0' );

  -- Alias \G07/\     
  \:52448\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \52448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$52448\,
                   R => '0',
                   S => SYSRESET );

  \=52448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$52448\,
                  I0 =>  \52445\,
                  I1 =>  \52446\,
                  I2 =>  \52449\,
                  I3 => \&52163\ );

  -- Alias \G07\      
  \=52449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52449\,
                  I0 =>  \52448\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM07\    
  \=52450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52450\,
                  I0 =>  \52448\,
                  I1 =>  \52448\,
                  I2 =>  \52448\,
                  I3 =>  '0' );

  \=52451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52451\,
                  I0 =>  \RGG/\,
                  I1 =>  \52448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL07\     
  \=52452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52452\,
                  I0 =>  \52457\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL07\    
  \=52453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52453\,
                  I0 =>  \52457\,
                  I1 =>  \52457\,
                  I2 =>  \52457\,
                  I3 =>  '0' );

  -- Alias \WL07/\    
  \=52454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52454\,
                  I0 =>  \52452\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL07/\    
  \=52457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52457\,
                  I0 =>  \52441\,
                  I1 =>  \52442\,
                  I2 =>  \52451\,
                  I3 => \&52423\ );

  -- Alias \52457\    
  \=52458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52458\,
                  I0 =>  \MDT07\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPGX+\   
  \=52461\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \52461\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAX+/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ROPER\    
  \=52462\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52462\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 => \&35422\ );

  -- Alias \ROPES\    
  \=52463\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&52463\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 => \&35441\ );

  -- ****************************************
  -- ***                                  ***
  -- ***  A10/1 - 4 BIT MODULE (3 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO12\     
  \=53101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53101\,
                  I0 =>  \XUY11/\,
                  I1 =>  \53110\,
                  I2 =>  \CI09/\,
                  I3 => \&53201\ );

  \=53102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53102\,
                  I0 =>  \A2XG/\,
                  I1 =>  \53120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53103\,
                   R => '0',
                   S => SYSRESET );

  \=53103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53103\,
                  I0 =>  \MONEX\,
                  I1 =>  \53102\,
                  I2 =>  \53104\,
                  I3 =>  '0' );

  \=53104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53104\,
                  I0 =>  \53103\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=53105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53105\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53106\,
                  I0 =>  \WL08/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53107\,
                   R => '0',
                   S => SYSRESET );

  \=53107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53107\,
                  I0 =>  \53105\,
                  I1 =>  \53106\,
                  I2 =>  \53108\,
                  I3 =>  '0' );

  \=53108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53108\,
                  I0 =>  \53107\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53109\,
                  I0 =>  \53103\,
                  I1 =>  \53107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY09/\   
  \=53110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53110\,
                  I0 =>  \53104\,
                  I1 =>  \53108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53111\,
                  I0 =>  \CI09/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA09/\  
  \=53112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53112\,
                  I0 =>  \53109\,
                  I1 =>  \CI09/\,
                  I2 =>  \53110\,
                  I3 =>  '0' );

  \=53113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53113\,
                  I0 =>  \53109\,
                  I1 =>  \53110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI10/\    
  \=53114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53114\,
                  I0 =>  \53109\,
                  I1 =>  \53112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB09/\  
  \=53115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53115\,
                  I0 =>  \53113\,
                  I1 =>  \53111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53117\,
                  I0 =>  \53112\,
                  I1 =>  \53115\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=53118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53118\,
                  I0 =>  \WAG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53119\,
                  I0 =>  \WL11/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A09/\     
  \:53120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53120\,
                   R => '0',
                   S => SYSRESET );

  \=53120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53120\,
                  I0 =>  \53118\,
                  I1 =>  \53119\,
                  I2 =>  \53121\,
                  I3 =>  '0' );

  \=53121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53121\,
                  I0 =>  \53120\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53122\,
                  I0 =>  \RAG/\,
                  I1 =>  \53120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53157\    
  \=53123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53123\,
                  I0 =>  \53117\,
                  I1 =>  \53122\,
                  I2 =>  \CH09\,
                  I3 => \&53133\ );

  \=53124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53124\,
                  I0 =>  \WLG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53125\,
                  I0 =>  \G12/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L09/\     
  \:53126\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53126\,
                   R => '0',
                   S => SYSRESET );

  \=53126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53126\,
                  I0 =>  \53124\,
                  I1 =>  \53125\,
                  I2 =>  \53127\,
                  I3 =>  '0' );

  \=53127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53127\,
                  I0 =>  \53126\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53128\,
                  I0 =>  \RLG/\,
                  I1 =>  \53126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53129\,
                  I0 =>  \WQG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53130\,
                   R => '0',
                   S => SYSRESET );

  \=53130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53130\,
                  I0 =>  \53129\,
                  I1 =>  \53131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53131\,
                  I0 =>  \53130\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53132\,
                  I0 =>  \RQG/\,
                  I1 =>  \53130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53157\    
  \=53133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53133\,
                  I0 =>  \53128\,
                  I1 =>  \53132\,
                  I2 =>  \53137\,
                  I3 => \&53158\ );

  \=53134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53134\,
                  I0 =>  \WZG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z09/\     
  \:53135\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53135\,
                   R => '0',
                   S => SYSRESET );

  \=53135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53135\,
                  I0 =>  \53134\,
                  I1 =>  \53136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53136\,
                  I0 =>  \53135\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53137\,
                  I0 =>  \RZG/\,
                  I1 =>  \53135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53138\,
                  I0 =>  \WBG/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53139\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53139\,
                   R => '0',
                   S => SYSRESET );

  \=53139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53139\,
                  I0 =>  \53138\,
                  I1 =>  \53140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53140\,
                  I0 =>  \53139\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53141\,
                  I0 =>  \RBLG/\,
                  I1 =>  \53139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53142\,
                  I0 =>  \53140\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53143\,
                  I0 =>  \WL08/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53144\,
                  I0 =>  \WL10/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53145\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53146\,
                  I0 =>  \WG1G/\,
                  I1 =>  \53154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53148\    
  \=53147\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53147\,
                  I0 =>  \SA09\,
                  I1 =>  \53143\,
                  I2 =>  \53144\,
                  I3 =>  '0' );

  -- Alias \G09/\     
  \:53148\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53148\,
                   R => '0',
                   S => SYSRESET );

  \=53148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53148\,
                  I0 =>  \53145\,
                  I1 =>  \53146\,
                  I2 =>  \53149\,
                  I3 => \&53147\ );

  -- Alias \G09\      
  \=53149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53149\,
                  I0 =>  \53148\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM09\    
  \=53150\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53150\,
                  I0 =>  \53148\,
                  I1 =>  \53148\,
                  I2 =>  \53148\,
                  I3 =>  '0' );

  \=53151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53151\,
                  I0 =>  \RGG/\,
                  I1 =>  \53148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL09\     
  \=53152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53152\,
                  I0 =>  \53157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL09\    
  \=53153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53153\,
                  I0 =>  \53157\,
                  I1 =>  \53157\,
                  I2 =>  \53157\,
                  I3 =>  '0' );

  -- Alias \WL09/\    
  \=53154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53154\,
                  I0 =>  \53152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL09/\    
  \=53157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53157\,
                  I0 =>  \53141\,
                  I1 =>  \53142\,
                  I2 =>  \53151\,
                  I3 => \&53123\ );

  -- Alias \53157\    
  \=53158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53158\,
                  I0 =>  \MDT09\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35149\ );

  -- Alias \PIPGY-\   
  \=53161\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53161\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAY-/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CO12\     
  \=53201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53201\,
                  I0 =>  \XUY12/\,
                  I1 =>  \53210\,
                  I2 =>  '0',
                  I3 => \&53463\ );

  \=53202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53202\,
                  I0 =>  \A2XG/\,
                  I1 =>  \53220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53203\,
                   R => '0',
                   S => SYSRESET );

  \=53203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53203\,
                  I0 =>  \MONEX\,
                  I1 =>  \53202\,
                  I2 =>  \53204\,
                  I3 =>  '0' );

  \=53204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53204\,
                  I0 =>  \53203\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=53205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53205\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53206\,
                  I0 =>  \WL09/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53207\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53207\,
                   R => '0',
                   S => SYSRESET );

  \=53207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53207\,
                  I0 =>  \53205\,
                  I1 =>  \53206\,
                  I2 =>  \53208\,
                  I3 =>  '0' );

  \=53208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53208\,
                  I0 =>  \53207\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53209\,
                  I0 =>  \53203\,
                  I1 =>  \53207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY10/\   
  \=53210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53210\,
                  I0 =>  \53204\,
                  I1 =>  \53208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53211\,
                  I0 =>  \CI10/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA10/\  
  \=53212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53212\,
                  I0 =>  \53209\,
                  I1 =>  \53210\,
                  I2 =>  \CI10/\,
                  I3 =>  '0' );

  \=53213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53213\,
                  I0 =>  \53209\,
                  I1 =>  \53210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI11/\    
  \=53214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53214\,
                  I0 =>  \53209\,
                  I1 =>  \53212\,
                  I2 =>  \CO10\,
                  I3 =>  '0' );

  -- Alias \SUMB10/\  
  \=53215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53215\,
                  I0 =>  \53213\,
                  I1 =>  \53211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53217\,
                  I0 =>  \53212\,
                  I1 =>  \53215\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=53218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53218\,
                  I0 =>  \WAG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53219\,
                  I0 =>  \WL12/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A10/\     
  \:53220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53220\,
                   R => '0',
                   S => SYSRESET );

  \=53220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53220\,
                  I0 =>  \53218\,
                  I1 =>  \53219\,
                  I2 =>  \53221\,
                  I3 =>  '0' );

  \=53221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53221\,
                  I0 =>  \53220\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53222\,
                  I0 =>  \RAG/\,
                  I1 =>  \53220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53257\    
  \=53223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53223\,
                  I0 =>  \53217\,
                  I1 =>  \53222\,
                  I2 =>  \CH10\,
                  I3 => \&53233\ );

  \=53224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53224\,
                  I0 =>  \WLG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53225\,
                  I0 =>  \G13/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L10/\     
  \:53226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53226\,
                   R => '0',
                   S => SYSRESET );

  \=53226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53226\,
                  I0 =>  \53224\,
                  I1 =>  \53225\,
                  I2 =>  \53227\,
                  I3 =>  '0' );

  \=53227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53227\,
                  I0 =>  \53226\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53228\,
                  I0 =>  \RLG/\,
                  I1 =>  \53226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53229\,
                  I0 =>  \WQG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53230\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53230\,
                   R => '0',
                   S => SYSRESET );

  \=53230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53230\,
                  I0 =>  \53229\,
                  I1 =>  \53231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53231\,
                  I0 =>  \53230\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53232\,
                  I0 =>  \RQG/\,
                  I1 =>  \53230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53257\    
  \=53233\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53233\,
                  I0 =>  \53228\,
                  I1 =>  \53232\,
                  I2 =>  \53237\,
                  I3 => \&53258\ );

  \=53234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53234\,
                  I0 =>  \WZG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z10/\     
  \:53235\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53235\,
                   R => '0',
                   S => SYSRESET );

  \=53235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53235\,
                  I0 =>  \53234\,
                  I1 =>  \53236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53236\,
                  I0 =>  \53235\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53237\,
                  I0 =>  \RZG/\,
                  I1 =>  \53235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53238\,
                  I0 =>  \WBG/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53239\,
                   R => '0',
                   S => SYSRESET );

  \=53239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53239\,
                  I0 =>  \53238\,
                  I1 =>  \53240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53240\,
                  I0 =>  \53239\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53241\,
                  I0 =>  \RBLG/\,
                  I1 =>  \53239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53242\,
                  I0 =>  \53240\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53243\,
                  I0 =>  \WL09/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53244\,
                  I0 =>  \WL11/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53245\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53246\,
                  I0 =>  \WG1G/\,
                  I1 =>  \53254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53248\    
  \=53247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53247\,
                  I0 =>  \SA10\,
                  I1 =>  \53243\,
                  I2 =>  \53244\,
                  I3 =>  '0' );

  -- Alias \G10/\     
  \:53248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53248\,
                   R => '0',
                   S => SYSRESET );

  \=53248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53248\,
                  I0 =>  \53245\,
                  I1 =>  \53246\,
                  I2 =>  \53249\,
                  I3 => \&53247\ );

  -- Alias \G10\      
  \=53249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53249\,
                  I0 =>  \53248\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM10\    
  \=53250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53250\,
                  I0 =>  \53248\,
                  I1 =>  \53248\,
                  I2 =>  \53248\,
                  I3 =>  '0' );

  \=53251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53251\,
                  I0 =>  \RGG/\,
                  I1 =>  \53248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL10\     
  \=53252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53252\,
                  I0 =>  \53257\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL10\    
  \=53253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53253\,
                  I0 =>  \53257\,
                  I1 =>  \53257\,
                  I2 =>  \53257\,
                  I3 =>  '0' );

  -- Alias \WL10/\    
  \=53254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53254\,
                  I0 =>  \53252\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL10/\    
  \=53257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53257\,
                  I0 =>  \53241\,
                  I1 =>  \53242\,
                  I2 =>  \53251\,
                  I3 => \&53223\ );

  -- Alias \53257\    
  \=53258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53258\,
                  I0 =>  \MDT10\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35141\ );

  -- Alias \PIPGZ+\   
  \=53261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53261\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAZ+/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPGZ-\   
  \=53262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53262\,
                  I0 =>  \PIPSAM/\,
                  I1 =>  \PIPAZ-/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A10/2 - 4 BIT MODULE (3 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO14\     
  \=53301\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53301\,
                  I0 =>  \XUY14/\,
                  I1 =>  \53310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53302\,
                  I0 =>  \A2XG/\,
                  I1 =>  \53320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53303\,
                   R => '0',
                   S => SYSRESET );

  \=53303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53303\,
                  I0 =>  \MONEX\,
                  I1 =>  \53302\,
                  I2 =>  \53304\,
                  I3 =>  '0' );

  \=53304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53304\,
                  I0 =>  \53303\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=53305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53305\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53306\,
                  I0 =>  \WL11/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53307\,
                   R => '0',
                   S => SYSRESET );

  \=53307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53307\,
                  I0 =>  \53305\,
                  I1 =>  \53306\,
                  I2 =>  \53308\,
                  I3 =>  '0' );

  \=53308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53308\,
                  I0 =>  \53307\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53309\,
                  I0 =>  \53303\,
                  I1 =>  \53307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY12/\   
  \=53310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53310\,
                  I0 =>  \53304\,
                  I1 =>  \53308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53311\,
                  I0 =>  \CI12/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA12/\  
  \=53312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53312\,
                  I0 =>  \53309\,
                  I1 =>  \53310\,
                  I2 =>  \CI12/\,
                  I3 => \&54463\ );

  \=53313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53313\,
                  I0 =>  \53309\,
                  I1 =>  \53310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI13/\    
  \=53314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53314\,
                  I0 =>  \53309\,
                  I1 =>  \53312\,
                  I2 =>  \CO12\,
                  I3 =>  '0' );

  -- Alias \SUMB12/\  
  \=53315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53315\,
                  I0 =>  \53313\,
                  I1 =>  \53311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53317\,
                  I0 =>  \53312\,
                  I1 =>  \53315\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=53318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53318\,
                  I0 =>  \WAG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53319\,
                  I0 =>  \WL14/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A12/\     
  \:53320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53320\,
                   R => '0',
                   S => SYSRESET );

  \=53320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53320\,
                  I0 =>  \53318\,
                  I1 =>  \53319\,
                  I2 =>  \53321\,
                  I3 =>  '0' );

  \=53321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53321\,
                  I0 =>  \53320\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53322\,
                  I0 =>  \RAG/\,
                  I1 =>  \53320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53357\    
  \=53323\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53323\,
                  I0 =>  \53317\,
                  I1 =>  \53322\,
                  I2 =>  \CH12\,
                  I3 => \&53333\ );

  \=53324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53324\,
                  I0 =>  \WLG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53325\,
                  I0 =>  \G15/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L12/\     
  \:53326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53326\,
                   R => '0',
                   S => SYSRESET );

  \=53326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53326\,
                  I0 =>  \53324\,
                  I1 =>  \53325\,
                  I2 =>  \53327\,
                  I3 =>  '0' );

  \=53327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53327\,
                  I0 =>  \53326\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53328\,
                  I0 =>  \RLG/\,
                  I1 =>  \53326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53329\,
                  I0 =>  \WQG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53330\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53330\,
                   R => '0',
                   S => SYSRESET );

  \=53330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53330\,
                  I0 =>  \53329\,
                  I1 =>  \53331\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53331\,
                  I0 =>  \53330\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53332\,
                  I0 =>  \RQG/\,
                  I1 =>  \53330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53357\    
  \=53333\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53333\,
                  I0 =>  \53328\,
                  I1 =>  \53332\,
                  I2 =>  \53337\,
                  I3 => \&53358\ );

  \=53334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53334\,
                  I0 =>  \WZG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z12/\     
  \:53335\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53335\,
                   R => '0',
                   S => SYSRESET );

  \=53335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53335\,
                  I0 =>  \53334\,
                  I1 =>  \53336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53336\,
                  I0 =>  \53335\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53337\,
                  I0 =>  \RZG/\,
                  I1 =>  \53335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53338\,
                  I0 =>  \WBG/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53339\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53339\,
                   R => '0',
                   S => SYSRESET );

  \=53339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53339\,
                  I0 =>  \53338\,
                  I1 =>  \53340\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53340\,
                  I0 =>  \53339\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53341\,
                  I0 =>  \RBHG/\,
                  I1 =>  \53339\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53342\,
                  I0 =>  \53340\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53343\,
                  I0 =>  \WL11/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53344\,
                  I0 =>  \WL13/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53345\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53346\,
                  I0 =>  \WG1G/\,
                  I1 =>  \53354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53348\    
  \=53347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53347\,
                  I0 =>  \SA12\,
                  I1 =>  \53343\,
                  I2 =>  \53344\,
                  I3 =>  '0' );

  -- Alias \G12/\     
  \:53348\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53348\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53348\,
                   R => '0',
                   S => SYSRESET );

  \=53348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53348\,
                  I0 =>  \53345\,
                  I1 =>  \53346\,
                  I2 =>  \53349\,
                  I3 => \&53347\ );

  -- Alias \G12\      
  \=53349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53349\,
                  I0 =>  \53348\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM12\    
  \=53350\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53350\,
                  I0 =>  \53348\,
                  I1 =>  \53348\,
                  I2 =>  \53348\,
                  I3 =>  '0' );

  \=53351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53351\,
                  I0 =>  \RGG/\,
                  I1 =>  \53348\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL12\     
  \=53352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53352\,
                  I0 =>  \53357\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL12\    
  \=53353\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53353\,
                  I0 =>  \53357\,
                  I1 =>  \53357\,
                  I2 =>  \53357\,
                  I3 =>  '0' );

  -- Alias \WL12/\    
  \=53354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53354\,
                  I0 =>  \53352\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL12/\    
  \=53357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53357\,
                  I0 =>  \53341\,
                  I1 =>  \53342\,
                  I2 =>  \53351\,
                  I3 => \&53323\ );

  -- Alias \53357\    
  \=53358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53358\,
                  I0 =>  \MDT12\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35122\ );

  -- Alias \PIPAX-/\  
  \=53361\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53361\,
                  I0 =>  \PIPAX-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPAY+/\  
  \=53362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53362\,
                  I0 =>  \PIPAY+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL15/\    
  \=53363\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53363\,
                  I0 =>  \BK16\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54423\ );

  -- Alias \CO14\     
  \=53401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53401\,
                  I0 =>  \XUY13/\,
                  I1 =>  \53410\,
                  I2 =>  \CI11/\,
                  I3 => \&53301\ );

  \=53402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53402\,
                  I0 =>  \A2XG/\,
                  I1 =>  \53420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53403\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53403\,
                   R => '0',
                   S => SYSRESET );

  \=53403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53403\,
                  I0 =>  \MONEX\,
                  I1 =>  \53402\,
                  I2 =>  \53404\,
                  I3 =>  '0' );

  \=53404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53404\,
                  I0 =>  \53403\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=53405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53405\,
                  I0 =>  \WYLOG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53406\,
                  I0 =>  \WL10/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53407\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53407\,
                   R => '0',
                   S => SYSRESET );

  \=53407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53407\,
                  I0 =>  \53405\,
                  I1 =>  \53406\,
                  I2 =>  \53408\,
                  I3 =>  '0' );

  \=53408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53408\,
                  I0 =>  \53407\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53409\,
                  I0 =>  \53403\,
                  I1 =>  \53407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY11/\   
  \=53410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53410\,
                  I0 =>  \53404\,
                  I1 =>  \53408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53411\,
                  I0 =>  \CI11/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA11/\  
  \=53412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53412\,
                  I0 =>  \53409\,
                  I1 =>  \CI11/\,
                  I2 =>  \53410\,
                  I3 =>  '0' );

  \=53413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53413\,
                  I0 =>  \53409\,
                  I1 =>  \53410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI12/\    
  \=53414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53414\,
                  I0 =>  \53409\,
                  I1 =>  \53412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB11/\  
  \=53415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53415\,
                  I0 =>  \53413\,
                  I1 =>  \53411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53417\,
                  I0 =>  \53412\,
                  I1 =>  \53415\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=53418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53418\,
                  I0 =>  \WAG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53419\,
                  I0 =>  \WL13/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A11/\     
  \:53420\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53420\,
                   R => '0',
                   S => SYSRESET );

  \=53420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53420\,
                  I0 =>  \53418\,
                  I1 =>  \53419\,
                  I2 =>  \53421\,
                  I3 =>  '0' );

  \=53421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53421\,
                  I0 =>  \53420\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53422\,
                  I0 =>  \RAG/\,
                  I1 =>  \53420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53457\    
  \=53423\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53423\,
                  I0 =>  \53417\,
                  I1 =>  \53422\,
                  I2 =>  \CH11\,
                  I3 => \&53433\ );

  \=53424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53424\,
                  I0 =>  \WLG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53425\,
                  I0 =>  \G14/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L11/\     
  \:53426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53426\,
                   R => '0',
                   S => SYSRESET );

  \=53426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53426\,
                  I0 =>  \53424\,
                  I1 =>  \53425\,
                  I2 =>  \53427\,
                  I3 =>  '0' );

  \=53427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53427\,
                  I0 =>  \53426\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53428\,
                  I0 =>  \RLG/\,
                  I1 =>  \53426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53429\,
                  I0 =>  \WQG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53430\,
                   R => '0',
                   S => SYSRESET );

  \=53430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53430\,
                  I0 =>  \53429\,
                  I1 =>  \53431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53431\,
                  I0 =>  \53430\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53432\,
                  I0 =>  \RQG/\,
                  I1 =>  \53430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53457\    
  \=53433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53433\,
                  I0 =>  \53428\,
                  I1 =>  \53432\,
                  I2 =>  \53437\,
                  I3 => \&53458\ );

  \=53434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53434\,
                  I0 =>  \WZG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z11/\     
  \:53435\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53435\,
                   R => '0',
                   S => SYSRESET );

  \=53435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53435\,
                  I0 =>  \53434\,
                  I1 =>  \53436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53436\,
                  I0 =>  \53435\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53437\,
                  I0 =>  \RZG/\,
                  I1 =>  \53435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53438\,
                  I0 =>  \WBG/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:53439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53439\,
                   R => '0',
                   S => SYSRESET );

  \=53439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53439\,
                  I0 =>  \53438\,
                  I1 =>  \53440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53440\,
                  I0 =>  \53439\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53441\,
                  I0 =>  \RBHG/\,
                  I1 =>  \53439\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53442\,
                  I0 =>  \53440\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53443\,
                  I0 =>  \WL10/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53444\,
                  I0 =>  \WL12/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53445\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=53446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53446\,
                  I0 =>  \WG1G/\,
                  I1 =>  \53454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \53448\    
  \=53447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53447\,
                  I0 =>  \SA11\,
                  I1 =>  \53443\,
                  I2 =>  \53444\,
                  I3 =>  '0' );

  -- Alias \G11/\     
  \:53448\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \53448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$53448\,
                   R => '0',
                   S => SYSRESET );

  \=53448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$53448\,
                  I0 =>  \53445\,
                  I1 =>  \53446\,
                  I2 =>  \53449\,
                  I3 => \&53447\ );

  -- Alias \G11\      
  \=53449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53449\,
                  I0 =>  \53448\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM11\    
  \=53450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53450\,
                  I0 =>  \53448\,
                  I1 =>  \53448\,
                  I2 =>  \53448\,
                  I3 =>  '0' );

  \=53451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53451\,
                  I0 =>  \RGG/\,
                  I1 =>  \53448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL11\     
  \=53452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53452\,
                  I0 =>  \53457\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL11\    
  \=53453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53453\,
                  I0 =>  \53457\,
                  I1 =>  \53457\,
                  I2 =>  \53457\,
                  I3 =>  '0' );

  -- Alias \WL11/\    
  \=53454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53454\,
                  I0 =>  \53452\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL11/\    
  \=53457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53457\,
                  I0 =>  \53441\,
                  I1 =>  \53442\,
                  I2 =>  \53451\,
                  I3 => \&53423\ );

  -- Alias \53457\    
  \=53458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53458\,
                  I0 =>  \MDT11\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35127\ );

  -- Alias \PIPAX+/\  
  \=53461\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \53461\,
                  I0 =>  \PIPAX+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CO04\     
  \=53462\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53462\,
                  I0 =>  \WHOMPA\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CO12\     
  \=53463\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&53463\,
                  I0 =>  \WHOMPA\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A11/1 - 4 BIT MODULE (4 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO16\     
  \=54101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54101\,
                  I0 =>  \XUY15/\,
                  I1 =>  \54110\,
                  I2 =>  \CI13/\,
                  I3 => \&54201\ );

  \=54102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54102\,
                  I0 =>  \A2XG/\,
                  I1 =>  \54120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54103\,
                   R => '0',
                   S => SYSRESET );

  \=54103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54103\,
                  I0 =>  \MONEX\,
                  I1 =>  \54102\,
                  I2 =>  \54104\,
                  I3 =>  '0' );

  \=54104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54104\,
                  I0 =>  \54103\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=54105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54105\,
                  I0 =>  \WYHIG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54106\,
                  I0 =>  \WL12/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54107\,
                   R => '0',
                   S => SYSRESET );

  \=54107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54107\,
                  I0 =>  \54105\,
                  I1 =>  \54106\,
                  I2 =>  \54108\,
                  I3 =>  '0' );

  \=54108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54108\,
                  I0 =>  \54107\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54109\,
                  I0 =>  \54103\,
                  I1 =>  \54107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY13/\   
  \=54110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54110\,
                  I0 =>  \54104\,
                  I1 =>  \54108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54111\,
                  I0 =>  \CI13/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA13/\  
  \=54112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54112\,
                  I0 =>  \54109\,
                  I1 =>  \CI13/\,
                  I2 =>  \54110\,
                  I3 =>  '0' );

  \=54113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54113\,
                  I0 =>  \54109\,
                  I1 =>  \54110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI14/\    
  \=54114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54114\,
                  I0 =>  \54109\,
                  I1 =>  \54112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB13/\  
  \=54115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54115\,
                  I0 =>  \54113\,
                  I1 =>  \54111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54117\,
                  I0 =>  \54112\,
                  I1 =>  \54115\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=54118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54118\,
                  I0 =>  \WAG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54119\,
                  I0 =>  \WL15/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A13/\     
  \:54120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54120\,
                   R => '0',
                   S => SYSRESET );

  \=54120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54120\,
                  I0 =>  \54118\,
                  I1 =>  \54119\,
                  I2 =>  \54121\,
                  I3 =>  '0' );

  \=54121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54121\,
                  I0 =>  \54120\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54122\,
                  I0 =>  \RAG/\,
                  I1 =>  \54120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54157\    
  \=54123\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54123\,
                  I0 =>  \54117\,
                  I1 =>  \54122\,
                  I2 =>  \CH13\,
                  I3 => \&54133\ );

  \=54124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54124\,
                  I0 =>  \WLG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54125\,
                  I0 =>  \WL01/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L13/\     
  \:54126\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54126\,
                   R => '0',
                   S => SYSRESET );

  \=54126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54126\,
                  I0 =>  \54124\,
                  I1 =>  \54125\,
                  I2 =>  \54127\,
                  I3 =>  '0' );

  \=54127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54127\,
                  I0 =>  \54126\,
                  I1 =>  \CLG2G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54128\,
                  I0 =>  \RLG/\,
                  I1 =>  \54126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54129\,
                  I0 =>  \WQG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54130\,
                   R => '0',
                   S => SYSRESET );

  \=54130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54130\,
                  I0 =>  \54129\,
                  I1 =>  \54131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54131\,
                  I0 =>  \54130\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54132\,
                  I0 =>  \RQG/\,
                  I1 =>  \54130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54157\    
  \=54133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54133\,
                  I0 =>  \54128\,
                  I1 =>  \54132\,
                  I2 =>  \54137\,
                  I3 => \&54158\ );

  \=54134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54134\,
                  I0 =>  \WZG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z13/\     
  \:54135\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54135\,
                   R => '0',
                   S => SYSRESET );

  \=54135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54135\,
                  I0 =>  \54134\,
                  I1 =>  \54136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54136\,
                  I0 =>  \54135\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54137\,
                  I0 =>  \RZG/\,
                  I1 =>  \54135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54138\,
                  I0 =>  \WBG/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54139\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54139\,
                   R => '0',
                   S => SYSRESET );

  \=54139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54139\,
                  I0 =>  \54138\,
                  I1 =>  \54140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54140\,
                  I0 =>  \54139\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54141\,
                  I0 =>  \RBHG/\,
                  I1 =>  \54139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54142\,
                  I0 =>  \54140\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54143\,
                  I0 =>  \WL12/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54144\,
                  I0 =>  \WL14/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54145\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54146\,
                  I0 =>  \WG1G/\,
                  I1 =>  \54154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54148\    
  \=54147\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54147\,
                  I0 =>  \SA13\,
                  I1 =>  \54143\,
                  I2 =>  \54144\,
                  I3 =>  '0' );

  -- Alias \G13/\     
  \:54148\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54148\,
                   R => '0',
                   S => SYSRESET );

  \=54148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54148\,
                  I0 =>  \54145\,
                  I1 =>  \54146\,
                  I2 =>  \54149\,
                  I3 => \&54147\ );

  -- Alias \G13\      
  \=54149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54149\,
                  I0 =>  \54148\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM13\    
  \=54150\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54150\,
                  I0 =>  \54148\,
                  I1 =>  \54148\,
                  I2 =>  \54148\,
                  I3 =>  '0' );

  \=54151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54151\,
                  I0 =>  \RGG/\,
                  I1 =>  \54148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL13\     
  \=54152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54152\,
                  I0 =>  \54157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL13\    
  \=54153\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54153\,
                  I0 =>  \54157\,
                  I1 =>  \54157\,
                  I2 =>  \54157\,
                  I3 =>  '0' );

  -- Alias \WL13/\    
  \=54154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54154\,
                  I0 =>  \54152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL13/\    
  \=54157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54157\,
                  I0 =>  \54141\,
                  I1 =>  \54142\,
                  I2 =>  \54151\,
                  I3 => \&54123\ );

  -- Alias \54157\    
  \=54158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54158\,
                  I0 =>  \MDT13\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35117\ );

  -- Alias \WHOMP/\   
  \:54161\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54161\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54161\,
                   R => '0',
                   S => SYSRESET );

  \=54161\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54161\,
                  I0 =>  \CLXC\,
                  I1 =>  \WHOMP\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA02/\  
  \=54162\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54162\,
                  I0 =>  \WHOMP\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA04/\  
  \=54163\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54163\,
                  I0 =>  \WHOMP\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CO16\     
  \=54201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54201\,
                  I0 =>  \XUY16/\,
                  I1 =>  \54210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54202\,
                  I0 =>  \A2XG/\,
                  I1 =>  \54220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54203\,
                   R => '0',
                   S => SYSRESET );

  \=54203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54203\,
                  I0 =>  \MONEX\,
                  I1 =>  \54202\,
                  I2 =>  \54204\,
                  I3 =>  '0' );

  \=54204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54204\,
                  I0 =>  \54203\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=54205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54205\,
                  I0 =>  \WYHIG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54206\,
                  I0 =>  \WL13/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54207\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54207\,
                   R => '0',
                   S => SYSRESET );

  \=54207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54207\,
                  I0 =>  \54205\,
                  I1 =>  \54206\,
                  I2 =>  \54208\,
                  I3 =>  '0' );

  \=54208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54208\,
                  I0 =>  \54207\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54209\,
                  I0 =>  \54203\,
                  I1 =>  \54207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY14/\   
  \=54210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54210\,
                  I0 =>  \54204\,
                  I1 =>  \54208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54211\,
                  I0 =>  \CI14/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA14/\  
  \=54212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54212\,
                  I0 =>  \54209\,
                  I1 =>  \54210\,
                  I2 =>  \CI14/\,
                  I3 =>  '0' );

  \=54213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54213\,
                  I0 =>  \54209\,
                  I1 =>  \54210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI15/\    
  \=54214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54214\,
                  I0 =>  \54209\,
                  I1 =>  \54212\,
                  I2 =>  \CO14\,
                  I3 =>  '0' );

  -- Alias \SUMB14/\  
  \=54215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54215\,
                  I0 =>  \54213\,
                  I1 =>  \54211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54217\,
                  I0 =>  \54212\,
                  I1 =>  \54215\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=54218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54218\,
                  I0 =>  \WAG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54219\,
                  I0 =>  \WL16/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A14/\     
  \:54220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54220\,
                   R => '0',
                   S => SYSRESET );

  \=54220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54220\,
                  I0 =>  \54218\,
                  I1 =>  \54219\,
                  I2 =>  \54221\,
                  I3 =>  '0' );

  \=54221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54221\,
                  I0 =>  \54220\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54222\,
                  I0 =>  \RAG/\,
                  I1 =>  \54220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54257\    
  \=54223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54223\,
                  I0 =>  \54217\,
                  I1 =>  \54222\,
                  I2 =>  \CH14\,
                  I3 => \&54233\ );

  \=54224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54224\,
                  I0 =>  \WLG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54225\,
                  I0 =>  \WL02/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L14/\     
  \:54226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54226\,
                   R => '0',
                   S => SYSRESET );

  \=54226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54226\,
                  I0 =>  \54224\,
                  I1 =>  \54225\,
                  I2 =>  \54227\,
                  I3 =>  '0' );

  \=54227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54227\,
                  I0 =>  \54226\,
                  I1 =>  \CLG2G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54228\,
                  I0 =>  \RLG/\,
                  I1 =>  \54226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54229\,
                  I0 =>  \WQG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54230\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54230\,
                   R => '0',
                   S => SYSRESET );

  \=54230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54230\,
                  I0 =>  \54229\,
                  I1 =>  \54231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54231\,
                  I0 =>  \54230\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54232\,
                  I0 =>  \RQG/\,
                  I1 =>  \54230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54257\    
  \=54233\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54233\,
                  I0 =>  \54228\,
                  I1 =>  \54232\,
                  I2 =>  \54237\,
                  I3 => \&54258\ );

  \=54234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54234\,
                  I0 =>  \WZG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z14/\     
  \:54235\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54235\,
                   R => '0',
                   S => SYSRESET );

  \=54235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54235\,
                  I0 =>  \54234\,
                  I1 =>  \54236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54236\,
                  I0 =>  \54235\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54237\,
                  I0 =>  \RZG/\,
                  I1 =>  \54235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54238\,
                  I0 =>  \WBG/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54239\,
                   R => '0',
                   S => SYSRESET );

  \=54239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54239\,
                  I0 =>  \54238\,
                  I1 =>  \54240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54240\,
                  I0 =>  \54239\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54241\,
                  I0 =>  \RBHG/\,
                  I1 =>  \54239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54242\,
                  I0 =>  \54240\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54243\,
                  I0 =>  \WL13/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54244\,
                  I0 =>  \WL16/\,
                  I1 =>  \WG4G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54245\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54246\,
                  I0 =>  \WG1G/\,
                  I1 =>  \54254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54248\    
  \=54247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54247\,
                  I0 =>  \SA14\,
                  I1 =>  \54243\,
                  I2 =>  \54244\,
                  I3 =>  '0' );

  -- Alias \G14/\     
  \:54248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54248\,
                   R => '0',
                   S => SYSRESET );

  \=54248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54248\,
                  I0 =>  \54245\,
                  I1 =>  \54246\,
                  I2 =>  \54249\,
                  I3 => \&54247\ );

  -- Alias \G14\      
  \=54249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54249\,
                  I0 =>  \54248\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM14\    
  \=54250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54250\,
                  I0 =>  \54248\,
                  I1 =>  \54248\,
                  I2 =>  \54248\,
                  I3 =>  '0' );

  \=54251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54251\,
                  I0 =>  \RGG/\,
                  I1 =>  \54248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL14\     
  \=54252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54252\,
                  I0 =>  \54257\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL14\    
  \=54253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54253\,
                  I0 =>  \54257\,
                  I1 =>  \54257\,
                  I2 =>  \54257\,
                  I3 =>  '0' );

  -- Alias \WL14/\    
  \=54254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54254\,
                  I0 =>  \54252\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL14/\    
  \=54257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54257\,
                  I0 =>  \54241\,
                  I1 =>  \54242\,
                  I2 =>  \54251\,
                  I3 => \&54223\ );

  -- Alias \54257\    
  \=54258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54258\,
                  I0 =>  \MDT14\,
                  I1 =>  \R1C\,
                  I2 =>  '0',
                  I3 => \&35251\ );

  -- Alias \GTRST/\   
  \=54261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54261\,
                  I0 =>  \GTRST\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WHOMP\    
  \:54262\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \54262\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54262\,
                   R => SYSRESET,
                   S => '0' );

  \=54262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54262\,
                  I0 =>  \WHOMP/\,
                  I1 =>  \DVXP1\,
                  I2 =>  '0',
                  I3 => \&54263\ );

  -- Alias \WHOMP\    
  \=54263\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54263\,
                  I0 =>  \NISQ\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A11/2 - 4 BIT MODULE (4 OF 4).  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \CO02\     
  \=54301\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54301\,
                  I0 =>  \XUY02/\,
                  I1 =>  \54310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54302\,
                  I0 =>  \A2XG/\,
                  I1 =>  \54320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54303\,
                   R => '0',
                   S => SYSRESET );

  \=54303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54303\,
                  I0 =>  \MONEX\,
                  I1 =>  \54302\,
                  I2 =>  \54304\,
                  I3 =>  '0' );

  \=54304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54304\,
                  I0 =>  \54303\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=54305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54305\,
                  I0 =>  \WYHIG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54306\,
                  I0 =>  \WL16/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54307\,
                   R => '0',
                   S => SYSRESET );

  \=54307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54307\,
                  I0 =>  \54305\,
                  I1 =>  \54306\,
                  I2 =>  \54308\,
                  I3 =>  '0' );

  \=54308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54308\,
                  I0 =>  \54307\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54309\,
                  I0 =>  \54303\,
                  I1 =>  \54307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY16/\   
  \=54310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54310\,
                  I0 =>  \54304\,
                  I1 =>  \54308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54311\,
                  I0 =>  \CI16/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA16/\  
  \=54312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54312\,
                  I0 =>  \54309\,
                  I1 =>  \54310\,
                  I2 =>  \CI16/\,
                  I3 => \&54363\ );

  \=54313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54313\,
                  I0 =>  \54309\,
                  I1 =>  \54310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAC/\     
  \=54314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54314\,
                  I0 =>  \54309\,
                  I1 =>  \54312\,
                  I2 =>  \CO16\,
                  I3 =>  '0' );

  -- Alias \SUMB16/\  
  \=54315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54315\,
                  I0 =>  \54313\,
                  I1 =>  \54311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54317\,
                  I0 =>  \54312\,
                  I1 =>  \54315\,
                  I2 =>  \RUG/\,
                  I3 =>  '0' );

  \=54318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54318\,
                  I0 =>  \WAG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54319\,
                  I0 =>  \G16SW/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A16/\     
  \:54320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54320\,
                   R => '0',
                   S => SYSRESET );

  \=54320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54320\,
                  I0 =>  \54318\,
                  I1 =>  \54319\,
                  I2 =>  \54321\,
                  I3 =>  '0' );

  \=54321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54321\,
                  I0 =>  \54320\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54322\,
                  I0 =>  \RAG/\,
                  I1 =>  \54320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54357\    
  \=54323\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54323\,
                  I0 =>  \54317\,
                  I1 =>  \54322\,
                  I2 =>  \CH16\,
                  I3 => \&54333\ );

  \=54324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54324\,
                  I0 =>  \WLG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54325\,
                  I0 =>  \G16/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L16/\     
  \:54326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54326\,
                   R => '0',
                   S => SYSRESET );

  \=54326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54326\,
                  I0 =>  \54324\,
                  I1 =>  \54325\,
                  I2 =>  \54327\,
                  I3 => \&36460\ );

  \=54327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54327\,
                  I0 =>  \54326\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL16\     
  \=54328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54328\,
                  I0 =>  \RLG/\,
                  I1 =>  \54326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54329\,
                  I0 =>  \WQG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54330\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54330\,
                   R => '0',
                   S => SYSRESET );

  \=54330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54330\,
                  I0 =>  \54329\,
                  I1 =>  \54331\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54331\,
                  I0 =>  \54330\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54332\,
                  I0 =>  \RQG/\,
                  I1 =>  \54330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54357\    
  \=54333\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54333\,
                  I0 =>  \54328\,
                  I1 =>  \54332\,
                  I2 =>  \54337\,
                  I3 => \&54358\ );

  \=54334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54334\,
                  I0 =>  \WZG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z16/\     
  \:54335\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54335\,
                   R => '0',
                   S => SYSRESET );

  \=54335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54335\,
                  I0 =>  \54334\,
                  I1 =>  \54336\,
                  I2 =>  '0',
                  I3 => \&39413\ );

  \=54336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54336\,
                  I0 =>  \54335\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54337\,
                  I0 =>  \RZG/\,
                  I1 =>  \54335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54338\,
                  I0 =>  \WBG/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54339\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54339\,
                   R => '0',
                   S => SYSRESET );

  \=54339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54339\,
                  I0 =>  \54338\,
                  I1 =>  \54340\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54340\,
                  I0 =>  \54339\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54341\,
                  I0 =>  \RBHG/\,
                  I1 =>  \54339\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54342\,
                  I0 =>  \54340\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54343\,
                  I0 =>  \WL14/\,
                  I1 =>  \WG3G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54344\,
                  I0 =>  \WL01/\,
                  I1 =>  \WG5G/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54345\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54346\,
                  I0 =>  \WG2G/\,
                  I1 =>  \54354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54348\    
  \=54347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54347\,
                  I0 =>  \SA16\,
                  I1 =>  \54343\,
                  I2 =>  \54344\,
                  I3 =>  '0' );

  -- Alias \G16/\     
  \:54348\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54348\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54348\,
                   R => '0',
                   S => SYSRESET );

  \=54348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54348\,
                  I0 =>  \54345\,
                  I1 =>  \54346\,
                  I2 =>  \54349\,
                  I3 => \&54347\ );

  -- Alias \G16\      
  \=54349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54349\,
                  I0 =>  \54348\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEM16\    
  \=54350\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54350\,
                  I0 =>  \54348\,
                  I1 =>  \54348\,
                  I2 =>  \54348\,
                  I3 =>  '0' );

  \=54351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54351\,
                  I0 =>  \RGG/\,
                  I1 =>  \54348\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL16\     
  \=54352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54352\,
                  I0 =>  \54357\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL16\    
  \=54353\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54353\,
                  I0 =>  \54357\,
                  I1 =>  \54357\,
                  I2 =>  \54357\,
                  I3 =>  '0' );

  -- Alias \WL16/\    
  \=54354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54354\,
                  I0 =>  \54352\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL16/\    
  \=54357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54357\,
                  I0 =>  \54341\,
                  I1 =>  \54342\,
                  I2 =>  \54351\,
                  I3 => \&54323\ );

  -- Alias \54357\    
  \=54358\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54358\,
                  I0 =>  \MDT16\,
                  I1 =>  \R1C\,
                  I2 =>  \US2SG\,
                  I3 => \&35106\ );

  -- Alias \PIPAZ+/\  
  \=54361\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54361\,
                  I0 =>  \PIPAZ+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPAZ-/\  
  \=54362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54362\,
                  I0 =>  \PIPAZ-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA16/\  
  \=54363\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54363\,
                  I0 =>  \WHOMPA\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CO02\     
  \=54401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54401\,
                  I0 =>  \XUY01/\,
                  I1 =>  \54410\,
                  I2 =>  \CI15/\,
                  I3 => \&54301\ );

  \=54402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54402\,
                  I0 =>  \A2XG/\,
                  I1 =>  \54420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54403\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54403\,
                   R => '0',
                   S => SYSRESET );

  \=54403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54403\,
                  I0 =>  \BXVX\,
                  I1 =>  \54402\,
                  I2 =>  \54404\,
                  I3 =>  '0' );

  \=54404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54404\,
                  I0 =>  \54403\,
                  I1 =>  \CLXC\,
                  I2 =>  \CUG\,
                  I3 =>  '0' );

  \=54405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54405\,
                  I0 =>  \WYHIG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54406\,
                  I0 =>  \WL14/\,
                  I1 =>  \WYDG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54407\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54407\,
                   R => '0',
                   S => SYSRESET );

  \=54407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54407\,
                  I0 =>  \54405\,
                  I1 =>  \54406\,
                  I2 =>  \54408\,
                  I3 =>  '0' );

  \=54408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54408\,
                  I0 =>  \54407\,
                  I1 =>  \CUG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54409\,
                  I0 =>  \54403\,
                  I1 =>  \54407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XUY15/\   
  \=54410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54410\,
                  I0 =>  \54404\,
                  I1 =>  \54408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54411\,
                  I0 =>  \CI15/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA15/\  
  \=54412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54412\,
                  I0 =>  \54409\,
                  I1 =>  \CI15/\,
                  I2 =>  \54410\,
                  I3 =>  '0' );

  \=54413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54413\,
                  I0 =>  \54409\,
                  I1 =>  \54410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI16/\    
  \=54414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54414\,
                  I0 =>  \54409\,
                  I1 =>  \54412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMB15/\  
  \=54415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54415\,
                  I0 =>  \54413\,
                  I1 =>  \54411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54417\,
                  I0 =>  \54412\,
                  I1 =>  \54415\,
                  I2 =>  \RULOG/\,
                  I3 =>  '0' );

  \=54418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54418\,
                  I0 =>  \WAG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54419\,
                  I0 =>  \G16SW/\,
                  I1 =>  \WALSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \A15/\     
  \:54420\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54420\,
                   R => '0',
                   S => SYSRESET );

  \=54420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54420\,
                  I0 =>  \54418\,
                  I1 =>  \54419\,
                  I2 =>  \54421\,
                  I3 =>  '0' );

  \=54421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54421\,
                  I0 =>  \54420\,
                  I1 =>  \CAG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54422\,
                  I0 =>  \RAG/\,
                  I1 =>  \54420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54457\    
  \=54423\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54423\,
                  I0 =>  \54417\,
                  I1 =>  \54422\,
                  I2 =>  \CH16\,
                  I3 => \&54433\ );

  \=54424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54424\,
                  I0 =>  \WLG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54425\,
                  I0 =>  \G01/\,
                  I1 =>  \G2LSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L15/\     
  \:54426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54426\,
                   R => '0',
                   S => SYSRESET );

  \=54426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54426\,
                  I0 =>  \54424\,
                  I1 =>  \54425\,
                  I2 =>  \54427\,
                  I3 =>  '0' );

  \=54427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54427\,
                  I0 =>  \54426\,
                  I1 =>  \CLG1G\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54429\,
                  I0 =>  \WQG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54430\,
                   R => '0',
                   S => SYSRESET );

  \=54430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54430\,
                  I0 =>  \54429\,
                  I1 =>  \54431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54431\,
                  I0 =>  \54430\,
                  I1 =>  \CQG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54432\,
                  I0 =>  \RQG/\,
                  I1 =>  \54430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54457\    
  \=54433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54433\,
                  I0 =>  '0',
                  I1 =>  \54432\,
                  I2 =>  \54437\,
                  I3 => \&54458\ );

  \=54434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54434\,
                  I0 =>  \WZG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \Z15/\     
  \:54435\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54435\,
                   R => '0',
                   S => SYSRESET );

  \=54435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54435\,
                  I0 =>  \54434\,
                  I1 =>  \54436\,
                  I2 =>  '0',
                  I3 => \&39433\ );

  \=54436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54436\,
                  I0 =>  \54435\,
                  I1 =>  \CZG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54437\,
                  I0 =>  \RZG/\,
                  I1 =>  \54435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54438\,
                  I0 =>  \WBG/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:54439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54439\,
                   R => '0',
                   S => SYSRESET );

  \=54439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54439\,
                  I0 =>  \54438\,
                  I1 =>  \54440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54440\,
                  I0 =>  \54439\,
                  I1 =>  \CBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54441\,
                  I0 =>  \RBHG/\,
                  I1 =>  \54439\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54442\,
                  I0 =>  \54440\,
                  I1 =>  \RCG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54443\,
                  I0 =>  '0',
                  I1 =>  \ONE\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54444\,
                  I0 =>  '0',
                  I1 =>  \ONE\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54445\,
                  I0 =>  \L2GDG/\,
                  I1 =>  \L14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54446\,
                  I0 =>  \WG1G/\,
                  I1 =>  \54454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \54448\    
  \=54447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54447\,
                  I0 =>  \SA16\,
                  I1 =>  \54443\,
                  I2 =>  \54444\,
                  I3 =>  '0' );

  -- Alias \G15/\     
  \:54448\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \54448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$54448\,
                   R => '0',
                   S => SYSRESET );

  \=54448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$54448\,
                  I0 =>  \54445\,
                  I1 =>  \54446\,
                  I2 =>  \54449\,
                  I3 => \&54447\ );

  -- Alias \G15\      
  \=54449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54449\,
                  I0 =>  \54448\,
                  I1 =>  \CGG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=54451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54451\,
                  I0 =>  \RGG/\,
                  I1 =>  \54448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WL15\     
  \=54452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54452\,
                  I0 =>  \54457\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL15\    
  \=54453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54453\,
                  I0 =>  \54457\,
                  I1 =>  \54457\,
                  I2 =>  \54457\,
                  I3 =>  '0' );

  -- Alias \WL15/\    
  \=54454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54454\,
                  I0 =>  \54452\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL15/\    
  \=54457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54457\,
                  I0 =>  \54441\,
                  I1 =>  \54442\,
                  I2 =>  \54451\,
                  I3 => \&53363\ );

  -- Alias \54457\    
  \=54458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54458\,
                  I0 =>  \MDT15\,
                  I1 =>  \R1C\,
                  I2 =>  \RL16\,
                  I3 =>  '0' );

  -- Alias \PIPAY-/\  
  \=54461\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \54461\,
                  I0 =>  \PIPAY-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA07/\  
  \=54462\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54462\,
                  I0 =>  \WHOMP\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SUMA12/\  
  \=54463\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&54463\,
                  I0 =>  \WHOMP\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A12/1 - PARITY AND S REGISTER.  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \G01A/\    
  \=34101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34101\,
                  I0 =>  \G01\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34102\,
                  I0 =>  \G02\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34103\,
                  I0 =>  \G03\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34104\,
                  I0 =>  \G01\,
                  I1 =>  \G02\,
                  I2 =>  \G03\,
                  I3 =>  '0' );

  \=34105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34105\,
                  I0 =>  \G01\,
                  I1 =>  \34102\,
                  I2 =>  \34103\,
                  I3 =>  '0' );

  \=34106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34106\,
                  I0 =>  \34101\,
                  I1 =>  \G02\,
                  I2 =>  \34103\,
                  I3 =>  '0' );

  \=34107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34107\,
                  I0 =>  \34101\,
                  I1 =>  \34102\,
                  I2 =>  \G03\,
                  I3 =>  '0' );

  -- Alias \PA03\     
  \=34108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34108\,
                  I0 =>  \34104\,
                  I1 =>  \34105\,
                  I2 =>  '0',
                  I3 => \&34109\ );

  -- Alias \34108\    
  \=34109\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34109\,
                  I0 =>  \34106\,
                  I1 =>  \34107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PA03/\    
  \=34110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34110\,
                  I0 =>  \34108\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34111\,
                  I0 =>  \G04\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34112\,
                  I0 =>  \G05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34113\,
                  I0 =>  \G06\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34114\,
                  I0 =>  \G04\,
                  I1 =>  \G05\,
                  I2 =>  \G06\,
                  I3 =>  '0' );

  \=34115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34115\,
                  I0 =>  \G04\,
                  I1 =>  \34112\,
                  I2 =>  \34113\,
                  I3 =>  '0' );

  \=34116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34116\,
                  I0 =>  \34111\,
                  I1 =>  \G05\,
                  I2 =>  \34113\,
                  I3 =>  '0' );

  \=34117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34117\,
                  I0 =>  \34111\,
                  I1 =>  \34112\,
                  I2 =>  \G06\,
                  I3 =>  '0' );

  -- Alias \PA06\     
  \=34118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34118\,
                  I0 =>  \34114\,
                  I1 =>  \34115\,
                  I2 =>  '0',
                  I3 => \&34119\ );

  -- Alias \34118\    
  \=34119\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34119\,
                  I0 =>  \34116\,
                  I1 =>  \34117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PA06/\    
  \=34120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34120\,
                  I0 =>  \34118\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34121\,
                  I0 =>  \34114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34122\,
                  I0 =>  \G07\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34123\,
                  I0 =>  \G08\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34124\,
                  I0 =>  \G09\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34125\,
                  I0 =>  \G07\,
                  I1 =>  \G08\,
                  I2 =>  \G09\,
                  I3 =>  '0' );

  \=34126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34126\,
                  I0 =>  \G07\,
                  I1 =>  \34123\,
                  I2 =>  \34124\,
                  I3 =>  '0' );

  \=34127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34127\,
                  I0 =>  \34122\,
                  I1 =>  \G08\,
                  I2 =>  \34124\,
                  I3 =>  '0' );

  \=34128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34128\,
                  I0 =>  \34122\,
                  I1 =>  \34123\,
                  I2 =>  \G09\,
                  I3 =>  '0' );

  -- Alias \PA09\     
  \=34129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34129\,
                  I0 =>  \34125\,
                  I1 =>  \34126\,
                  I2 =>  '0',
                  I3 => \&34130\ );

  -- Alias \34129\    
  \=34130\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34130\,
                  I0 =>  \34127\,
                  I1 =>  \34128\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PA09/\    
  \=34131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34131\,
                  I0 =>  \34129\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34132\,
                  I0 =>  \34125\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34133\,
                  I0 =>  \G10\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34134\,
                  I0 =>  \G11\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34135\,
                  I0 =>  \G12\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34136\,
                  I0 =>  \G10\,
                  I1 =>  \G11\,
                  I2 =>  \G12\,
                  I3 =>  '0' );

  \=34137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34137\,
                  I0 =>  \G10\,
                  I1 =>  \34134\,
                  I2 =>  \34135\,
                  I3 =>  '0' );

  \=34138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34138\,
                  I0 =>  \34133\,
                  I1 =>  \G11\,
                  I2 =>  \34135\,
                  I3 =>  '0' );

  \=34139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34139\,
                  I0 =>  \34133\,
                  I1 =>  \34134\,
                  I2 =>  \G12\,
                  I3 =>  '0' );

  -- Alias \PA12\     
  \=34140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34140\,
                  I0 =>  \34136\,
                  I1 =>  \34137\,
                  I2 =>  '0',
                  I3 => \&34141\ );

  -- Alias \34140\    
  \=34141\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34141\,
                  I0 =>  \34138\,
                  I1 =>  \34139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34142\,
                  I0 =>  \34136\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PA12/\    
  \=34143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34143\,
                  I0 =>  \34140\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34144\,
                  I0 =>  \G13\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34145\,
                  I0 =>  \G14\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G16A/\    
  \=34146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34146\,
                  I0 =>  \G16\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34147\,
                  I0 =>  \G13\,
                  I1 =>  \G14\,
                  I2 =>  \G16\,
                  I3 =>  '0' );

  \=34148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34148\,
                  I0 =>  \G13\,
                  I1 =>  \34145\,
                  I2 =>  \34146\,
                  I3 =>  '0' );

  \=34149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34149\,
                  I0 =>  \34144\,
                  I1 =>  \G14\,
                  I2 =>  \34146\,
                  I3 =>  '0' );

  \=34150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34150\,
                  I0 =>  \34144\,
                  I1 =>  \34145\,
                  I2 =>  \G16\,
                  I3 =>  '0' );

  -- Alias \PA15\     
  \=34151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34151\,
                  I0 =>  \34147\,
                  I1 =>  \34148\,
                  I2 =>  '0',
                  I3 => \&34152\ );

  -- Alias \34151\    
  \=34152\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34152\,
                  I0 =>  \34149\,
                  I1 =>  \34150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PA15/\    
  \=34153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34153\,
                  I0 =>  \34151\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34154\,
                  I0 =>  \34147\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GNZRO\    
  \=34155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34155\,
                  I0 =>  \34142\,
                  I1 =>  \34154\,
                  I2 =>  '0',
                  I3 => \&34156\ );

  -- Alias \34155\    
  \=34156\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34156\,
                  I0 =>  \34121\,
                  I1 =>  \34132\,
                  I2 =>  '0',
                  I3 => \&34157\ );

  -- Alias \GNZRO\    
  \=34157\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34157\,
                  I0 =>  \G15\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSC/\     
  \=34158\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34158\,
                  I0 =>  '0',
                  I1 =>  \BRXP3\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WG/\      
  \=34159\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34159\,
                  I0 =>  '0',
                  I1 =>  \BRXP3\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34201\,
                  I0 =>  \TSUDO/\,
                  I1 =>  \T7PHS4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34202\,
                  I0 =>  \34201\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34203\,
                  I0 =>  \34105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34204\,
                  I0 =>  \34155\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EXTPLS\   
  \=34205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34205\,
                  I0 =>  \34203\,
                  I1 =>  \34204\,
                  I2 =>  \34202\,
                  I3 =>  '0' );

  -- Alias \RELPLS\   
  \=34206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34206\,
                  I0 =>  \34204\,
                  I1 =>  \34202\,
                  I2 =>  \G01A/\,
                  I3 => \&34207\ );

  -- Alias \34206\    
  \=34207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34207\,
                  I0 =>  \34102\,
                  I1 =>  \G03\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \34209\    
  \=34208\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34208\,
                  I0 =>  \34205\,
                  I1 =>  \34206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34209\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34209\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34209\,
                   R => '0',
                   S => SYSRESET );

  \=34209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34209\,
                  I0 =>  \34215\,
                  I1 =>  \34210\,
                  I2 =>  '0',
                  I3 => \&34208\ );

  \=34210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34210\,
                  I0 =>  \34209\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34211\,
                  I0 =>  \RAD\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RADRZ\    
  \=34212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34212\,
                  I0 =>  \34209\,
                  I1 =>  \34211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RADRG\    
  \=34213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34213\,
                  I0 =>  \34211\,
                  I1 =>  \34210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \34215\    
  \=34214\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34214\,
                  I0 =>  \34204\,
                  I1 =>  \G01\,
                  I2 =>  \34202\,
                  I3 =>  '0' );

  -- Alias \INHPLS\   
  \=34215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34215\,
                  I0 =>  \G02\,
                  I1 =>  \34103\,
                  I2 =>  '0',
                  I3 => \&34214\ );

  \=34216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34216\,
                  I0 =>  \34204\,
                  I1 =>  \G02\,
                  I2 =>  '0',
                  I3 => \&34217\ );

  -- Alias \34216\    
  \=34217\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34217\,
                  I0 =>  \G01\,
                  I1 =>  \G03\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEQZRO/\  
  \=34218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34218\,
                  I0 =>  \34216\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34219\,
                  I0 =>  \EB9\,
                  I1 =>  \S10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34220\,
                  I0 =>  \EB10\,
                  I1 =>  \S09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAD09\    
  \=34221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34221\,
                  I0 =>  \S09/\,
                  I1 =>  \34219\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAD10\    
  \=34222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34222\,
                  I0 =>  \S10/\,
                  I1 =>  \34220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAD11\    
  \=34223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34223\,
                  I0 =>  \S10/\,
                  I1 =>  \S09/\,
                  I2 =>  \EB11/\,
                  I3 =>  '0' );

  -- Alias \EAD09/\   
  \=34224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34224\,
                  I0 =>  \34221\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAD10/\   
  \=34225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34225\,
                  I0 =>  \34222\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EAD11/\   
  \=34226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34226\,
                  I0 =>  \34223\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34227\,
                  I0 =>  \PA03\,
                  I1 =>  \PA06\,
                  I2 =>  \PA09\,
                  I3 =>  '0' );

  \=34228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34228\,
                  I0 =>  \PA03\,
                  I1 =>  \PA06/\,
                  I2 =>  \PA09/\,
                  I3 =>  '0' );

  \=34229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34229\,
                  I0 =>  \PA03/\,
                  I1 =>  \PA06\,
                  I2 =>  \PA09/\,
                  I3 =>  '0' );

  \=34230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34230\,
                  I0 =>  \PA03/\,
                  I1 =>  \PA06/\,
                  I2 =>  \PA09\,
                  I3 =>  '0' );

  -- Alias \PB09\     
  \=34231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34231\,
                  I0 =>  \34227\,
                  I1 =>  \34228\,
                  I2 =>  '0',
                  I3 => \&34232\ );

  -- Alias \34231\    
  \=34232\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34232\,
                  I0 =>  \34229\,
                  I1 =>  \34230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PB09/\    
  \=34233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34233\,
                  I0 =>  \34231\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34234\,
                  I0 =>  \PA12\,
                  I1 =>  \PA15\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34235\,
                  I0 =>  \PA12/\,
                  I1 =>  \PA15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PB15\     
  \=34236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34236\,
                  I0 =>  \34234\,
                  I1 =>  \34235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PB15/\    
  \=34237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34237\,
                  I0 =>  \34236\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34238\,
                  I0 =>  \34233\,
                  I1 =>  \34236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34239\,
                  I0 =>  \34231\,
                  I1 =>  \34237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PC15\     
  \=34240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34240\,
                  I0 =>  \34238\,
                  I1 =>  \34239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MGP/\     
  \=34241\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34241\,
                  I0 =>  \34240\,
                  I1 =>  \34240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PC15/\    
  \=34242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34242\,
                  I0 =>  \34240\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GEMP\     
  \=34243\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34243\,
                  I0 =>  \34242\,
                  I1 =>  \34242\,
                  I2 =>  \34242\,
                  I3 =>  '0' );

  -- Alias \MSP\      
  \=34244\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34244\,
                  I0 =>  \34245\,
                  I1 =>  \34245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34245\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34245\,
                   R => '0',
                   S => SYSRESET );

  \=34245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34245\,
                  I0 =>  \34246\,
                  I1 =>  \MONPAR\,
                  I2 =>  \SAP\,
                  I3 =>  '0' );

  \=34246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34246\,
                  I0 =>  \CGG\,
                  I1 =>  \34245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34247\,
                  I0 =>  \34242\,
                  I1 =>  \34245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34248\,
                  I0 =>  \34246\,
                  I1 =>  \34240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \34251\    
  \=34250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34250\,
                  I0 =>  \TPARG/\,
                  I1 =>  \8XP5\,
                  I2 =>  \34247\,
                  I3 =>  '0' );

  -- Alias \PALE\     
  \=34251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34251\,
                  I0 =>  \SCAD\,
                  I1 =>  \34248\,
                  I2 =>  \GOJAM\,
                  I3 => \&34250\ );

  -- Alias \MPAL/\    
  \=34252\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34252\,
                  I0 =>  \34251\,
                  I1 =>  \34251\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BRXP3\    
  \=34253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34253\,
                  I0 =>  \IC15/\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSCDBL/\  
  \=34254\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34254\,
                  I0 =>  \SCADBL\,
                  I1 =>  \SCADBL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************************
  -- ***                                  ***
  -- ***  A12/2 - PARITY AND S REGISTER.  ***
  -- ***                                  ***
  -- ****************************************

  -- Alias \G01ED\    
  \=34301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34301\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34302\,
                  I0 =>  \WL08/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34303\,
                   R => '0',
                   S => SYSRESET );

  \=34303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34303\,
                  I0 =>  \34302\,
                  I1 =>  \34304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34304\,
                  I0 =>  \34303\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S08\      
  \=34306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34306\,
                  I0 =>  \34303\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S08/\     
  \=34307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34307\,
                  I0 =>  \34304\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G02ED\    
  \=34309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34309\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34310\,
                  I0 =>  \WL09/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34311\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34311\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34311\,
                   R => '0',
                   S => SYSRESET );

  \=34311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34311\,
                  I0 =>  \34310\,
                  I1 =>  \34312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34312\,
                  I0 =>  \34311\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S09\      
  \=34314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34314\,
                  I0 =>  \34311\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S09/\     
  \=34315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34315\,
                  I0 =>  \34312\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G03ED\    
  \=34317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34317\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34318\,
                  I0 =>  \WL10/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34319\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34319\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34319\,
                   R => '0',
                   S => SYSRESET );

  \=34319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34319\,
                  I0 =>  \34318\,
                  I1 =>  \34320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34320\,
                  I0 =>  \34319\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S10\      
  \=34322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34322\,
                  I0 =>  \34319\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S10/\     
  \=34323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34323\,
                  I0 =>  \34320\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G04ED\    
  \=34325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34325\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34326\,
                  I0 =>  \WL11/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34327\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34327\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34327\,
                   R => '0',
                   S => SYSRESET );

  \=34327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34327\,
                  I0 =>  \34326\,
                  I1 =>  \34328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34328\,
                  I0 =>  \34327\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T12A\     
  \=34329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34329\,
                  I0 =>  \T12/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S11\      
  \=34330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34330\,
                  I0 =>  \34327\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S11/\     
  \=34331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34331\,
                  I0 =>  \34328\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G05ED\    
  \=34333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34333\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34334\,
                  I0 =>  \WL12/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34335\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34335\,
                   R => '0',
                   S => SYSRESET );

  \=34335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34335\,
                  I0 =>  \8XP5\,
                  I1 =>  \34334\,
                  I2 =>  \34336\,
                  I3 =>  '0' );

  \=34336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34336\,
                  I0 =>  \34335\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S12\      
  \=34338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34338\,
                  I0 =>  \34335\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S12/\     
  \=34339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34339\,
                  I0 =>  \34336\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHIFT/\   
  \=34340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34340\,
                  I0 =>  \SHINC\,
                  I1 =>  \SHANC\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G06ED\    
  \=34341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34341\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G07ED\    
  \=34342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34342\,
                  I0 =>  \WEDOPG/\,
                  I1 =>  \WL14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34343\,
                  I0 =>  \OCTAD2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34344\,
                  I0 =>  \XB0/\,
                  I1 =>  \T02/\,
                  I2 =>  \34343\,
                  I3 =>  '0' );

  \=34345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34345\,
                  I0 =>  \34343\,
                  I1 =>  \T02/\,
                  I2 =>  \XB1/\,
                  I3 =>  '0' );

  \=34346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34346\,
                  I0 =>  \34343\,
                  I1 =>  \T02/\,
                  I2 =>  \XB2/\,
                  I3 =>  '0' );

  \=34347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34347\,
                  I0 =>  \34343\,
                  I1 =>  \T02/\,
                  I2 =>  \XB3/\,
                  I3 =>  '0' );

  -- Alias \CYR/\     
  \:34348\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34348\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34348\,
                   R => '0',
                   S => SYSRESET );

  \=34348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34348\,
                  I0 =>  \34344\,
                  I1 =>  \34349\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34349\,
                  I0 =>  \34348\,
                  I1 =>  \34329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SR/\      
  \:34350\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34350\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34350\,
                   R => '0',
                   S => SYSRESET );

  \=34350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34350\,
                  I0 =>  \34345\,
                  I1 =>  \34351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34351\,
                  I0 =>  \34350\,
                  I1 =>  \34329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CYL/\     
  \:34352\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34352\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34352\,
                   R => '0',
                   S => SYSRESET );

  \=34352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34352\,
                  I0 =>  \34346\,
                  I1 =>  \34353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34353\,
                  I0 =>  \34352\,
                  I1 =>  \34329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EDOP/\    
  \:34354\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34354\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34354\,
                   R => '0',
                   S => SYSRESET );

  \=34354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34354\,
                  I0 =>  \34347\,
                  I1 =>  \34355\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34355\,
                  I0 =>  \34354\,
                  I1 =>  \34329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34356\,
                  I0 =>  \34349\,
                  I1 =>  \34351\,
                  I2 =>  '0',
                  I3 => \&34357\ );

  -- Alias \34356\    
  \=34357\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34357\,
                  I0 =>  \34353\,
                  I1 =>  \34355\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GINH\     
  \=34358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34358\,
                  I0 =>  \34356\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHIFT\    
  \=34362\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34362\,
                  I0 =>  \34340\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34401\,
                  I0 =>  \WL01/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34402\,
                   R => '0',
                   S => SYSRESET );

  \=34402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34402\,
                  I0 =>  \34401\,
                  I1 =>  \34403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34403\,
                  I0 =>  \34402\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S01\      
  \=34404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34404\,
                  I0 =>  \34402\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S01/\     
  \=34406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34406\,
                  I0 =>  \34403\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34408\,
                  I0 =>  \WL02/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34409\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34409\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34409\,
                   R => '0',
                   S => SYSRESET );

  \=34409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34409\,
                  I0 =>  \34408\,
                  I1 =>  \34410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34410\,
                  I0 =>  \34409\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S02\      
  \=34411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34411\,
                  I0 =>  \34409\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S02/\     
  \=34413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34413\,
                  I0 =>  \34410\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34415\,
                  I0 =>  \WL03/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34416\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34416\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34416\,
                   R => '0',
                   S => SYSRESET );

  \=34416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34416\,
                  I0 =>  \34415\,
                  I1 =>  \34417\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34417\,
                  I0 =>  \34416\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S03\      
  \=34418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34418\,
                  I0 =>  \34416\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S03/\     
  \=34420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34420\,
                  I0 =>  \34417\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34422\,
                  I0 =>  \WL04/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34423\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34423\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34423\,
                   R => '0',
                   S => SYSRESET );

  \=34423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34423\,
                  I0 =>  \34422\,
                  I1 =>  \34424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34424\,
                  I0 =>  \34423\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S04\      
  \=34425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34425\,
                  I0 =>  \34423\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S04/\     
  \=34427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34427\,
                  I0 =>  \34424\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34429\,
                  I0 =>  \WL05/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34430\,
                   R => '0',
                   S => SYSRESET );

  \=34430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34430\,
                  I0 =>  \34429\,
                  I1 =>  \34431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34431\,
                  I0 =>  \34430\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S05\      
  \=34432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34432\,
                  I0 =>  \34430\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S05/\     
  \=34434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34434\,
                  I0 =>  \34431\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34436\,
                  I0 =>  \WL06/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34437\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34437\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34437\,
                   R => '0',
                   S => SYSRESET );

  \=34437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34437\,
                  I0 =>  \34436\,
                  I1 =>  \34438\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34438\,
                  I0 =>  \34437\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S06\      
  \=34439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34439\,
                  I0 =>  \34437\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S06/\     
  \=34441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34441\,
                  I0 =>  \34438\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34443\,
                  I0 =>  \WL07/\,
                  I1 =>  \WSG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:34444\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \34444\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$34444\,
                   R => '0',
                   S => SYSRESET );

  \=34444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$34444\,
                  I0 =>  \34443\,
                  I1 =>  \34445\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34445\,
                  I0 =>  \34444\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WGA/\     
  \=34446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34446\,
                  I0 =>  \34467\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S07\      
  \=34447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34447\,
                  I0 =>  \34444\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S07/\     
  \=34449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34449\,
                  I0 =>  \34445\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL03/\    
  \=34450\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34450\,
                  I0 =>  \R6\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35359\ );

  -- Alias \RL04/\    
  \=34451\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34451\,
                  I0 =>  \CAD4\,
                  I1 =>  \RPTAD4\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL05/\    
  \=34452\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34452\,
                  I0 =>  \CAD5\,
                  I1 =>  \RPTAD5\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL06/\    
  \=34453\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&34453\,
                  I0 =>  \CAD6\,
                  I1 =>  \RPTAD6\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34462\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34462\,
                  I0 =>  \L02/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L02A/\    
  \=34463\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34463\,
                  I0 =>  \34462\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34464\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34464\,
                  I0 =>  \L15/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \L15A/\    
  \=34465\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34465\,
                  I0 =>  \34464\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \G01A\     
  \=34466\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34466\,
                  I0 =>  \G01A/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=34467\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \34467\,
                  I0 =>  \WG/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *************************
  -- ***                   ***
  -- ***  A13/1 - ALARMS.  ***
  -- ***                   ***
  -- *************************

  \=41101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41101\,
                  I0 =>  \MSTRT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41102\,
                  I0 =>  \F05B/\,
                  I1 =>  \41101\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41103\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41103\,
                   R => '0',
                   S => SYSRESET );

  \=41103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41103\,
                  I0 =>  \41102\,
                  I1 =>  \41104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41104\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41104\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41104\,
                   R => SYSRESET,
                   S => '0' );

  \=41104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41104\,
                  I0 =>  \41103\,
                  I1 =>  \41101\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSTRTP\   
  \=41105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41105\,
                  I0 =>  \F05A/\,
                  I1 =>  \41103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MPIPAL/\  
  \=41106\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41106\,
                  I0 =>  \PIPAFL\,
                  I1 =>  \PIPAFL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41107\,
                   R => '0',
                   S => SYSRESET );

  \=41107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41107\,
                  I0 =>  \IIP\,
                  I1 =>  \41108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41108\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41108\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41108\,
                   R => SYSRESET,
                   S => '0' );

  \=41108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41108\,
                  I0 =>  \41107\,
                  I1 =>  \F14B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41109\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41109\,
                   R => '0',
                   S => SYSRESET );

  \=41109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41109\,
                  I0 =>  \IIP/\,
                  I1 =>  \41110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41110\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41110\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41110\,
                   R => SYSRESET,
                   S => '0' );

  \=41110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41110\,
                  I0 =>  \41109\,
                  I1 =>  \F14B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41111\,
                  I0 =>  \F14H\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41112\,
                  I0 =>  \41108\,
                  I1 =>  \41111\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41113\,
                  I0 =>  \41111\,
                  I1 =>  \41110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRPTAL/\  
  \=41114\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41114\,
                  I0 =>  \41112\,
                  I1 =>  \41112\,
                  I2 =>  \41113\,
                  I3 => \&41115\ );

  -- Alias \MRPTAL/\  
  \=41115\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41115\,
                  I0 =>  \41113\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \41117\    
  \=41116\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41116\,
                  I0 =>  \PALE\,
                  I1 =>  \41112\,
                  I2 =>  \41113\,
                  I3 =>  '0' );

  -- Alias \CKTAL/\   
  \=41117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41117\,
                  I0 =>  \41125\,
                  I1 =>  \41126\,
                  I2 =>  \WATCHP\,
                  I3 => \&41116\ );

  -- Alias \ALGA\     
  \=41118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41118\,
                  I0 =>  \NHALGA\,
                  I1 =>  \41117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41119\,
                  I0 =>  \TCF0\,
                  I1 =>  \TC0\,
                  I2 =>  '0',
                  I3 => \&41120\ );

  -- Alias \41119\    
  \=41120\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41120\,
                  I0 =>  \INKL\,
                  I1 =>  \T04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41121\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41121\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41121\,
                   R => SYSRESET,
                   S => '0' );

  \=41121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41121\,
                  I0 =>  \TC0\,
                  I1 =>  \TCF0\,
                  I2 =>  \41122\,
                  I3 =>  '0' );

  \:41122\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41122\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41122\,
                   R => '0',
                   S => SYSRESET );

  \=41122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41122\,
                  I0 =>  \41121\,
                  I1 =>  \F10B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41123\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41123\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41123\,
                   R => SYSRESET,
                   S => '0' );

  \=41123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41123\,
                  I0 =>  \41119\,
                  I1 =>  \41124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41124\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41124\,
                   R => '0',
                   S => SYSRESET );

  \=41124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41124\,
                  I0 =>  \41123\,
                  I1 =>  \F10B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41125\,
                  I0 =>  \F10A/\,
                  I1 =>  \41122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41126\,
                  I0 =>  \F10A/\,
                  I1 =>  \41124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MTCAL/\   
  \=41127\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41127\,
                  I0 =>  \41125\,
                  I1 =>  \41125\,
                  I2 =>  \41126\,
                  I3 => \&41128\ );

  -- Alias \MTCAL/\   
  \=41128\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41128\,
                  I0 =>  \41126\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41129\,
                  I0 =>  \G01A\,
                  I1 =>  \G16A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41130\,
                  I0 =>  \SUMA16/\,
                  I1 =>  \SUMB16/\,
                  I2 =>  \G01A/\,
                  I3 =>  '0' );

  -- Alias \G16SW/\   
  \=41131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41131\,
                  I0 =>  \41129\,
                  I1 =>  \41130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \41134\    
  \=41132\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41132\,
                  I0 =>  \BMAGZM\,
                  I1 =>  \INLNKP\,
                  I2 =>  \INLNKM\,
                  I3 => \&41133\ );

  -- Alias \41134\    
  \=41133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41133\,
                  I0 =>  \RNRADP\,
                  I1 =>  \RNRADM\,
                  I2 =>  \GYROD\,
                  I3 => \&41135\ );

  -- Alias \CTPLS/\   
  \=41134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41134\,
                  I0 =>  \CDUXD\,
                  I1 =>  \CDUYD\,
                  I2 =>  \CDUZD\,
                  I3 => \&41132\ );

  -- Alias \41134\    
  \=41135\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41135\,
                  I0 =>  \TRUND\,
                  I1 =>  \SHAFTD\,
                  I2 =>  \THRSTD\,
                  I3 => \&41136\ );

  -- Alias \41134\    
  \=41136\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41136\,
                  I0 =>  \EMSD\,
                  I1 =>  \OTLNKM\,
                  I2 =>  \ALTM\,
                  I3 => \&49435\ );

  \=41137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41137\,
                  I0 =>  \41134\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41138\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41138\,
                   R => '0',
                   S => SYSRESET );

  \=41138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41138\,
                  I0 =>  \41137\,
                  I1 =>  \41139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41139\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41139\,
                   R => SYSRESET,
                   S => '0' );

  \=41139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41139\,
                  I0 =>  \41138\,
                  I1 =>  \INKL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41140\,
                  I0 =>  \NOTEST\,
                  I1 =>  \41138\,
                  I2 =>  \T09/\,
                  I3 =>  '0' );

  \:41141\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41141\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41141\,
                   R => '0',
                   S => SYSRESET );

  \=41141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41141\,
                  I0 =>  \41140\,
                  I1 =>  \41142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41142\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41142\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41142\,
                   R => SYSRESET,
                   S => '0' );

  \=41142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41142\,
                  I0 =>  \41141\,
                  I1 =>  \INKL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41143\,
                  I0 =>  \T03/\,
                  I1 =>  \41141\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MCTRAL/\  
  \=41144\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41144\,
                  I0 =>  \41143\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41145\ );

  -- Alias \MCTRAL/\  
  \=41145\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41145\,
                  I0 =>  \41143\,
                  I1 =>  \41151\,
                  I2 =>  \41151\,
                  I3 =>  '0' );

  \=41146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41146\,
                  I0 =>  \41143\,
                  I1 =>  \41151\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \DOFILT\   
  \=41147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41147\,
                  I0 =>  \41146\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41148\,
                  I0 =>  \T03/\,
                  I1 =>  \INKL\,
                  I2 =>  \CTROR\,
                  I3 =>  '0' );

  \:41149\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41149\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41149\,
                   R => '0',
                   S => SYSRESET );

  \=41149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41149\,
                  I0 =>  \41148\,
                  I1 =>  \41150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41150\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41150\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41150\,
                   R => SYSRESET,
                   S => '0' );

  \=41150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41150\,
                  I0 =>  \41149\,
                  I1 =>  \F07A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41151\,
                  I0 =>  \41150\,
                  I1 =>  \F07B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41152\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41152\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41152\,
                   R => '0',
                   S => SYSRESET );

  \=41152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41152\,
                  I0 =>  \DLKRPT\,
                  I1 =>  \41153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41153\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41153\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41153\,
                   R => SYSRESET,
                   S => '0' );

  \=41153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41153\,
                  I0 =>  \41152\,
                  I1 =>  \DRPRST\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \DLKPLS\   
  \=41154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41154\,
                  I0 =>  \T10/\,
                  I1 =>  \41152\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41201\,
                  I0 =>  \VFAIL\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41202\,
                  I0 =>  \F05B/\,
                  I1 =>  \41201\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41203\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41203\,
                   R => '0',
                   S => SYSRESET );

  \=41203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41203\,
                  I0 =>  \41202\,
                  I1 =>  \41204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41204\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41204\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41204\,
                   R => SYSRESET,
                   S => '0' );

  \=41204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41204\,
                  I0 =>  \41203\,
                  I1 =>  \41201\,
                  I2 =>  \NHVFAL\,
                  I3 =>  '0' );

  \=41205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41205\,
                  I0 =>  \F05A/\,
                  I1 =>  \41203\,
                  I2 =>  \NHVFAL\,
                  I3 =>  '0' );

  \=41206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41206\,
                  I0 =>  \F05A/\,
                  I1 =>  \41203\,
                  I2 =>  \STNDBY/\,
                  I3 =>  '0' );

  -- Alias \MVFAIL/\  
  \=41207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41207\,
                  I0 =>  \41205\,
                  I1 =>  \41205\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \41211\    
  \=41208\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41208\,
                  I0 =>  \41206\,
                  I1 =>  \DOFILT\,
                  I2 =>  \SCADBL\,
                  I3 =>  '0' );

  \=41209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41209\,
                  I0 =>  \F14B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41210\,
                  I0 =>  \41209\,
                  I1 =>  \SB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41211\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41211\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41211\,
                   R => '0',
                   S => SYSRESET );

  \=41211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41211\,
                  I0 =>  \ALTEST\,
                  I1 =>  \41212\,
                  I2 =>  '0',
                  I3 => \&41208\ );

  \:41212\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41212\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41212\,
                   R => SYSRESET,
                   S => '0' );

  \=41212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41212\,
                  I0 =>  \41211\,
                  I1 =>  \41210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41213\,
                  I0 =>  \41209\,
                  I1 =>  \41211\,
                  I2 =>  \SB0/\,
                  I3 =>  '0' );

  \:41214\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41214\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41214\,
                   R => '0',
                   S => SYSRESET );

  \=41214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41214\,
                  I0 =>  \41213\,
                  I1 =>  \41215\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41215\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41215\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41215\,
                   R => SYSRESET,
                   S => '0' );

  \=41215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41215\,
                  I0 =>  \41214\,
                  I1 =>  \F08B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FILTIN\   
  \=41216\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41216\,
                  I0 =>  \41214\,
                  I1 =>  \41214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \41218\    
  \=41217\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41217\,
                  I0 =>  \FS01\,
                  I1 =>  \P02\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41218\,
                  I0 =>  \P03/\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 => \&41217\ );

  -- Alias \SYNC4/\   
  \=41219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41219\,
                  I0 =>  \41218\,
                  I1 =>  \41218\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41220\,
                  I0 =>  \CT/\,
                  I1 =>  \P02/\,
                  I2 =>  \P03\,
                  I3 =>  '0' );

  -- Alias \SYNC14/\  
  \=41221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41221\,
                  I0 =>  \41220\,
                  I1 =>  \41220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSCAFL/\  
  \=41222\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41222\,
                  I0 =>  \SCAFAL\,
                  I1 =>  \SCAFAL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWARNF/\  
  \=41223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41223\,
                  I0 =>  \FLTOUT\,
                  I1 =>  \FLTOUT\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41224\,
                  I0 =>  \FLTOUT\,
                  I1 =>  \SCAFAL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41225\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41225\,
                   R => '0',
                   S => SYSRESET );

  \=41225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41225\,
                  I0 =>  \FLTOUT\,
                  I1 =>  \SCAFAL\,
                  I2 =>  \41226\,
                  I3 =>  '0' );

  -- Alias \AGCWAR\   
  \:41226\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41226\,
                   R => SYSRESET,
                   S => '0' );

  \=41226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41226\,
                  I0 =>  \41225\,
                  I1 =>  \CCH33\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WARN\     
  \=41227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41227\,
                  I0 =>  \41224\,
                  I1 =>  \41224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CGCWAR\   
  \=41228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41228\,
                  I0 =>  \WARN\,
                  I1 =>  \WARN\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41229\,
                  I0 =>  \TEMPIN/\,
                  I1 =>  \TMPOUT\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TMPCAU\   
  \=41230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41230\,
                  I0 =>  \41229\,
                  I1 =>  \41229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MOSCAL/\  
  \=41231\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&41231\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41232\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41232\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41232\,
                   R => '0',
                   S => SYSRESET );

  \=41232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41232\,
                  I0 =>  \STRT2\,
                  I1 =>  \41233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OSCALM\   
  \:41233\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41233\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41233\,
                   R => SYSRESET,
                   S => '0' );

  \=41233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41233\,
                  I0 =>  \41232\,
                  I1 =>  \CCH33\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41234\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41234\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41234\,
                   R => '0',
                   S => SYSRESET );

  \=41234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41234\,
                  I0 =>  \SBY\,
                  I1 =>  \41235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41235\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41235\,
                   R => SYSRESET,
                   S => '0' );

  \=41235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41235\,
                  I0 =>  \41234\,
                  I1 =>  \T10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBYEXT\   
  \=41236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41236\,
                  I0 =>  \41234\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41237\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41237\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41237\,
                   R => SYSRESET,
                   S => '0' );

  \=41237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41237\,
                  I0 =>  \GOJAM\,
                  I1 =>  \41238\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41238\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41238\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41238\,
                   R => '0',
                   S => SYSRESET );

  \=41238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41238\,
                  I0 =>  \41237\,
                  I1 =>  \ERRST\,
                  I2 =>  \41236\,
                  I3 =>  '0' );

  \=41239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41239\,
                  I0 =>  \ALTEST\,
                  I1 =>  \41238\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RESTRT\   
  \=41240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41240\,
                  I0 =>  \41239\,
                  I1 =>  \41239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F08B/\    
  \=41241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41241\,
                  I0 =>  \F08B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CON3\     
  \=41242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41242\,
                  I0 =>  \CON2\,
                  I1 =>  \FS10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SCADBL\   
  \=41243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41243\,
                  I0 =>  \CON3\,
                  I1 =>  \2FSFAL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=41245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \41245\,
                  I0 =>  \41204\,
                  I1 =>  \F05A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STRT1\    
  \:41246\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \41246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41246\,
                   R => SYSRESET,
                   S => '0' );

  \=41246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41246\,
                  I0 =>  \41247\,
                  I1 =>  \41245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:41247\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \41247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$41247\,
                   R => '0',
                   S => SYSRESET );

  \=41247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$41247\,
                  I0 =>  \41205\,
                  I1 =>  \41246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *********************************************
  -- ***                                       ***
  -- ***  A14/1 - MEMORY TIMING & ADDRESSING.  ***
  -- ***                                       ***
  -- *********************************************

  -- Alias \ROP/\     
  \=42101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42101\,
                  I0 =>  \S11\,
                  I1 =>  \S11\,
                  I2 =>  '0',
                  I3 => \&42102\ );

  -- Alias \42101\    
  \=42102\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42102\,
                  I0 =>  \S12\,
                  I1 =>  \S12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42103\,
                  I0 =>  \T08/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42104\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42104\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42104\,
                   R => '0',
                   S => SYSRESET );

  \=42104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42104\,
                  I0 =>  \42103\,
                  I1 =>  \42105\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42105\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42105\,
                   R => SYSRESET,
                   S => '0' );

  \=42105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42105\,
                  I0 =>  \42104\,
                  I1 =>  \T09\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=42106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42106\,
                  I0 =>  \42101\,
                  I1 =>  \42104\,
                  I2 =>  \T08\,
                  I3 =>  '0' );

  \:42107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42107\,
                   R => '0',
                   S => SYSRESET );

  \=42107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42107\,
                  I0 =>  \42106\,
                  I1 =>  \42109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IHENV\    
  \=42108\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42108\,
                  I0 =>  \42107\,
                  I1 =>  \42107\,
                  I2 =>  \42107\,
                  I3 =>  '0' );

  \:42109\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42109\,
                   R => SYSRESET,
                   S => '0' );

  \=42109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42109\,
                  I0 =>  \42107\,
                  I1 =>  \42110\,
                  I2 =>  \TIMR\,
                  I3 =>  '0' );

  \=42110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42110\,
                  I0 =>  '0',
                  I1 =>  \T01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42111\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42111\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42111\,
                   R => '0',
                   S => SYSRESET );

  \=42111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42111\,
                  I0 =>  \TIMR\,
                  I1 =>  \42110\,
                  I2 =>  \42112\,
                  I3 =>  '0' );

  \:42112\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42112\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42112\,
                   R => SYSRESET,
                   S => '0' );

  \=42112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42112\,
                  I0 =>  \42111\,
                  I1 =>  \42113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42113\,
                  I0 =>  \PHS4/\,
                  I1 =>  \42101\,
                  I2 =>  \T10/\,
                  I3 =>  '0' );

  \=42114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42114\,
                  I0 =>  \S09\,
                  I1 =>  \42112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42115\,
                  I0 =>  \42112\,
                  I1 =>  \S09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SETAB/\   
  \=42116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42116\,
                  I0 =>  \42114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SETCD/\   
  \=42117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42117\,
                  I0 =>  \42115\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SETAB\    
  \=42118\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42118\,
                  I0 =>  \42116\,
                  I1 =>  \42116\,
                  I2 =>  \42116\,
                  I3 =>  '0' );

  -- Alias \SETCD\    
  \=42119\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42119\,
                  I0 =>  \42117\,
                  I1 =>  \42117\,
                  I2 =>  \42117\,
                  I3 =>  '0' );

  -- Alias \42122\    
  \=42120\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42120\,
                  I0 =>  \42101\,
                  I1 =>  \T06/\,
                  I2 =>  \DV3764\,
                  I3 =>  '0' );

  -- Alias \SBF\      
  \=42121\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42121\,
                  I0 =>  \42123\,
                  I1 =>  \42123\,
                  I2 =>  \42123\,
                  I3 =>  '0' );

  -- Alias \SBFSET\   
  \=42122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42122\,
                  I0 =>  \MNHSBF\,
                  I1 =>  \MP1\,
                  I2 =>  \PHS4/\,
                  I3 => \&42120\ );

  \:42123\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42123\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42123\,
                   R => '0',
                   S => SYSRESET );

  \=42123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42123\,
                  I0 =>  \42124\,
                  I1 =>  \42122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STBF\     
  \:42124\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42124\,
                   R => SYSRESET,
                   S => '0' );

  \=42124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42124\,
                  I0 =>  \GOJAM\,
                  I1 =>  \42125\,
                  I2 =>  \42123\,
                  I3 =>  '0' );

  \=42125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42125\,
                  I0 =>  \T07/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42126\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42126\,
                   R => SYSRESET,
                   S => '0' );

  \=42126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42126\,
                  I0 =>  \42127\,
                  I1 =>  \T08\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \:42127\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42127\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42127\,
                   R => '0',
                   S => SYSRESET );

  \=42127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42127\,
                  I0 =>  \42128\,
                  I1 =>  \42126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42128\,
                  I0 =>  \T05/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42129\,
                  I0 =>  \S09\,
                  I1 =>  \42127\,
                  I2 =>  \S08\,
                  I3 =>  '0' );

  \=42130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42130\,
                  I0 =>  \CLEARA\,
                  I1 =>  \42129\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42131\,
                  I0 =>  \42127\,
                  I1 =>  \S09\,
                  I2 =>  \S08/\,
                  I3 =>  '0' );

  \=42132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42132\,
                  I0 =>  \CLEARB\,
                  I1 =>  \42131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RESETA\   
  \=42133\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42133\,
                  I0 =>  \42130\,
                  I1 =>  \42130\,
                  I2 =>  \42130\,
                  I3 =>  '0' );

  -- Alias \RESETB\   
  \=42134\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42134\,
                  I0 =>  \42132\,
                  I1 =>  \42132\,
                  I2 =>  \42132\,
                  I3 =>  '0' );

  \=42135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42135\,
                  I0 =>  \42127\,
                  I1 =>  \S08\,
                  I2 =>  \S09/\,
                  I3 =>  '0' );

  \=42136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42136\,
                  I0 =>  \CLEARC\,
                  I1 =>  \42135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42137\,
                  I0 =>  \42127\,
                  I1 =>  \S09/\,
                  I2 =>  \S08/\,
                  I3 =>  '0' );

  \=42138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42138\,
                  I0 =>  \42137\,
                  I1 =>  \CLEARD\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RESETC\   
  \=42139\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42139\,
                  I0 =>  \42136\,
                  I1 =>  \42136\,
                  I2 =>  \42136\,
                  I3 =>  '0' );

  -- Alias \RESETD\   
  \=42140\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42140\,
                  I0 =>  \42138\,
                  I1 =>  \42138\,
                  I2 =>  \42138\,
                  I3 =>  '0' );

  -- Alias \42143\    
  \=42141\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42141\,
                  I0 =>  \PHS2/\,
                  I1 =>  \MP1\,
                  I2 =>  '0',
                  I3 => \&42142\ );

  -- Alias \42143\    
  \=42142\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42142\,
                  I0 =>  \GOJ1\,
                  I1 =>  \GOJAM\,
                  I2 =>  \TCSAJ3\,
                  I3 =>  '0' );

  -- Alias \TPGF\     
  \=42143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42143\,
                  I0 =>  \42101\,
                  I1 =>  \T08/\,
                  I2 =>  \DV3764\,
                  I3 => \&42141\ );

  \=42144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42144\,
                  I0 =>  \T02/\,
                  I1 =>  \42101\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42145\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42145\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42145\,
                   R => '0',
                   S => SYSRESET );

  \=42145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42145\,
                  I0 =>  \42144\,
                  I1 =>  \42146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STRGAT\   
  \:42146\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42146\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42146\,
                   R => SYSRESET,
                   S => '0' );

  \=42146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42146\,
                  I0 =>  \42145\,
                  I1 =>  \T08\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=42147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42147\,
                  I0 =>  \42101\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42148\,
                  I0 =>  \T02/\,
                  I1 =>  \42147\,
                  I2 =>  \42155\,
                  I3 =>  '0' );

  -- Alias \42150\    
  \=42149\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42149\,
                  I0 =>  \42148\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42150\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42150\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42150\,
                   R => '0',
                   S => SYSRESET );

  \=42150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42150\,
                  I0 =>  \42148\,
                  I1 =>  \42151\,
                  I2 =>  \42151\,
                  I3 => \&42149\ );

  \:42151\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42151\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42151\,
                   R => SYSRESET,
                   S => '0' );

  \=42151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42151\,
                  I0 =>  \42150\,
                  I1 =>  \T07\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \CLROPE\   
  \=42152\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42152\,
                  I0 =>  \42150\,
                  I1 =>  \42150\,
                  I2 =>  \42150\,
                  I3 =>  '0' );

  \=42154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42154\,
                  I0 =>  \42101\,
                  I1 =>  \T10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42155\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42155\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42155\,
                   R => '0',
                   S => SYSRESET );

  \=42155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42155\,
                  I0 =>  \42154\,
                  I1 =>  \42156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42156\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42156\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42156\,
                   R => SYSRESET,
                   S => '0' );

  \=42156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42156\,
                  I0 =>  \42155\,
                  I1 =>  \T03\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \WHOMPA\   
  \=42157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42157\,
                  I0 =>  '0',
                  I1 =>  \WHOMP/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42201\,
                  I0 =>  \T12/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42202\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42202\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42202\,
                   R => '0',
                   S => SYSRESET );

  \=42202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42202\,
                  I0 =>  \42203\,
                  I1 =>  \42201\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42203\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42203\,
                   R => SYSRESET,
                   S => '0' );

  \=42203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42203\,
                  I0 =>  \T01\,
                  I1 =>  \42202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42204\,
                  I0 =>  \T12A\,
                  I1 =>  \42202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42205\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42205\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42205\,
                   R => SYSRESET,
                   S => '0' );

  \=42205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42205\,
                  I0 =>  \42204\,
                  I1 =>  \TIMR\,
                  I2 =>  \42206\,
                  I3 =>  '0' );

  \:42206\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42206\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42206\,
                   R => '0',
                   S => SYSRESET );

  \=42206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42206\,
                  I0 =>  \42205\,
                  I1 =>  \42211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WEX\      
  \=42207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42207\,
                  I0 =>  \42206\,
                  I1 =>  \42206\,
                  I2 =>  \42206\,
                  I3 =>  '0' );

  -- Alias \WEY\      
  \=42208\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42208\,
                  I0 =>  \42209\,
                  I1 =>  \42209\,
                  I2 =>  \42209\,
                  I3 =>  '0' );

  \:42209\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42209\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42209\,
                   R => '0',
                   S => SYSRESET );

  \=42209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42209\,
                  I0 =>  \42210\,
                  I1 =>  \42214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42210\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42210\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42210\,
                   R => SYSRESET,
                   S => '0' );

  \=42210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42210\,
                  I0 =>  \TIMR\,
                  I1 =>  \42204\,
                  I2 =>  \42209\,
                  I3 =>  '0' );

  \=42211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42211\,
                  I0 =>  \42212\,
                  I1 =>  \T10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42212\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42212\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42212\,
                   R => '0',
                   S => SYSRESET );

  \=42212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42212\,
                  I0 =>  \42213\,
                  I1 =>  \42216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42213\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42213\,
                   R => SYSRESET,
                   S => '0' );

  \=42213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42213\,
                  I0 =>  \TIMR\,
                  I1 =>  \T11\,
                  I2 =>  \42212\,
                  I3 =>  '0' );

  \=42214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42214\,
                  I0 =>  \T10/\,
                  I1 =>  \42225\,
                  I2 =>  \PHS4/\,
                  I3 =>  '0' );

  \=42215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42215\,
                  I0 =>  \PHS4/\,
                  I1 =>  \T02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42216\,
                  I0 =>  \42225\,
                  I1 =>  \T10/\,
                  I2 =>  \PHS3/\,
                  I3 =>  '0' );

  \=42217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42217\,
                  I0 =>  \42225\,
                  I1 =>  \T10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42218\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42218\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42218\,
                   R => SYSRESET,
                   S => '0' );

  \=42218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42218\,
                  I0 =>  \TIMR\,
                  I1 =>  \42215\,
                  I2 =>  \42219\,
                  I3 =>  '0' );

  -- Alias \RSTK/\    
  \:42219\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42219\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42219\,
                   R => '0',
                   S => SYSRESET );

  \=42219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42219\,
                  I0 =>  \42218\,
                  I1 =>  \42216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42220\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42220\,
                   R => SYSRESET,
                   S => '0' );

  \=42220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42220\,
                  I0 =>  \TIMR\,
                  I1 =>  \T01\,
                  I2 =>  \42221\,
                  I3 =>  '0' );

  \:42221\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42221\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42221\,
                   R => '0',
                   S => SYSRESET );

  \=42221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42221\,
                  I0 =>  \42220\,
                  I1 =>  \42217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZID\      
  \=42222\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42222\,
                  I0 =>  \42221\,
                  I1 =>  \42221\,
                  I2 =>  \42221\,
                  I3 => \&42223\ );

  -- Alias \ZID\      
  \=42223\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42223\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  \STRT2\,
                  I3 =>  '0' );

  \=42224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42224\,
                  I0 =>  \T05/\,
                  I1 =>  \42252\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FNERAS/\  
  \:42225\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42225\,
                   R => '0',
                   S => SYSRESET );

  \=42225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42225\,
                  I0 =>  \42224\,
                  I1 =>  \42226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42226\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42226\,
                   R => SYSRESET,
                   S => '0' );

  \=42226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42226\,
                  I0 =>  \42225\,
                  I1 =>  \T12A\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=42227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42227\,
                  I0 =>  \42252\,
                  I1 =>  \T03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42228\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42228\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42228\,
                   R => '0',
                   S => SYSRESET );

  \=42228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42228\,
                  I0 =>  \42227\,
                  I1 =>  \42229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42229\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42229\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42229\,
                   R => SYSRESET,
                   S => '0' );

  \=42229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42229\,
                  I0 =>  \42228\,
                  I1 =>  \42232\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \SETEK\    
  \=42230\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42230\,
                  I0 =>  \42228\,
                  I1 =>  \42228\,
                  I2 =>  \42228\,
                  I3 => \&42231\ );

  -- Alias \SETEK\    
  \=42231\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42231\,
                  I0 =>  \STRT2\,
                  I1 =>  \STRT2\,
                  I2 =>  \STRT2\,
                  I3 =>  '0' );

  \=42232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42232\,
                  I0 =>  \T06/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42233\,
                  I0 =>  \PHS3/\,
                  I1 =>  \42252\,
                  I2 =>  \T03/\,
                  I3 =>  '0' );

  \:42234\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42234\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42234\,
                   R => '0',
                   S => SYSRESET );

  \=42234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42234\,
                  I0 =>  \42233\,
                  I1 =>  \42235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42235\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42235\,
                   R => SYSRESET,
                   S => '0' );

  \=42235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42235\,
                  I0 =>  \42234\,
                  I1 =>  \GOJAM\,
                  I2 =>  \42241\,
                  I3 =>  '0' );

  -- Alias \REY\      
  \=42236\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42236\,
                  I0 =>  \42234\,
                  I1 =>  \42234\,
                  I2 =>  \42234\,
                  I3 =>  '0' );

  -- Alias \REX\      
  \=42237\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42237\,
                  I0 =>  \42238\,
                  I1 =>  \42238\,
                  I2 =>  \42238\,
                  I3 =>  '0' );

  \:42238\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42238\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42238\,
                   R => '0',
                   S => SYSRESET );

  \=42238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42238\,
                  I0 =>  \42240\,
                  I1 =>  \42239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42239\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42239\,
                   R => SYSRESET,
                   S => '0' );

  \=42239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42239\,
                  I0 =>  \42238\,
                  I1 =>  \42241\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=42240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42240\,
                  I0 =>  \42252\,
                  I1 =>  \T03/\,
                  I2 =>  \PHS4/\,
                  I3 =>  '0' );

  -- Alias \REDRST\   
  \=42241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42241\,
                  I0 =>  \42242\,
                  I1 =>  \T05\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42242\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42242\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42242\,
                   R => '0',
                   S => SYSRESET );

  \=42242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42242\,
                  I0 =>  \42244\,
                  I1 =>  \42243\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:42243\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42243\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42243\,
                   R => SYSRESET,
                   S => '0' );

  \=42243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42243\,
                  I0 =>  \42242\,
                  I1 =>  \T06\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42244\,
                  I0 =>  \T05/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBESET\   
  \=42245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42245\,
                  I0 =>  \T04/\,
                  I1 =>  \42252\,
                  I2 =>  \SCAD\,
                  I3 =>  '0' );

  \:42246\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \42246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42246\,
                   R => '0',
                   S => SYSRESET );

  \=42246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42246\,
                  I0 =>  \42247\,
                  I1 =>  \42245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STBE\     
  \:42247\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \42247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$42247\,
                   R => SYSRESET,
                   S => '0' );

  \=42247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$42247\,
                  I0 =>  \GOJAM\,
                  I1 =>  \T05\,
                  I2 =>  \42246\,
                  I3 =>  '0' );

  -- Alias \TPGE\     
  \=42248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42248\,
                  I0 =>  \SCAD\,
                  I1 =>  \42252\,
                  I2 =>  \GOJAM\,
                  I3 => \&42250\ );

  -- Alias \TPARG/\   
  \=42249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42249\,
                  I0 =>  \TPGF\,
                  I1 =>  \42248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \42248\    
  \=42250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42250\,
                  I0 =>  \T05/\,
                  I1 =>  \PHS3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBE\      
  \=42251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42251\,
                  I0 =>  \42246\,
                  I1 =>  \42246\,
                  I2 =>  \42246\,
                  I3 =>  '0' );

  -- Alias \ERAS/\    
  \=42252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42252\,
                  I0 =>  \42254\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ERAS\     
  \=42254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42254\,
                  I0 =>  \TCSAJ3\,
                  I1 =>  \S11\,
                  I2 =>  \S12\,
                  I3 => \&42255\ );

  -- Alias \42254\    
  \=42255\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42255\,
                  I0 =>  \INOUT\,
                  I1 =>  \CHINC\,
                  I2 =>  \GOJ1\,
                  I3 => \&42256\ );

  -- Alias \ERAS\     
  \=42256\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42256\,
                  I0 =>  \MP1\,
                  I1 =>  \MAMU\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOTEST/\  
  \=42257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42257\,
                  I0 =>  \PSEUDO\,
                  I1 =>  \NISQL/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *********************************************
  -- ***                                       ***
  -- ***  A14/2 - MEMORY TIMING & ADDRESSING.  ***
  -- ***                                       ***
  -- *********************************************

  -- Alias \XB0\      
  \=42301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42301\,
                  I0 =>  \S01\,
                  I1 =>  \S02\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- Alias \XB0/\     
  \=42302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42302\,
                  I0 =>  \42301\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB0E\     
  \=42306\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42306\,
                  I0 =>  \42302\,
                  I1 =>  \42302\,
                  I2 =>  \42302\,
                  I3 =>  '0' );

  -- Alias \XB1\      
  \=42307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42307\,
                  I0 =>  \S01/\,
                  I1 =>  \S02\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- Alias \XB1/\     
  \=42308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42308\,
                  I0 =>  \42307\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB1E\     
  \=42311\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42311\,
                  I0 =>  \42308\,
                  I1 =>  \42308\,
                  I2 =>  \42308\,
                  I3 =>  '0' );

  -- Alias \XB2\      
  \=42312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42312\,
                  I0 =>  \S01\,
                  I1 =>  \S02/\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- Alias \XB2/\     
  \=42313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42313\,
                  I0 =>  \42312\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB2E\     
  \=42316\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42316\,
                  I0 =>  \42313\,
                  I1 =>  \42313\,
                  I2 =>  \42313\,
                  I3 =>  '0' );

  -- Alias \XB3\      
  \=42317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42317\,
                  I0 =>  \S01/\,
                  I1 =>  \S02/\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- Alias \XB3/\     
  \=42318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42318\,
                  I0 =>  \42317\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB3E\     
  \=42321\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42321\,
                  I0 =>  \42318\,
                  I1 =>  \42318\,
                  I2 =>  \42318\,
                  I3 =>  '0' );

  -- Alias \XB4\      
  \=42322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42322\,
                  I0 =>  \S01\,
                  I1 =>  \S02\,
                  I2 =>  \S03/\,
                  I3 =>  '0' );

  -- Alias \XB4/\     
  \=42323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42323\,
                  I0 =>  \42322\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB4E\     
  \=42326\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42326\,
                  I0 =>  \42323\,
                  I1 =>  \42323\,
                  I2 =>  \42323\,
                  I3 =>  '0' );

  -- Alias \XB5\      
  \=42327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42327\,
                  I0 =>  \S01/\,
                  I1 =>  \S02\,
                  I2 =>  \S03/\,
                  I3 =>  '0' );

  -- Alias \XB5/\     
  \=42328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42328\,
                  I0 =>  \42327\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB5E\     
  \=42331\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42331\,
                  I0 =>  \42328\,
                  I1 =>  \42328\,
                  I2 =>  \42328\,
                  I3 =>  '0' );

  -- Alias \XB6\      
  \=42332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42332\,
                  I0 =>  \S02/\,
                  I1 =>  \S03/\,
                  I2 =>  \S01\,
                  I3 =>  '0' );

  -- Alias \XB6/\     
  \=42333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42333\,
                  I0 =>  \42332\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB6E\     
  \=42336\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42336\,
                  I0 =>  \42333\,
                  I1 =>  \42333\,
                  I2 =>  \42333\,
                  I3 =>  '0' );

  -- Alias \XB7\      
  \=42337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42337\,
                  I0 =>  \S02/\,
                  I1 =>  \S03/\,
                  I2 =>  \S01/\,
                  I3 =>  '0' );

  -- Alias \XB7/\     
  \=42339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42339\,
                  I0 =>  \42337\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XB7E\     
  \=42341\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42341\,
                  I0 =>  \42339\,
                  I1 =>  \42339\,
                  I2 =>  \42339\,
                  I3 =>  '0' );

  -- Alias \YB0\      
  \=42342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42342\,
                  I0 =>  \S07\,
                  I1 =>  \S08\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB0/\     
  \=42343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42343\,
                  I0 =>  \42342\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB0E\     
  \=42345\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42345\,
                  I0 =>  \42343\,
                  I1 =>  \42343\,
                  I2 =>  \42343\,
                  I3 =>  '0' );

  -- Alias \YB1\      
  \=42346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42346\,
                  I0 =>  \S08\,
                  I1 =>  \S07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB1/\     
  \=42347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42347\,
                  I0 =>  \42346\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB1E\     
  \=42348\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42348\,
                  I0 =>  \42347\,
                  I1 =>  \42347\,
                  I2 =>  \42347\,
                  I3 =>  '0' );

  -- Alias \YB2\      
  \=42349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42349\,
                  I0 =>  \S07\,
                  I1 =>  \S08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB2/\     
  \=42350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42350\,
                  I0 =>  \42349\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB2E\     
  \=42351\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42351\,
                  I0 =>  \42350\,
                  I1 =>  \42350\,
                  I2 =>  \42350\,
                  I3 =>  '0' );

  -- Alias \YB3\      
  \=42352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42352\,
                  I0 =>  \S07/\,
                  I1 =>  \S08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB3/\     
  \=42353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42353\,
                  I0 =>  \42352\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \YB3E\     
  \=42354\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42354\,
                  I0 =>  \42353\,
                  I1 =>  \42353\,
                  I2 =>  \42353\,
                  I3 =>  '0' );

  -- Alias \RILP1\    
  \=42355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42355\,
                  I0 =>  \42342\,
                  I1 =>  \42352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RILP1/\   
  \=42356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42356\,
                  I0 =>  \42355\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CXB1/\    
  \=42357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42357\,
                  I0 =>  \XB1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT0\      
  \=42401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42401\,
                  I0 =>  \S06\,
                  I1 =>  \S05\,
                  I2 =>  \S04\,
                  I3 =>  '0' );

  -- Alias \XT0/\     
  \=42402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42402\,
                  I0 =>  \42401\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT0E\     
  \=42404\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42404\,
                  I0 =>  \42402\,
                  I1 =>  \42402\,
                  I2 =>  \42402\,
                  I3 =>  '0' );

  -- Alias \XT1\      
  \=42405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42405\,
                  I0 =>  \S06\,
                  I1 =>  \S05\,
                  I2 =>  \S04/\,
                  I3 =>  '0' );

  -- Alias \XT1/\     
  \=42406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42406\,
                  I0 =>  \42405\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT1E\     
  \=42408\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42408\,
                  I0 =>  \42406\,
                  I1 =>  \42406\,
                  I2 =>  \42406\,
                  I3 =>  '0' );

  -- Alias \XT2\      
  \=42409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42409\,
                  I0 =>  \S06\,
                  I1 =>  \S05/\,
                  I2 =>  \S04\,
                  I3 =>  '0' );

  -- Alias \XT2/\     
  \=42410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42410\,
                  I0 =>  \42409\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT2E\     
  \=42412\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42412\,
                  I0 =>  \42410\,
                  I1 =>  \42410\,
                  I2 =>  \42410\,
                  I3 =>  '0' );

  -- Alias \XT3\      
  \=42413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42413\,
                  I0 =>  \S06\,
                  I1 =>  \S05/\,
                  I2 =>  \S04/\,
                  I3 =>  '0' );

  -- Alias \XT3/\     
  \=42414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42414\,
                  I0 =>  \42413\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT3E\     
  \=42416\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42416\,
                  I0 =>  \42414\,
                  I1 =>  \42414\,
                  I2 =>  \42414\,
                  I3 =>  '0' );

  -- Alias \XT4\      
  \=42417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42417\,
                  I0 =>  \S06/\,
                  I1 =>  \S05\,
                  I2 =>  \S04\,
                  I3 =>  '0' );

  -- Alias \XT4/\     
  \=42418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42418\,
                  I0 =>  \42417\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT4E\     
  \=42420\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42420\,
                  I0 =>  \42418\,
                  I1 =>  \42418\,
                  I2 =>  \42418\,
                  I3 =>  '0' );

  -- Alias \XT5\      
  \=42421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42421\,
                  I0 =>  \S06/\,
                  I1 =>  \S05\,
                  I2 =>  \S04/\,
                  I3 =>  '0' );

  -- Alias \XT5/\     
  \=42423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42423\,
                  I0 =>  \42421\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT5E\     
  \=42424\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42424\,
                  I0 =>  \42423\,
                  I1 =>  \42423\,
                  I2 =>  \42423\,
                  I3 =>  '0' );

  -- Alias \XT6\      
  \=42425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42425\,
                  I0 =>  \S06/\,
                  I1 =>  \S05/\,
                  I2 =>  \S04\,
                  I3 =>  '0' );

  -- Alias \RB1\      
  \=42426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42426\,
                  I0 =>  \RB1/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT6/\     
  \=42427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42427\,
                  I0 =>  \42425\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT6E\     
  \=42428\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42428\,
                  I0 =>  \42427\,
                  I1 =>  \42427\,
                  I2 =>  \42427\,
                  I3 =>  '0' );

  -- Alias \XT7\      
  \=42429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42429\,
                  I0 =>  \S06/\,
                  I1 =>  \S05/\,
                  I2 =>  \S04/\,
                  I3 =>  '0' );

  -- Alias \XT7/\     
  \=42431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42431\,
                  I0 =>  \42429\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XT7E\     
  \=42432\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42432\,
                  I0 =>  \42431\,
                  I1 =>  \42431\,
                  I2 =>  \42431\,
                  I3 =>  '0' );

  \=42433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42433\,
                  I0 =>  \42401\,
                  I1 =>  \42413\,
                  I2 =>  '0',
                  I3 => \&42434\ );

  -- Alias \42433\    
  \=42434\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42434\,
                  I0 =>  \42421\,
                  I1 =>  \42425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42435\,
                  I0 =>  \42433\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42436\,
                  I0 =>  \42440\,
                  I1 =>  \RILP1\,
                  I2 =>  \42433\,
                  I3 =>  '0' );

  \=42437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42437\,
                  I0 =>  \42442\,
                  I1 =>  \RILP1\,
                  I2 =>  \42435\,
                  I3 =>  '0' );

  \=42438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42438\,
                  I0 =>  \42442\,
                  I1 =>  \RILP1/\,
                  I2 =>  \42433\,
                  I3 =>  '0' );

  \=42439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42439\,
                  I0 =>  \42435\,
                  I1 =>  \RILP1/\,
                  I2 =>  \42440\,
                  I3 =>  '0' );

  \=42440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42440\,
                  I0 =>  \XB0\,
                  I1 =>  \XB3\,
                  I2 =>  '0',
                  I3 => \&42441\ );

  -- Alias \42440\    
  \=42441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42441\,
                  I0 =>  \XB5\,
                  I1 =>  \XB6\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42442\,
                  I0 =>  \42440\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42443\,
                  I0 =>  \42436\,
                  I1 =>  \42437\,
                  I2 =>  '0',
                  I3 => \&42444\ );

  -- Alias \42443\    
  \=42444\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42444\,
                  I0 =>  \42438\,
                  I1 =>  \42439\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42445\,
                  I0 =>  \42443\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ILP\      
  \=42446\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42446\,
                  I0 =>  \42445\,
                  I1 =>  \42445\,
                  I2 =>  \42445\,
                  I3 =>  '0' );

  -- Alias \ILP/\     
  \=42447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42447\,
                  I0 =>  \42443\,
                  I1 =>  \42443\,
                  I2 =>  \42443\,
                  I3 =>  '0' );

  \=42448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42448\,
                  I0 =>  \RSC/\,
                  I1 =>  \RT/\,
                  I2 =>  \SCAD/\,
                  I3 =>  '0' );

  -- Alias \RSCG/\    
  \=42449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42449\,
                  I0 =>  \42448\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=42451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42451\,
                  I0 =>  \WSC/\,
                  I1 =>  '0',
                  I2 =>  \SCAD/\,
                  I3 =>  '0' );

  -- Alias \WSCG/\    
  \=42452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42452\,
                  I0 =>  \42451\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \R1C\      
  \=42454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42454\,
                  I0 =>  \R1C/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBYREL/\  
  \=42457\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&42457\,
                  I0 =>  \SBY\,
                  I1 =>  \SBY\,
                  I2 =>  \SBY\,
                  I3 =>  '0' );

  -- Alias \NOTEST\   
  \=42459\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \42459\,
                  I0 =>  '0',
                  I1 =>  \NOTEST/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *******************************
  -- ***                         ***
  -- ***  A15/1 - RUPT SERVICE.  ***
  -- ***                         ***
  -- *******************************

  \=35101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35101\,
                  I0 =>  \WL16/\,
                  I1 =>  \WFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FB16/\    
  \:35102\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35102\,
                   R => '0',
                   S => SYSRESET );

  \=35102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35102\,
                  I0 =>  \35101\,
                  I1 =>  \35151\,
                  I2 =>  \35104\,
                  I3 =>  '0' );

  -- Alias \FB16\     
  \:35104\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35104\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35104\,
                   R => SYSRESET,
                   S => '0' );

  \=35104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35104\,
                  I0 =>  \35102\,
                  I1 =>  \CFBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BK16\     
  \=35105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35105\,
                  I0 =>  \35102\,
                  I1 =>  \RFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL16/\    
  \=35106\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35106\,
                  I0 =>  \35105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35107\,
                  I0 =>  \WL14/\,
                  I1 =>  \WFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FB14/\    
  \:35108\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35108\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35108\,
                   R => '0',
                   S => SYSRESET );

  \=35108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35108\,
                  I0 =>  \35107\,
                  I1 =>  \35152\,
                  I2 =>  \35110\,
                  I3 =>  '0' );

  -- Alias \FB14\     
  \:35110\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35110\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35110\,
                   R => SYSRESET,
                   S => '0' );

  \=35110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35110\,
                  I0 =>  \35108\,
                  I1 =>  \CFBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35111\,
                  I0 =>  \35108\,
                  I1 =>  \RFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35113\,
                  I0 =>  \WL13/\,
                  I1 =>  \WFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FB13/\    
  \:35114\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35114\,
                   R => '0',
                   S => SYSRESET );

  \=35114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35114\,
                  I0 =>  \35113\,
                  I1 =>  \35153\,
                  I2 =>  \35115\,
                  I3 =>  '0' );

  -- Alias \FB13\     
  \:35115\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35115\,
                   R => SYSRESET,
                   S => '0' );

  \=35115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35115\,
                  I0 =>  \35114\,
                  I1 =>  \CFBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35116\,
                  I0 =>  \35114\,
                  I1 =>  \RFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL13/\    
  \=35117\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35117\,
                  I0 =>  \35116\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35118\,
                  I0 =>  \WL12/\,
                  I1 =>  \WFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FB12/\    
  \:35119\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35119\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35119\,
                   R => '0',
                   S => SYSRESET );

  \=35119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35119\,
                  I0 =>  \35118\,
                  I1 =>  \35154\,
                  I2 =>  \35120\,
                  I3 =>  '0' );

  -- Alias \FB12\     
  \:35120\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35120\,
                   R => SYSRESET,
                   S => '0' );

  \=35120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35120\,
                  I0 =>  \35119\,
                  I1 =>  \CFBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35121\,
                  I0 =>  \35119\,
                  I1 =>  \RFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL12/\    
  \=35122\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35122\,
                  I0 =>  \RSTRT\,
                  I1 =>  \35121\,
                  I2 =>  \RPTA12\,
                  I3 =>  '0' );

  \=35123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35123\,
                  I0 =>  \WFBG/\,
                  I1 =>  \WL11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FB11/\    
  \:35124\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35124\,
                   R => '0',
                   S => SYSRESET );

  \=35124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35124\,
                  I0 =>  \35123\,
                  I1 =>  \35155\,
                  I2 =>  \35125\,
                  I3 =>  '0' );

  -- Alias \FB11\     
  \:35125\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35125\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35125\,
                   R => SYSRESET,
                   S => '0' );

  \=35125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35125\,
                  I0 =>  \35124\,
                  I1 =>  \CFBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35126\,
                  I0 =>  \35124\,
                  I1 =>  \RFBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL11/\    
  \=35127\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35127\,
                  I0 =>  \35126\,
                  I1 =>  \35132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35128\,
                  I0 =>  \WL11/\,
                  I1 =>  \WEBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35129\,
                  I0 =>  \WL03/\,
                  I1 =>  \WBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EB11/\    
  \:35130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35130\,
                   R => '0',
                   S => SYSRESET );

  \=35130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35130\,
                  I0 =>  \35128\,
                  I1 =>  \35129\,
                  I2 =>  \35131\,
                  I3 => \&35150\ );

  -- Alias \EB11\     
  \:35131\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35131\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35131\,
                   R => SYSRESET,
                   S => '0' );

  \=35131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35131\,
                  I0 =>  \35130\,
                  I1 =>  \CEBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35132\,
                  I0 =>  \REBG/\,
                  I1 =>  \35130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BBK3\     
  \=35133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35133\,
                  I0 =>  \35130\,
                  I1 =>  \RBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35137\    
  \=35134\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35134\,
                  I0 =>  \35157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35135\,
                  I0 =>  \WL10/\,
                  I1 =>  \WEBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35136\,
                  I0 =>  \WL02/\,
                  I1 =>  \WBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EB10/\    
  \:35137\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35137\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35137\,
                   R => '0',
                   S => SYSRESET );

  \=35137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35137\,
                  I0 =>  \35135\,
                  I1 =>  \35136\,
                  I2 =>  \35138\,
                  I3 => \&35134\ );

  -- Alias \EB10\     
  \:35138\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35138\,
                   R => SYSRESET,
                   S => '0' );

  \=35138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35138\,
                  I0 =>  \35137\,
                  I1 =>  \CEBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35139\,
                  I0 =>  \REBG/\,
                  I1 =>  \35137\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BBK2\     
  \=35140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35140\,
                  I0 =>  \35137\,
                  I1 =>  \RBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL10/\    
  \=35141\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35141\,
                  I0 =>  \35139\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35145\    
  \=35142\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35142\,
                  I0 =>  \35158\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35143\,
                  I0 =>  \WL09/\,
                  I1 =>  \WEBG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35144\,
                  I0 =>  \WL01/\,
                  I1 =>  \WBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EB9/\     
  \:35145\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35145\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35145\,
                   R => '0',
                   S => SYSRESET );

  \=35145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35145\,
                  I0 =>  \35143\,
                  I1 =>  \35144\,
                  I2 =>  \35146\,
                  I3 => \&35142\ );

  -- Alias \EB9\      
  \:35146\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35146\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35146\,
                   R => SYSRESET,
                   S => '0' );

  \=35146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35146\,
                  I0 =>  \35145\,
                  I1 =>  \CEBG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35147\,
                  I0 =>  \REBG/\,
                  I1 =>  \35145\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BBK1\     
  \=35148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35148\,
                  I0 =>  \35145\,
                  I1 =>  \RBBEG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL09/\    
  \=35149\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35149\,
                  I0 =>  \35147\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35130\    
  \=35150\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35150\,
                  I0 =>  \35156\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35151\,
                  I0 =>  \SUMA16/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB16/\,
                  I3 =>  '0' );

  \=35152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35152\,
                  I0 =>  \SUMA14/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB14/\,
                  I3 =>  '0' );

  \=35153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35153\,
                  I0 =>  \SUMA13/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB13/\,
                  I3 =>  '0' );

  \=35154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35154\,
                  I0 =>  \SUMA12/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB12/\,
                  I3 =>  '0' );

  \=35155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35155\,
                  I0 =>  \SUMA11/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB11/\,
                  I3 =>  '0' );

  \=35156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35156\,
                  I0 =>  \SUMA03/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB03/\,
                  I3 =>  '0' );

  \=35157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35157\,
                  I0 =>  \SUMA02/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB02/\,
                  I3 =>  '0' );

  \=35158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35158\,
                  I0 =>  \SUMA01/\,
                  I1 =>  \U2BBKG/\,
                  I2 =>  \SUMB01/\,
                  I3 =>  '0' );

  \=35201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35201\,
                  I0 =>  \S12/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35203\,
                  I0 =>  \35124\,
                  I1 =>  \35201\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35204\,
                  I0 =>  \S11/\,
                  I1 =>  \S12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F11/\     
  \=35205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35205\,
                  I0 =>  \35203\,
                  I1 =>  \35204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F11\      
  \=35206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35206\,
                  I0 =>  \35205\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F13\      
  \=35207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35207\,
                  I0 =>  \35201\,
                  I1 =>  \35114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F12/\     
  \=35208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35208\,
                  I0 =>  \35201\,
                  I1 =>  \35120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F12\      
  \=35209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35209\,
                  I0 =>  \35208\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F13/\     
  \=35210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35210\,
                  I0 =>  \35207\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35211\,
                  I0 =>  \E5\,
                  I1 =>  \35102\,
                  I2 =>  \E7/\,
                  I3 =>  '0' );

  \=35212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35212\,
                  I0 =>  \E7/\,
                  I1 =>  \35108\,
                  I2 =>  \E6\,
                  I3 =>  '0' );

  -- Alias \F16\      
  \=35213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35213\,
                  I0 =>  \35108\,
                  I1 =>  \35102\,
                  I2 =>  \E7/\,
                  I3 => \&35214\ );

  -- Alias \35213\    
  \=35214\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35214\,
                  I0 =>  \35201\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F14\      
  \=35215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35215\,
                  I0 =>  \35201\,
                  I1 =>  \35211\,
                  I2 =>  \35108\,
                  I3 =>  '0' );

  -- Alias \F15\      
  \=35216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35216\,
                  I0 =>  \35102\,
                  I1 =>  \35212\,
                  I2 =>  \35201\,
                  I3 =>  '0' );

  -- Alias \F14/\     
  \=35217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35217\,
                  I0 =>  \35215\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F15/\     
  \=35218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35218\,
                  I0 =>  \35216\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F16/\     
  \=35219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35219\,
                  I0 =>  \35213\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35220\,
                  I0 =>  \XB4/\,
                  I1 =>  \XT4/\,
                  I2 =>  \KRPTA/\,
                  I3 =>  '0' );

  \=35221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35221\,
                  I0 =>  \KRPTA/\,
                  I1 =>  \XB0/\,
                  I2 =>  \XT5/\,
                  I3 =>  '0' );

  \:35222\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35222\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35222\,
                   R => '0',
                   S => SYSRESET );

  \=35222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35222\,
                  I0 =>  \RADRPT\,
                  I1 =>  \35223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35223\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35223\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35223\,
                   R => SYSRESET,
                   S => '0' );

  \=35223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35223\,
                  I0 =>  \35222\,
                  I1 =>  \35220\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \:35224\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35224\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35224\,
                   R => '0',
                   S => SYSRESET );

  \=35224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35224\,
                  I0 =>  \HNDRPT\,
                  I1 =>  \35225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35225\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35225\,
                   R => SYSRESET,
                   S => '0' );

  \=35225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35225\,
                  I0 =>  \35224\,
                  I1 =>  \35221\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \PRPOR3\   
  \=35226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35226\,
                  I0 =>  \PRPOR1\,
                  I1 =>  \35222\,
                  I2 =>  \DNRPTA\,
                  I3 =>  '0' );

  -- Alias \PRPOR4\   
  \=35227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35227\,
                  I0 =>  \PRPOR1\,
                  I1 =>  \DNRPTA\,
                  I2 =>  '0',
                  I3 => \&35228\ );

  -- Alias \35227\    
  \=35228\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35228\,
                  I0 =>  \35223\,
                  I1 =>  \35224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35229\,
                  I0 =>  \35225\,
                  I1 =>  \35223\,
                  I2 =>  '0',
                  I3 => \&35230\ );

  -- Alias \35229\    
  \=35230\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35230\,
                  I0 =>  \PRPOR1\,
                  I1 =>  \DNRPTA\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35231\,
                  I0 =>  \PRPOR2\,
                  I1 =>  \35226\,
                  I2 =>  \35227\,
                  I3 =>  '0' );

  -- Alias \RPTAD6\   
  \=35232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35232\,
                  I0 =>  \35231\,
                  I1 =>  \RRPA1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RPTA12\   
  \=35233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35233\,
                  I0 =>  \RRPA1/\,
                  I1 =>  \35229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35234\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35234\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35234\,
                   R => SYSRESET,
                   S => '0' );

  \=35234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35234\,
                  I0 =>  \35229\,
                  I1 =>  \35235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RUPTOR/\  
  \:35235\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35235\,
                   R => '0',
                   S => SYSRESET );

  \=35235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35235\,
                  I0 =>  \35234\,
                  I1 =>  \T10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35236\,
                  I0 =>  \C37M\,
                  I1 =>  \C40M\,
                  I2 =>  \C41M\,
                  I3 => \&35237\ );

  -- Alias \35236\    
  \=35237\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35237\,
                  I0 =>  \C42M\,
                  I1 =>  \C43M\,
                  I2 =>  \C44M\,
                  I3 =>  '0' );

  \=35238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35238\,
                  I0 =>  \INCSET/\,
                  I1 =>  \35236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MINC/\    
  \:35239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35239\,
                   R => '0',
                   S => SYSRESET );

  \=35239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35239\,
                  I0 =>  \35238\,
                  I1 =>  \35240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MINC\     
  \:35240\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35240\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35240\,
                   R => SYSRESET,
                   S => '0' );

  \=35240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35240\,
                  I0 =>  \35239\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35241\,
                  I0 =>  \C32P\,
                  I1 =>  \C33P\,
                  I2 =>  \C34P\,
                  I3 => \&35242\ );

  -- Alias \35241\    
  \=35242\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35242\,
                  I0 =>  \C35P\,
                  I1 =>  \C36P\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35243\,
                  I0 =>  \INCSET/\,
                  I1 =>  \35241\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PCDU/\    
  \:35244\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35244\,
                   R => '0',
                   S => SYSRESET );

  \=35244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35244\,
                  I0 =>  \35243\,
                  I1 =>  \35245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PCDU\     
  \:35245\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35245\,
                   R => SYSRESET,
                   S => '0' );

  \=35245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35245\,
                  I0 =>  \35244\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35246\,
                  I0 =>  \C32M\,
                  I1 =>  \C33M\,
                  I2 =>  \C34M\,
                  I3 => \&35247\ );

  -- Alias \35246\    
  \=35247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35247\,
                  I0 =>  \C35M\,
                  I1 =>  \C36M\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35248\,
                  I0 =>  \INCSET/\,
                  I1 =>  \35246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MCDU/\    
  \:35249\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35249\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35249\,
                   R => '0',
                   S => SYSRESET );

  \=35249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35249\,
                  I0 =>  \35248\,
                  I1 =>  \35250\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MCDU\     
  \:35250\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35250\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35250\,
                   R => SYSRESET,
                   S => '0' );

  \=35250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35250\,
                  I0 =>  \35249\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL14/\    
  \=35251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35251\,
                  I0 =>  \35111\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *******************************
  -- ***                         ***
  -- ***  A15/2 - RUPT SERVICE.  ***
  -- ***                         ***
  -- *******************************

  -- Alias \WOVR/\    
  \=35301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35301\,
                  I0 =>  \WOVR\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35302\,
                  I0 =>  \35301\,
                  I1 =>  \OVF/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35303\,
                  I0 =>  \35302\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \KRPTA/\   
  \=35304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35304\,
                  I0 =>  \KRPT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35306\,
                  I0 =>  \XT0/\,
                  I1 =>  \XB4/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  -- Alias \T6RPT\    
  \=35307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35307\,
                  I0 =>  \CA3/\,
                  I1 =>  \XB1/\,
                  I2 =>  \ZOUT/\,
                  I3 =>  '0' );

  \:35308\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35308\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35308\,
                   R => '0',
                   S => SYSRESET );

  \=35308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35308\,
                  I0 =>  \35307\,
                  I1 =>  \35309\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35309\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35309\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35309\,
                   R => SYSRESET,
                   S => '0' );

  \=35309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35309\,
                  I0 =>  \35308\,
                  I1 =>  \GOJAM\,
                  I2 =>  \35306\,
                  I3 =>  '0' );

  \=35310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35310\,
                  I0 =>  \XB0/\,
                  I1 =>  \XT1/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \=35311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35311\,
                  I0 =>  \CA3/\,
                  I1 =>  \XB0/\,
                  I2 =>  \35303\,
                  I3 =>  '0' );

  \:35312\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35312\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35312\,
                   R => '0',
                   S => SYSRESET );

  \=35312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35312\,
                  I0 =>  \35311\,
                  I1 =>  \35313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35313\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35313\,
                   R => SYSRESET,
                   S => '0' );

  \=35313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35313\,
                  I0 =>  \35312\,
                  I1 =>  \35310\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=35314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35314\,
                  I0 =>  \35309\,
                  I1 =>  \35312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35315\,
                  I0 =>  \XT1/\,
                  I1 =>  \XB4/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \=35316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35316\,
                  I0 =>  \CA2/\,
                  I1 =>  \XB6/\,
                  I2 =>  \35303\,
                  I3 =>  '0' );

  \:35317\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35317\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35317\,
                   R => '0',
                   S => SYSRESET );

  \=35317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35317\,
                  I0 =>  \35316\,
                  I1 =>  \35318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35318\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35318\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35318\,
                   R => SYSRESET,
                   S => '0' );

  \=35318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35318\,
                  I0 =>  \35317\,
                  I1 =>  \35315\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=35319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35319\,
                  I0 =>  \35309\,
                  I1 =>  \35317\,
                  I2 =>  \35313\,
                  I3 =>  '0' );

  \=35320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35320\,
                  I0 =>  \35309\,
                  I1 =>  \35318\,
                  I2 =>  \35313\,
                  I3 =>  '0' );

  \=35321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35321\,
                  I0 =>  \35320\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35322\,
                  I0 =>  \CA2/\,
                  I1 =>  \XB7/\,
                  I2 =>  \35303\,
                  I3 =>  '0' );

  \:35323\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35323\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35323\,
                   R => '0',
                   S => SYSRESET );

  \=35323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35323\,
                  I0 =>  \35322\,
                  I1 =>  \35326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35324\,
                  I0 =>  \35321\,
                  I1 =>  \35323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35325\,
                  I0 =>  \XT2/\,
                  I1 =>  \XB0/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \:35326\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35326\,
                   R => SYSRESET,
                   S => '0' );

  \=35326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35326\,
                  I0 =>  \35323\,
                  I1 =>  \35325\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \KY1RST\   
  \=35327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35327\,
                  I0 =>  \XB4/\,
                  I1 =>  \XT2/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \:35328\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35328\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35328\,
                   R => '0',
                   S => SYSRESET );

  \=35328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35328\,
                  I0 =>  \KYRPT1\,
                  I1 =>  \35329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35329\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35329\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35329\,
                   R => SYSRESET,
                   S => '0' );

  \=35329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35329\,
                  I0 =>  \35328\,
                  I1 =>  \35327\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=35330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35330\,
                  I0 =>  \35321\,
                  I1 =>  \35328\,
                  I2 =>  \35326\,
                  I3 =>  '0' );

  \=35331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35331\,
                  I0 =>  \35321\,
                  I1 =>  \35329\,
                  I2 =>  \35326\,
                  I3 =>  '0' );

  \=35332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35332\,
                  I0 =>  \35331\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \KY2RST\   
  \=35333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35333\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB0/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \:35334\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35334\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35334\,
                   R => '0',
                   S => SYSRESET );

  \=35334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35334\,
                  I0 =>  \KYRPT2\,
                  I1 =>  \MKRPT\,
                  I2 =>  \35335\,
                  I3 =>  '0' );

  \:35335\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35335\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35335\,
                   R => SYSRESET,
                   S => '0' );

  \=35335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35335\,
                  I0 =>  \35334\,
                  I1 =>  \35333\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=35336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35336\,
                  I0 =>  \35332\,
                  I1 =>  \35334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35339\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB4/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \:35340\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35340\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35340\,
                   R => '0',
                   S => SYSRESET );

  \=35340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35340\,
                  I0 =>  \UPRUPT\,
                  I1 =>  \35341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:35341\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35341\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35341\,
                   R => SYSRESET,
                   S => '0' );

  \=35341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35341\,
                  I0 =>  \35340\,
                  I1 =>  \35339\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=35342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35342\,
                  I0 =>  \35332\,
                  I1 =>  \35340\,
                  I2 =>  \35335\,
                  I3 =>  '0' );

  \=35343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35343\,
                  I0 =>  \35332\,
                  I1 =>  \35341\,
                  I2 =>  \35335\,
                  I3 =>  '0' );

  -- Alias \PRPOR1\   
  \=35344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35344\,
                  I0 =>  \35343\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DRPRST\   
  \=35345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35345\,
                  I0 =>  \XB0/\,
                  I1 =>  \XT4/\,
                  I2 =>  \35304\,
                  I3 =>  '0' );

  \:35346\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \35346\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35346\,
                   R => '0',
                   S => SYSRESET );

  \=35346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35346\,
                  I0 =>  \DLKPLS\,
                  I1 =>  \35347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DNRPTA\   
  \:35347\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \35347\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$35347\,
                   R => SYSRESET,
                   S => '0' );

  \=35347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$35347\,
                  I0 =>  \35346\,
                  I1 =>  \35345\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \PRPOR2\   
  \=35348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35348\,
                  I0 =>  \35344\,
                  I1 =>  \35346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RRPA1/\   
  \=35349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35349\,
                  I0 =>  \RRPA\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35351\    
  \=35350\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35350\,
                  I0 =>  \35309\,
                  I1 =>  \35319\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35351\,
                  I0 =>  \35330\,
                  I1 =>  \35342\,
                  I2 =>  \PRPOR3\,
                  I3 => \&35350\ );

  -- Alias \RPTAD3\   
  \=35352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35352\,
                  I0 =>  \35349\,
                  I1 =>  \35351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35354\    
  \=35353\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35353\,
                  I0 =>  \35314\,
                  I1 =>  \35319\,
                  I2 =>  \35336\,
                  I3 =>  '0' );

  \=35354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35354\,
                  I0 =>  \35342\,
                  I1 =>  \PRPOR4\,
                  I2 =>  '0',
                  I3 => \&35353\ );

  -- Alias \RPTAD4\   
  \=35355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35355\,
                  I0 =>  \35349\,
                  I1 =>  \35354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \35357\    
  \=35356\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35356\,
                  I0 =>  \35330\,
                  I1 =>  \35324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35357\,
                  I0 =>  \35336\,
                  I1 =>  \35342\,
                  I2 =>  '0',
                  I3 => \&35356\ );

  -- Alias \RPTAD5\   
  \=35358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35358\,
                  I0 =>  \35349\,
                  I1 =>  \35357\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RL03/\    
  \=35359\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35359\,
                  I0 =>  \RPTAD3\,
                  I1 =>  \BBK3\,
                  I2 =>  \CAD3\,
                  I3 =>  '0' );

  -- Alias \RL02/\    
  \=35360\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35360\,
                  I0 =>  \CAD2\,
                  I1 =>  \BBK2\,
                  I2 =>  \R6\,
                  I3 =>  '0' );

  \=35401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35401\,
                  I0 =>  \STRGAT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR412\   
  \=35403\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35403\,
                  I0 =>  \35401\,
                  I1 =>  \35408\,
                  I2 =>  \35408\,
                  I3 => \&35404\ );

  -- Alias \STR412\   
  \=35404\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35404\,
                  I0 =>  \35401\,
                  I1 =>  \35405\,
                  I2 =>  \35405\,
                  I3 =>  '0' );

  \=35405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35405\,
                  I0 =>  \F11\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR311\   
  \=35406\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35406\,
                  I0 =>  \35401\,
                  I1 =>  \35414\,
                  I2 =>  \35414\,
                  I3 => \&35407\ );

  -- Alias \STR311\   
  \=35407\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35407\,
                  I0 =>  \35401\,
                  I1 =>  \35405\,
                  I2 =>  \35405\,
                  I3 =>  '0' );

  \=35408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35408\,
                  I0 =>  \S10\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR210\   
  \=35409\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35409\,
                  I0 =>  \35401\,
                  I1 =>  \35408\,
                  I2 =>  \35408\,
                  I3 => \&35410\ );

  -- Alias \STR210\   
  \=35410\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35410\,
                  I0 =>  \35401\,
                  I1 =>  \35411\,
                  I2 =>  \35411\,
                  I3 =>  '0' );

  \=35411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35411\,
                  I0 =>  \F11/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR19\    
  \=35412\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35412\,
                  I0 =>  \35401\,
                  I1 =>  \35414\,
                  I2 =>  \35414\,
                  I3 => \&35413\ );

  -- Alias \STR19\    
  \=35413\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35413\,
                  I0 =>  \35401\,
                  I1 =>  \35411\,
                  I2 =>  \35411\,
                  I3 =>  '0' );

  \=35414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35414\,
                  I0 =>  \S10/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35415\,
                  I0 =>  \F16\,
                  I1 =>  \F15\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35416\,
                  I0 =>  \35415\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35417\,
                  I0 =>  \35416\,
                  I1 =>  \35423\,
                  I2 =>  \35430\,
                  I3 =>  '0' );

  \=35418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35418\,
                  I0 =>  \35417\,
                  I1 =>  \35432\,
                  I2 =>  \35445\,
                  I3 =>  '0' );

  \=35419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35419\,
                  I0 =>  \35418\,
                  I1 =>  \F12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35420\,
                  I0 =>  \35419\,
                  I1 =>  \35427\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR14\    
  \=35421\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35421\,
                  I0 =>  \35420\,
                  I1 =>  \35420\,
                  I2 =>  \35420\,
                  I3 =>  '0' );

  -- Alias \ROPER\    
  \=35422\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35422\,
                  I0 =>  \35426\,
                  I1 =>  \35426\,
                  I2 =>  \35426\,
                  I3 =>  '0' );

  \=35423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35423\,
                  I0 =>  \F14/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35424\,
                  I0 =>  \35416\,
                  I1 =>  \35423\,
                  I2 =>  \35431\,
                  I3 =>  '0' );

  \=35425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35425\,
                  I0 =>  \35416\,
                  I1 =>  \35437\,
                  I2 =>  \35430\,
                  I3 =>  '0' );

  \=35426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35426\,
                  I0 =>  \35417\,
                  I1 =>  \35424\,
                  I2 =>  \35425\,
                  I3 =>  '0' );

  \=35427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35427\,
                  I0 =>  \35433\,
                  I1 =>  \F12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35428\,
                  I0 =>  \35419\,
                  I1 =>  \35447\,
                  I2 =>  \35440\,
                  I3 =>  '0' );

  -- Alias \LOMOD\    
  \=35429\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35429\,
                  I0 =>  \35428\,
                  I1 =>  \35428\,
                  I2 =>  \35428\,
                  I3 =>  '0' );

  \=35430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35430\,
                  I0 =>  \F13/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35431\,
                  I0 =>  \F13\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35432\,
                  I0 =>  \35416\,
                  I1 =>  \35437\,
                  I2 =>  \35431\,
                  I3 =>  '0' );

  \=35433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35433\,
                  I0 =>  \35424\,
                  I1 =>  \35438\,
                  I2 =>  \35452\,
                  I3 =>  '0' );

  \=35434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35434\,
                  I0 =>  \35446\,
                  I1 =>  \F12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35435\,
                  I0 =>  \35434\,
                  I1 =>  \35440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR58\    
  \=35436\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35436\,
                  I0 =>  \35435\,
                  I1 =>  \35435\,
                  I2 =>  \35435\,
                  I3 =>  '0' );

  \=35437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35437\,
                  I0 =>  \F14\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35438\,
                  I0 =>  \35443\,
                  I1 =>  \35423\,
                  I2 =>  \35430\,
                  I3 =>  '0' );

  \=35439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35439\,
                  I0 =>  \35438\,
                  I1 =>  \35432\,
                  I2 =>  \35444\,
                  I3 =>  '0' );

  \=35440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35440\,
                  I0 =>  \35418\,
                  I1 =>  \F12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ROPES\    
  \=35441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35441\,
                  I0 =>  \35439\,
                  I1 =>  \35439\,
                  I2 =>  \35439\,
                  I3 =>  '0' );

  \=35442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35442\,
                  I0 =>  \F16\,
                  I1 =>  \F15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35443\,
                  I0 =>  \35442\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35444\,
                  I0 =>  \35443\,
                  I1 =>  \35423\,
                  I2 =>  \35431\,
                  I3 =>  '0' );

  \=35445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35445\,
                  I0 =>  \35443\,
                  I1 =>  \35437\,
                  I2 =>  \35430\,
                  I3 =>  '0' );

  \=35446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35446\,
                  I0 =>  \35425\,
                  I1 =>  \35444\,
                  I2 =>  \35453\,
                  I3 =>  '0' );

  \=35447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35447\,
                  I0 =>  \35433\,
                  I1 =>  \F12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35448\,
                  I0 =>  \35427\,
                  I1 =>  \35455\,
                  I2 =>  \35434\,
                  I3 =>  '0' );

  -- Alias \HIMOD\    
  \=35449\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35449\,
                  I0 =>  \35448\,
                  I1 =>  \35448\,
                  I2 =>  \35448\,
                  I3 =>  '0' );

  \=35450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35450\,
                  I0 =>  \F15\,
                  I1 =>  \F16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35451\,
                  I0 =>  \35450\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35452\,
                  I0 =>  \35443\,
                  I1 =>  \35437\,
                  I2 =>  \35431\,
                  I3 =>  '0' );

  \=35453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35453\,
                  I0 =>  \35451\,
                  I1 =>  \35423\,
                  I2 =>  \35430\,
                  I3 =>  '0' );

  \=35454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35454\,
                  I0 =>  \35445\,
                  I1 =>  \35452\,
                  I2 =>  \35453\,
                  I3 =>  '0' );

  \=35455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35455\,
                  I0 =>  \35446\,
                  I1 =>  \F12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=35456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \35456\,
                  I0 =>  \35447\,
                  I1 =>  \35455\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STR912\   
  \=35457\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35457\,
                  I0 =>  \35456\,
                  I1 =>  \35456\,
                  I2 =>  \35456\,
                  I3 =>  '0' );

  -- Alias \ROPET\    
  \=35458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35458\,
                  I0 =>  \35454\,
                  I1 =>  \35454\,
                  I2 =>  \35454\,
                  I3 =>  '0' );

  -- Alias \RL01/\    
  \=35460\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&35460\,
                  I0 =>  \CAD1\,
                  I1 =>  \BBK1\,
                  I2 =>  \RB1F\,
                  I3 =>  '0' );

  -- **************************
  -- ***                    ***
  -- ***  A16/1 - INOUT I.  ***
  -- ***                    ***
  -- **************************

  \=43101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43101\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43102\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43102\,
                   R => '0',
                   S => SYSRESET );

  \=43102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43102\,
                  I0 =>  \43101\,
                  I1 =>  \43103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43103\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43103\,
                   R => SYSRESET,
                   S => '0' );

  \=43103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43103\,
                  I0 =>  \43102\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43104\,
                  I0 =>  \43217\,
                  I1 =>  \43102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+X+P\   
  \=43105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43105\,
                  I0 =>  \43102\,
                  I1 =>  \43102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR01/\  
  \=43106\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43106\,
                  I0 =>  \43258\,
                  I1 =>  \43104\,
                  I2 =>  \CH3201\,
                  I3 => \&43407\ );

  \=43107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43107\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43108\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43108\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43108\,
                   R => '0',
                   S => SYSRESET );

  \=43108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43108\,
                  I0 =>  \43107\,
                  I1 =>  \43109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43109\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43109\,
                   R => SYSRESET,
                   S => '0' );

  \=43109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43109\,
                  I0 =>  \43108\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43110\,
                  I0 =>  \43217\,
                  I1 =>  \43108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-X-P\   
  \=43111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43111\,
                  I0 =>  \43108\,
                  I1 =>  \43108\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR02/\  
  \=43112\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43112\,
                  I0 =>  \43253\,
                  I1 =>  \43110\,
                  I2 =>  \CH3202\,
                  I3 => \&43408\ );

  \=43113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43113\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43114\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43114\,
                   R => '0',
                   S => SYSRESET );

  \=43114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43114\,
                  I0 =>  \43113\,
                  I1 =>  \43115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43115\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43115\,
                   R => SYSRESET,
                   S => '0' );

  \=43115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43115\,
                  I0 =>  \43114\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43116\,
                  I0 =>  \43217\,
                  I1 =>  \43114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-X+P\   
  \=43117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43117\,
                  I0 =>  \43114\,
                  I1 =>  \43114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR03/\  
  \=43118\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43118\,
                  I0 =>  \43248\,
                  I1 =>  \43116\,
                  I2 =>  \CH3203\,
                  I3 => \&43419\ );

  \=43119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43119\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43120\,
                   R => '0',
                   S => SYSRESET );

  \=43120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43120\,
                  I0 =>  \43119\,
                  I1 =>  \43121\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43121\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43121\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43121\,
                   R => SYSRESET,
                   S => '0' );

  \=43121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43121\,
                  I0 =>  \43120\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43122\,
                  I0 =>  \43217\,
                  I1 =>  \43120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+X-P\   
  \=43123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43123\,
                  I0 =>  \43120\,
                  I1 =>  \43120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR04/\  
  \=43124\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43124\,
                  I0 =>  \43243\,
                  I1 =>  \43122\,
                  I2 =>  \CH3204\,
                  I3 => \&43420\ );

  \=43125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43125\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43126\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43126\,
                   R => '0',
                   S => SYSRESET );

  \=43126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43126\,
                  I0 =>  \43125\,
                  I1 =>  \43127\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43127\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43127\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43127\,
                   R => SYSRESET,
                   S => '0' );

  \=43127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43127\,
                  I0 =>  \43126\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43128\,
                  I0 =>  \43217\,
                  I1 =>  \43126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+X+Y\   
  \=43129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43129\,
                  I0 =>  \43126\,
                  I1 =>  \43126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR05/\  
  \=43130\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43130\,
                  I0 =>  \43238\,
                  I1 =>  \43128\,
                  I2 =>  \CH3205\,
                  I3 => \&43425\ );

  \=43131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43131\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43132\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43132\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43132\,
                   R => '0',
                   S => SYSRESET );

  \=43132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43132\,
                  I0 =>  \43131\,
                  I1 =>  \43133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43133\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43133\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43133\,
                   R => SYSRESET,
                   S => '0' );

  \=43133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43133\,
                  I0 =>  \43132\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43134\,
                  I0 =>  \43217\,
                  I1 =>  \43132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-X-Y\   
  \=43135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43135\,
                  I0 =>  \43132\,
                  I1 =>  \43132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR06/\  
  \=43136\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43136\,
                  I0 =>  \43233\,
                  I1 =>  \43134\,
                  I2 =>  \CH3206\,
                  I3 => \&43437\ );

  \=43137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43137\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43138\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43138\,
                   R => '0',
                   S => SYSRESET );

  \=43138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43138\,
                  I0 =>  \43137\,
                  I1 =>  \43139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43139\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43139\,
                   R => SYSRESET,
                   S => '0' );

  \=43139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43139\,
                  I0 =>  \43138\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43140\,
                  I0 =>  \43217\,
                  I1 =>  \43138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-X+Y\   
  \=43141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43141\,
                  I0 =>  \43138\,
                  I1 =>  \43138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR07/\  
  \=43142\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43142\,
                  I0 =>  \43222\,
                  I1 =>  \43140\,
                  I2 =>  \CH3207\,
                  I3 => \&43439\ );

  \=43143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43143\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \43149\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43144\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43144\,
                   R => '0',
                   S => SYSRESET );

  \=43144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43144\,
                  I0 =>  \43143\,
                  I1 =>  \43145\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43145\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43145\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43145\,
                   R => SYSRESET,
                   S => '0' );

  \=43145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43145\,
                  I0 =>  \43144\,
                  I1 =>  \43154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43146\,
                  I0 =>  \43217\,
                  I1 =>  \43144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+X-Y\   
  \=43147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43147\,
                  I0 =>  \43144\,
                  I1 =>  \43144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR08/\  
  \=43148\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43148\,
                  I0 =>  \43204\,
                  I1 =>  \43146\,
                  I2 =>  \CH3208\,
                  I3 => \&44348\ );

  -- Alias \WCH05/\   
  \=43149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43149\,
                  I0 =>  \43151\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43151\,
                  I0 =>  \XB5/\,
                  I1 =>  \XT0/\,
                  I2 =>  \WCHG/\,
                  I3 =>  '0' );

  \=43152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43152\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XB5/\,
                  I2 =>  \XT0/\,
                  I3 =>  '0' );

  \=43153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43153\,
                  I0 =>  \43152\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH05\    
  \=43154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43154\,
                  I0 =>  \43153\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43156\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \WCH12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43157\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43157\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43157\,
                   R => '0',
                   S => SYSRESET );

  \=43157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43157\,
                  I0 =>  \43156\,
                  I1 =>  \43158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43158\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43158\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43158\,
                   R => SYSRESET,
                   S => '0' );

  \=43158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43158\,
                  I0 =>  \43157\,
                  I1 =>  \CCH12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1208\   
  \=43159\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43159\,
                  I0 =>  \RCH12/\,
                  I1 =>  \43157\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TVCNAB\   
  \=43160\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43160\,
                  I0 =>  \43157\,
                  I1 =>  \43157\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43201\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43202\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43202\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43202\,
                   R => '0',
                   S => SYSRESET );

  \=43202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43202\,
                  I0 =>  \43201\,
                  I1 =>  \43203\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43203\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43203\,
                   R => SYSRESET,
                   S => '0' );

  \=43203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43203\,
                  I0 =>  \43202\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43204\,
                  I0 =>  \43214\,
                  I1 =>  \43202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+Y-R\   
  \=43205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43205\,
                  I0 =>  \43202\,
                  I1 =>  \43202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43206\,
                  I0 =>  \XB6/\,
                  I1 =>  \WCHG/\,
                  I2 =>  \XT0/\,
                  I3 =>  '0' );

  -- Alias \WCH06/\   
  \=43207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43207\,
                  I0 =>  \43206\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43209\,
                  I0 =>  \XT0/\,
                  I1 =>  \CCHG/\,
                  I2 =>  \XB6/\,
                  I3 =>  '0' );

  \=43210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43210\,
                  I0 =>  \GOJAM\,
                  I1 =>  \43209\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH06\    
  \=43211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43211\,
                  I0 =>  \43210\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43213\,
                  I0 =>  \XB6/\,
                  I1 =>  \XT0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH06/\   
  \=43214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43214\,
                  I0 =>  \43213\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43216\,
                  I0 =>  \XT0/\,
                  I1 =>  \XB5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH05/\   
  \=43217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43217\,
                  I0 =>  \43216\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43219\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43220\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43220\,
                   R => '0',
                   S => SYSRESET );

  \=43220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43220\,
                  I0 =>  \43219\,
                  I1 =>  \43221\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43221\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43221\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43221\,
                   R => SYSRESET,
                   S => '0' );

  \=43221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43221\,
                  I0 =>  \43220\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43222\,
                  I0 =>  \43214\,
                  I1 =>  \43220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-Y+R\   
  \=43223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43223\,
                  I0 =>  \43220\,
                  I1 =>  \43220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43224\,
                  I0 =>  \WCH12/\,
                  I1 =>  \CHWL07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43225\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43225\,
                   R => '0',
                   S => SYSRESET );

  \=43225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43225\,
                  I0 =>  \43224\,
                  I1 =>  \43226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43226\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43226\,
                   R => SYSRESET,
                   S => '0' );

  \=43226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43226\,
                  I0 =>  \43225\,
                  I1 =>  \CCH12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1207\   
  \=43227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43227\,
                  I0 =>  \RCH12/\,
                  I1 =>  \43225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1207\   
  \=43228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43228\,
                  I0 =>  \43225\,
                  I1 =>  \43225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1207/\  
  \=43229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43229\,
                  I0 =>  \43226\,
                  I1 =>  \43226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43230\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43231\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43231\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43231\,
                   R => '0',
                   S => SYSRESET );

  \=43231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43231\,
                  I0 =>  \43230\,
                  I1 =>  \43232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43232\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43232\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43232\,
                   R => SYSRESET,
                   S => '0' );

  \=43232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43232\,
                  I0 =>  \43231\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43233\,
                  I0 =>  \43214\,
                  I1 =>  \43231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-Y-R\   
  \=43234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43234\,
                  I0 =>  \43231\,
                  I1 =>  \43231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43235\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43236\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43236\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43236\,
                   R => '0',
                   S => SYSRESET );

  \=43236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43236\,
                  I0 =>  \43235\,
                  I1 =>  \43237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43237\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43237\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43237\,
                   R => SYSRESET,
                   S => '0' );

  \=43237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43237\,
                  I0 =>  \43236\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43238\,
                  I0 =>  \43214\,
                  I1 =>  \43236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+Y+R\   
  \=43239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43239\,
                  I0 =>  \43236\,
                  I1 =>  \43236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43240\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43241\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43241\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43241\,
                   R => '0',
                   S => SYSRESET );

  \=43241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43241\,
                  I0 =>  \43240\,
                  I1 =>  \43242\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43242\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43242\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43242\,
                   R => SYSRESET,
                   S => '0' );

  \=43242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43242\,
                  I0 =>  \43241\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43243\,
                  I0 =>  \43214\,
                  I1 =>  \43241\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+Z-R\   
  \=43244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43244\,
                  I0 =>  \43241\,
                  I1 =>  \43241\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43245\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43246\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43246\,
                   R => '0',
                   S => SYSRESET );

  \=43246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43246\,
                  I0 =>  \43245\,
                  I1 =>  \43247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43247\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43247\,
                   R => SYSRESET,
                   S => '0' );

  \=43247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43247\,
                  I0 =>  \43246\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43248\,
                  I0 =>  \43214\,
                  I1 =>  \43246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-Z+R\   
  \=43249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43249\,
                  I0 =>  \43246\,
                  I1 =>  \43246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43250\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43251\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43251\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43251\,
                   R => '0',
                   S => SYSRESET );

  \=43251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43251\,
                  I0 =>  \43250\,
                  I1 =>  \43252\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43252\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43252\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43252\,
                   R => SYSRESET,
                   S => '0' );

  \=43252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43252\,
                  I0 =>  \43251\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43253\,
                  I0 =>  \43214\,
                  I1 =>  \43251\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC-Z-R\   
  \=43254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43254\,
                  I0 =>  \43251\,
                  I1 =>  \43251\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43255\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \43207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43256\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43256\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43256\,
                   R => '0',
                   S => SYSRESET );

  \=43256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43256\,
                  I0 =>  \43255\,
                  I1 =>  \43257\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43257\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43257\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43257\,
                   R => SYSRESET,
                   S => '0' );

  \=43257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43257\,
                  I0 =>  \43256\,
                  I1 =>  \43211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43258\,
                  I0 =>  \43214\,
                  I1 =>  \43256\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RC+Z+R\   
  \=43259\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43259\,
                  I0 =>  \43256\,
                  I1 =>  \43256\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- **************************
  -- ***                    ***
  -- ***  A16/2 - INOUT I.  ***
  -- ***                    ***
  -- **************************

  \=43301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43301\,
                  I0 =>  \43356\,
                  I1 =>  \43303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZOPCDU\   
  \=43302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43302\,
                  I0 =>  \43303\,
                  I1 =>  \43303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43303\,
                   R => '0',
                   S => SYSRESET );

  \=43303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43303\,
                  I0 =>  \43305\,
                  I1 =>  \43304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43304\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43304\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43304\,
                   R => SYSRESET,
                   S => '0' );

  \=43304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43304\,
                  I0 =>  \43303\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43305\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43306\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43307\,
                   R => '0',
                   S => SYSRESET );

  \=43307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43307\,
                  I0 =>  \43306\,
                  I1 =>  \43308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43308\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43308\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43308\,
                   R => SYSRESET,
                   S => '0' );

  \=43308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43308\,
                  I0 =>  \43307\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43309\,
                  I0 =>  \43356\,
                  I1 =>  \43307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ENEROP\   
  \=43310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43310\,
                  I0 =>  \43307\,
                  I1 =>  \43307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43311\,
                  I0 =>  \43356\,
                  I1 =>  \43313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STARON\   
  \=43312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43312\,
                  I0 =>  \43313\,
                  I1 =>  \43313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43313\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43313\,
                   R => '0',
                   S => SYSRESET );

  \=43313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43313\,
                  I0 =>  \43315\,
                  I1 =>  \43314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43314\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43314\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43314\,
                   R => SYSRESET,
                   S => '0' );

  \=43314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43314\,
                  I0 =>  \43313\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43315\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43316\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43317\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43317\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43317\,
                   R => '0',
                   S => SYSRESET );

  \=43317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43317\,
                  I0 =>  \43316\,
                  I1 =>  \43318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43318\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43318\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43318\,
                   R => SYSRESET,
                   S => '0' );

  \=43318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43318\,
                  I0 =>  \43317\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43319\,
                  I0 =>  \43356\,
                  I1 =>  \43317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \COARSE\   
  \=43320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43320\,
                  I0 =>  \43317\,
                  I1 =>  \43317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43321\,
                  I0 =>  \43356\,
                  I1 =>  \43323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZIMCDU\   
  \=43322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43322\,
                  I0 =>  \43323\,
                  I1 =>  \43323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43323\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43323\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43323\,
                   R => '0',
                   S => SYSRESET );

  \=43323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43323\,
                  I0 =>  \43325\,
                  I1 =>  \43324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43324\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43324\,
                   R => SYSRESET,
                   S => '0' );

  \=43324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43324\,
                  I0 =>  \43323\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43325\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43326\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43327\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43327\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43327\,
                   R => '0',
                   S => SYSRESET );

  \=43327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43327\,
                  I0 =>  \43326\,
                  I1 =>  \43328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43328\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43328\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43328\,
                   R => SYSRESET,
                   S => '0' );

  \=43328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43328\,
                  I0 =>  \43327\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43329\,
                  I0 =>  \43356\,
                  I1 =>  \43327\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ENERIM\   
  \=43330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43330\,
                  I0 =>  \43327\,
                  I1 =>  \43327\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1209\   
  \=43331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43331\,
                  I0 =>  \43356\,
                  I1 =>  \43333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S4BTAK\   
  \=43332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43332\,
                  I0 =>  \43333\,
                  I1 =>  \43333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43333\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43333\,
                   R => '0',
                   S => SYSRESET );

  \=43333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43333\,
                  I0 =>  \43335\,
                  I1 =>  \43334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43334\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43334\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43334\,
                   R => SYSRESET,
                   S => '0' );

  \=43334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43334\,
                  I0 =>  \43333\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43335\,
                  I0 =>  \CHWL09/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43336\,
                  I0 =>  \CHWL10/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43337\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43337\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43337\,
                   R => '0',
                   S => SYSRESET );

  \=43337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43337\,
                  I0 =>  \43336\,
                  I1 =>  \43338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43338\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43338\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43338\,
                   R => SYSRESET,
                   S => '0' );

  \=43338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43338\,
                  I0 =>  \43337\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1210\   
  \=43339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43339\,
                  I0 =>  \43356\,
                  I1 =>  \43337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZEROPT\   
  \=43340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43340\,
                  I0 =>  \43337\,
                  I1 =>  \43337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1211\   
  \=43341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43341\,
                  I0 =>  \43356\,
                  I1 =>  \43343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DISDAC\   
  \=43342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43342\,
                  I0 =>  \43343\,
                  I1 =>  \43343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43343\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43343\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43343\,
                   R => '0',
                   S => SYSRESET );

  \=43343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43343\,
                  I0 =>  \43345\,
                  I1 =>  \43344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43344\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43344\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43344\,
                   R => SYSRESET,
                   S => '0' );

  \=43344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43344\,
                  I0 =>  \43343\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43345\,
                  I0 =>  \CHWL11/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WCH12/\   
  \=43346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43346\,
                  I0 =>  \43349\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43349\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XB2/\,
                  I2 =>  \XT1/\,
                  I3 =>  '0' );

  \=43350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43350\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XT1/\,
                  I2 =>  \XB2/\,
                  I3 =>  '0' );

  \=43351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43351\,
                  I0 =>  \43350\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH12\    
  \=43352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43352\,
                  I0 =>  \43351\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43355\,
                  I0 =>  \XT1/\,
                  I1 =>  \XB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH12/\   
  \=43356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43356\,
                  I0 =>  \43355\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ISSWAR\   
  \=43401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43401\,
                  I0 =>  \43404\,
                  I1 =>  \43404\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43402\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43404\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43403\,
                   R => SYSRESET,
                   S => '0' );

  \=43403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43403\,
                  I0 =>  \43404\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43404\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43404\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43404\,
                   R => '0',
                   S => SYSRESET );

  \=43404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43404\,
                  I0 =>  \43405\,
                  I1 =>  \43403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43405\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43406\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR01/\  
  \=43407\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43407\,
                  I0 =>  \43301\,
                  I1 =>  \43402\,
                  I2 =>  \CH1501\,
                  I3 => \&44306\ );

  -- Alias \CHOR02/\  
  \=43408\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43408\,
                  I0 =>  \43309\,
                  I1 =>  \43411\,
                  I2 =>  \CH1502\,
                  I3 => \&44312\ );

  \:43409\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43409\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43409\,
                   R => '0',
                   S => SYSRESET );

  \=43409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43409\,
                  I0 =>  \43406\,
                  I1 =>  \43410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43410\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43410\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43410\,
                   R => SYSRESET,
                   S => '0' );

  \=43410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43410\,
                  I0 =>  \43409\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43411\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43409\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \COMACT\   
  \=43412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43412\,
                  I0 =>  \43409\,
                  I1 =>  \43409\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \UPLACT\   
  \=43413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43413\,
                  I0 =>  \43416\,
                  I1 =>  \43416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43414\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43415\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43415\,
                   R => SYSRESET,
                   S => '0' );

  \=43415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43415\,
                  I0 =>  \43416\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43416\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43416\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43416\,
                   R => '0',
                   S => SYSRESET );

  \=43416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43416\,
                  I0 =>  \43417\,
                  I1 =>  \43415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43417\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43418\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR03/\  
  \=43419\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43419\,
                  I0 =>  \43311\,
                  I1 =>  \43414\,
                  I2 =>  \CH1503\,
                  I3 => \&44318\ );

  -- Alias \CHOR04/\  
  \=43420\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43420\,
                  I0 =>  \43319\,
                  I1 =>  \43423\,
                  I2 =>  \CH1504\,
                  I3 => \&44324\ );

  \:43421\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43421\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43421\,
                   R => '0',
                   S => SYSRESET );

  \=43421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43421\,
                  I0 =>  \43418\,
                  I1 =>  \43422\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43422\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43422\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43422\,
                   R => SYSRESET,
                   S => '0' );

  \=43422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43422\,
                  I0 =>  \43421\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43423\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43421\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TMPOUT\   
  \=43424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43424\,
                  I0 =>  \43421\,
                  I1 =>  \43421\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR05/\  
  \=43425\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43425\,
                  I0 =>  \43321\,
                  I1 =>  \43428\,
                  I2 =>  \CH0705\,
                  I3 => \&44330\ );

  -- Alias \43427\    
  \=43426\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43426\,
                  I0 =>  \FLASH\,
                  I1 =>  \FLASH\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \KYRLS\    
  \=43427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43427\,
                  I0 =>  \43430\,
                  I1 =>  \43430\,
                  I2 =>  '0',
                  I3 => \&43426\ );

  \=43428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43428\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43429\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43429\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43429\,
                   R => SYSRESET,
                   S => '0' );

  \=43429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43429\,
                  I0 =>  \43430\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43430\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43430\,
                   R => '0',
                   S => SYSRESET );

  \=43430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43430\,
                  I0 =>  \43431\,
                  I1 =>  \43429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43431\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43432\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43433\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43433\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43433\,
                   R => SYSRESET,
                   S => '0' );

  \=43433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43433\,
                  I0 =>  \43434\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43434\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43434\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43434\,
                   R => '0',
                   S => SYSRESET );

  \=43434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43434\,
                  I0 =>  \43432\,
                  I1 =>  \43433\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \VNFLSH\   
  \=43435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43435\,
                  I0 =>  \43434\,
                  I1 =>  \43434\,
                  I2 =>  '0',
                  I3 => \&43438\ );

  \=43436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43436\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43434\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR06/\  
  \=43437\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43437\,
                  I0 =>  \43329\,
                  I1 =>  \43436\,
                  I2 =>  \CH0706\,
                  I3 => \&44336\ );

  -- Alias \43435\    
  \=43438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43438\,
                  I0 =>  \FLASH/\,
                  I1 =>  \FLASH/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR07/\  
  \=43439\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43439\,
                  I0 =>  \CH1207\,
                  I1 =>  \43442\,
                  I2 =>  \CH0707\,
                  I3 => \&44342\ );

  -- Alias \43441\    
  \=43440\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&43440\,
                  I0 =>  \FLASH\,
                  I1 =>  \FLASH\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OPEROR\   
  \=43441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43441\,
                  I0 =>  \43444\,
                  I1 =>  \43444\,
                  I2 =>  '0',
                  I3 => \&43440\ );

  \=43442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43442\,
                  I0 =>  \RCH11/\,
                  I1 =>  \43444\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43443\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43443\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43443\,
                   R => SYSRESET,
                   S => '0' );

  \=43443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43443\,
                  I0 =>  \43444\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43444\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43444\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43444\,
                   R => '0',
                   S => SYSRESET );

  \=43444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43444\,
                  I0 =>  \43445\,
                  I1 =>  \43443\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43445\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43446\,
                  I0 =>  \CHWL12/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43447\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43447\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43447\,
                   R => '0',
                   S => SYSRESET );

  \=43447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43447\,
                  I0 =>  \43446\,
                  I1 =>  \43448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43448\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43448\,
                   R => SYSRESET,
                   S => '0' );

  \=43448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43448\,
                  I0 =>  \43447\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1212\   
  \=43449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43449\,
                  I0 =>  \43356\,
                  I1 =>  \43447\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MROLGT\   
  \=43450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43450\,
                  I0 =>  \43447\,
                  I1 =>  \43447\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S4BSEQ\   
  \=43451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43451\,
                  I0 =>  \43454\,
                  I1 =>  \43454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1213\   
  \=43452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43452\,
                  I0 =>  \43356\,
                  I1 =>  \43454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43453\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43453\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43453\,
                   R => SYSRESET,
                   S => '0' );

  \=43453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43453\,
                  I0 =>  \43454\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43454\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43454\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43454\,
                   R => '0',
                   S => SYSRESET );

  \=43454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43454\,
                  I0 =>  \43455\,
                  I1 =>  \43453\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43455\,
                  I0 =>  \CHWL13/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=43456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43456\,
                  I0 =>  \CHWL14/\,
                  I1 =>  \43346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43457\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \43457\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43457\,
                   R => '0',
                   S => SYSRESET );

  \=43457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43457\,
                  I0 =>  \43456\,
                  I1 =>  \43458\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:43458\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \43458\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$43458\,
                   R => SYSRESET,
                   S => '0' );

  \=43458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$43458\,
                  I0 =>  \43457\,
                  I1 =>  \43352\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1214\   
  \=43459\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43459\,
                  I0 =>  \43356\,
                  I1 =>  \43457\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \S4BOFF\   
  \=43460\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \43460\,
                  I0 =>  \43457\,
                  I1 =>  \43457\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ***************************
  -- ***                     ***
  -- ***  A17/1 - INOUT II.  ***
  -- ***                     ***
  -- ***************************

  \=44101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44101\,
                  I0 =>  \ULLTHR\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44102\,
                  I0 =>  \IN3301\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR01/\  
  \=44103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44103\,
                  I0 =>  \44102\,
                  I1 =>  \44101\,
                  I2 =>  \44201\,
                  I3 => \&43106\ );

  \=44104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44104\,
                  I0 =>  \SMSEPR\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44105\,
                  I0 =>  \RRPONA\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR02/\  
  \=44106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44106\,
                  I0 =>  \44105\,
                  I1 =>  \44104\,
                  I2 =>  \44202\,
                  I3 => \&43112\ );

  \=44107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44107\,
                  I0 =>  \SPSRDY\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44108\,
                  I0 =>  \RRRLSC\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR03/\  
  \=44109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44109\,
                  I0 =>  \44108\,
                  I1 =>  \44107\,
                  I2 =>  \44203\,
                  I3 => \&43118\ );

  \=44110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44110\,
                  I0 =>  \S4BSAB\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44111\,
                  I0 =>  \ZEROP\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR04/\  
  \=44112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44112\,
                  I0 =>  \44111\,
                  I1 =>  \44110\,
                  I2 =>  \44204\,
                  I3 => \&43124\ );

  \=44113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44113\,
                  I0 =>  \LFTOFF\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44114\,
                  I0 =>  \OPMSW2\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR05/\  
  \=44115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44115\,
                  I0 =>  \44114\,
                  I1 =>  \44113\,
                  I2 =>  \44205\,
                  I3 => \&43130\ );

  \=44116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44116\,
                  I0 =>  \GUIREL\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44117\,
                  I0 =>  \OPMSW3\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR06/\  
  \=44118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44118\,
                  I0 =>  \44117\,
                  I1 =>  \44116\,
                  I2 =>  \44215\,
                  I3 => \&43136\ );

  \=44119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44119\,
                  I0 =>  \OPCDFL\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44120\,
                  I0 =>  \STRPRS\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR07/\  
  \=44121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44121\,
                  I0 =>  \44120\,
                  I1 =>  \44119\,
                  I2 =>  \44216\,
                  I3 => \&43142\ );

  \=44122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44122\,
                  I0 =>  \IN3008\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44123\,
                  I0 =>  \LVDAGD\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR08/\  
  \=44124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44124\,
                  I0 =>  \44123\,
                  I1 =>  \44122\,
                  I2 =>  \44217\,
                  I3 => \&43148\ );

  \=44125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44125\,
                  I0 =>  \IMUOPR\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44126\,
                  I0 =>  \LRRLSC\,
                  I1 =>  \44158\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR09/\  
  \=44127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44127\,
                  I0 =>  \44126\,
                  I1 =>  \44125\,
                  I2 =>  \44218\,
                  I3 => \&44354\ );

  \=44128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44128\,
                  I0 =>  \CTLSAT\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR10/\  
  \=44129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44129\,
                  I0 =>  \CH3310\,
                  I1 =>  \44128\,
                  I2 =>  \44219\,
                  I3 => \&44360\ );

  \=44130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44130\,
                  I0 =>  \IMUCAG\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44131\,
                  I0 =>  \LEMATT\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR11/\  
  \=44132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44132\,
                  I0 =>  \44131\,
                  I1 =>  \44130\,
                  I2 =>  \44220\,
                  I3 => \&44406\ );

  \=44133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44133\,
                  I0 =>  \CDUFAL\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44134\,
                  I0 =>  \IN3212\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR12/\  
  \=44135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44135\,
                  I0 =>  \44134\,
                  I1 =>  \44133\,
                  I2 =>  \44232\,
                  I3 => \&44412\ );

  \=44136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44136\,
                  I0 =>  \IMUFAL\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44137\,
                  I0 =>  \IN3213\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR13/\  
  \=44138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44138\,
                  I0 =>  \44137\,
                  I1 =>  \44136\,
                  I2 =>  \44233\,
                  I3 => \&44418\ );

  \=44139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44139\,
                  I0 =>  \ISSTOR\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44140\,
                  I0 =>  \IN3214\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR14/\  
  \=44141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44141\,
                  I0 =>  \44140\,
                  I1 =>  \44139\,
                  I2 =>  \44234\,
                  I3 => \&44424\ );

  \=44142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44142\,
                  I0 =>  \TEMPIN\,
                  I1 =>  \44146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44143\,
                  I0 =>  \IN3216\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR16/\  
  \=44144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44144\,
                  I0 =>  \44143\,
                  I1 =>  \44142\,
                  I2 =>  \44235\,
                  I3 => \&44430\ );

  \=44145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44145\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH30/\   
  \=44146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44146\,
                  I0 =>  \44145\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44149\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH31/\   
  \=44150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44150\,
                  I0 =>  \44149\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44153\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH32/\   
  \=44154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44154\,
                  I0 =>  \44153\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44157\,
                  I0 =>  \XB3/\,
                  I1 =>  \XT3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH33/\   
  \=44158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44158\,
                  I0 =>  \44157\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44201\,
                  I0 =>  \MANR+P\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44202\,
                  I0 =>  \MANR-P\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44203\,
                  I0 =>  \MANR+Y\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44204\,
                  I0 =>  \MANR-Y\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44205\,
                  I0 =>  \MANR+R\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44206\,
                  I0 =>  \MANR+P\,
                  I1 =>  \MANR-P\,
                  I2 =>  \MANR+Y\,
                  I3 => \&44207\ );

  -- Alias \44206\    
  \=44207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44207\,
                  I0 =>  \MANR-Y\,
                  I1 =>  \MANR+R\,
                  I2 =>  \MANR-R\,
                  I3 =>  '0' );

  \=44208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44208\,
                  I0 =>  \44213\,
                  I1 =>  \44206\,
                  I2 =>  \F05A/\,
                  I3 =>  '0' );

  \:44209\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44209\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44209\,
                   R => '0',
                   S => SYSRESET );

  \=44209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44209\,
                  I0 =>  \44208\,
                  I1 =>  \44210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44210\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44210\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44210\,
                   R => SYSRESET,
                   S => '0' );

  \=44210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44210\,
                  I0 =>  \44209\,
                  I1 =>  \44206\,
                  I2 =>  \F05D\,
                  I3 =>  '0' );

  -- Alias \TRP31A\   
  \=44211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44211\,
                  I0 =>  \44209\,
                  I1 =>  \F05B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44212\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44212\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44212\,
                   R => SYSRESET,
                   S => '0' );

  \=44212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44212\,
                  I0 =>  \44213\,
                  I1 =>  \GOJAM\,
                  I2 =>  \44211\,
                  I3 =>  '0' );

  \:44213\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44213\,
                   R => '0',
                   S => SYSRESET );

  \=44213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44213\,
                  I0 =>  \44214\,
                  I1 =>  \44212\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44214\,
                  I0 =>  \CHWL12/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44215\,
                  I0 =>  \MANR-R\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44216\,
                  I0 =>  \TRAN+X\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44217\,
                  I0 =>  \TRAN-X\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44218\,
                  I0 =>  \TRAN+Y\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44219\,
                  I0 =>  \TRAN-Y\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44220\,
                  I0 =>  \TRAN+Z\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44221\,
                  I0 =>  \TRAN+X\,
                  I1 =>  \TRAN-X\,
                  I2 =>  \TRAN+Y\,
                  I3 => \&44222\ );

  -- Alias \44221\    
  \=44222\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44222\,
                  I0 =>  \TRAN-Y\,
                  I1 =>  \TRAN+Z\,
                  I2 =>  \TRAN-Z\,
                  I3 =>  '0' );

  \=44223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44223\,
                  I0 =>  \44228\,
                  I1 =>  \F05A/\,
                  I2 =>  \44221\,
                  I3 =>  '0' );

  \:44224\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44224\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44224\,
                   R => '0',
                   S => SYSRESET );

  \=44224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44224\,
                  I0 =>  \44223\,
                  I1 =>  \44225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44225\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44225\,
                   R => SYSRESET,
                   S => '0' );

  \=44225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44225\,
                  I0 =>  \44224\,
                  I1 =>  \44221\,
                  I2 =>  \F05D\,
                  I3 =>  '0' );

  -- Alias \TRP31B\   
  \=44226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44226\,
                  I0 =>  \44224\,
                  I1 =>  \F05B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44227\,
                  I0 =>  \CHWL13/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44228\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44228\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44228\,
                   R => '0',
                   S => SYSRESET );

  \=44228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44228\,
                  I0 =>  \44227\,
                  I1 =>  \44229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44229\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44229\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44229\,
                   R => SYSRESET,
                   S => '0' );

  \=44229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44229\,
                  I0 =>  \44228\,
                  I1 =>  \GOJAM\,
                  I2 =>  \44226\,
                  I3 =>  '0' );

  \=44230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44230\,
                  I0 =>  \44211\,
                  I1 =>  \44226\,
                  I2 =>  \44253\,
                  I3 =>  '0' );

  -- Alias \HNDRPT\   
  \=44231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44231\,
                  I0 =>  \TPOR/\,
                  I1 =>  \44230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44232\,
                  I0 =>  \TRAN-Z\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44233\,
                  I0 =>  \HOLFUN\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44234\,
                  I0 =>  \FREFUN\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44235\,
                  I0 =>  \GCAPCL\,
                  I1 =>  \44150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3201\   
  \=44236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44236\,
                  I0 =>  \MNIM+P\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3206\   
  \=44237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44237\,
                  I0 =>  \44154\,
                  I1 =>  \MNIM-R\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3202\   
  \=44238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44238\,
                  I0 =>  \MNIM-P\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3207\   
  \=44239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44239\,
                  I0 =>  \44154\,
                  I1 =>  \TRST9\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3203\   
  \=44240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44240\,
                  I0 =>  \MNIM+Y\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3208\   
  \=44241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44241\,
                  I0 =>  \44154\,
                  I1 =>  \TRST10\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3204\   
  \=44242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44242\,
                  I0 =>  \MNIM-Y\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3209\   
  \=44243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44243\,
                  I0 =>  \44154\,
                  I1 =>  \PCHGOF\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3205\   
  \=44244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44244\,
                  I0 =>  \MNIM+R\,
                  I1 =>  \44154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3210\   
  \=44245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44245\,
                  I0 =>  \44154\,
                  I1 =>  \ROLGOF\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \44248\    
  \=44246\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44246\,
                  I0 =>  \ROLGOF\,
                  I1 =>  \PCHGOF\,
                  I2 =>  \TRST10\,
                  I3 => \&44247\ );

  -- Alias \44248\    
  \=44247\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44247\,
                  I0 =>  \TRST9\,
                  I1 =>  \MNIM-R\,
                  I2 =>  \MNIM+R\,
                  I3 => \&44249\ );

  \=44248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44248\,
                  I0 =>  \MNIM-Y\,
                  I1 =>  \MNIM+Y\,
                  I2 =>  \MNIM-P\,
                  I3 => \&44246\ );

  -- Alias \44248\    
  \=44249\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44249\,
                  I0 =>  \MNIM+P\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44250\,
                  I0 =>  \44255\,
                  I1 =>  \F05A/\,
                  I2 =>  \44248\,
                  I3 =>  '0' );

  \:44251\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44251\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44251\,
                   R => '0',
                   S => SYSRESET );

  \=44251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44251\,
                  I0 =>  \44250\,
                  I1 =>  \44252\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44252\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44252\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44252\,
                   R => SYSRESET,
                   S => '0' );

  \=44252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44252\,
                  I0 =>  \44251\,
                  I1 =>  \F05D\,
                  I2 =>  \44248\,
                  I3 =>  '0' );

  -- Alias \TRP32\    
  \=44253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44253\,
                  I0 =>  \F05B/\,
                  I1 =>  \44251\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44254\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44254\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44254\,
                   R => SYSRESET,
                   S => '0' );

  \=44254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44254\,
                  I0 =>  \44255\,
                  I1 =>  \44253\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \:44255\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44255\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44255\,
                   R => '0',
                   S => SYSRESET );

  \=44255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44255\,
                  I0 =>  \44256\,
                  I1 =>  \44254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44256\,
                  I0 =>  \CHWL14/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3316\   
  \=44257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44257\,
                  I0 =>  \OSCALM\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3314\   
  \=44258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44258\,
                  I0 =>  \AGCWAR\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3313\   
  \=44259\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44259\,
                  I0 =>  \PIPAFL\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ***************************
  -- ***                     ***
  -- ***  A17/2 - INOUT II.  ***
  -- ***                     ***
  -- ***************************

  \=44301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44301\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44302\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44302\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44302\,
                   R => '0',
                   S => SYSRESET );

  \=44302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44302\,
                  I0 =>  \44301\,
                  I1 =>  \44303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44303\,
                   R => SYSRESET,
                   S => '0' );

  \=44303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44303\,
                  I0 =>  \44302\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44304\,
                  I0 =>  \44441\,
                  I1 =>  \44302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB01\   
  \=44305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44305\,
                  I0 =>  \44302\,
                  I1 =>  \44302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR01/\  
  \=44306\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44306\,
                  I0 =>  \CH1301\,
                  I1 =>  \44304\,
                  I2 =>  \CH1401\,
                  I3 => \&48201\ );

  \=44307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44307\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44308\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44308\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44308\,
                   R => '0',
                   S => SYSRESET );

  \=44308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44308\,
                  I0 =>  \44307\,
                  I1 =>  \44309\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44309\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44309\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44309\,
                   R => SYSRESET,
                   S => '0' );

  \=44309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44309\,
                  I0 =>  \44308\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44310\,
                  I0 =>  \44441\,
                  I1 =>  \44308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB02\   
  \=44311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44311\,
                  I0 =>  \44308\,
                  I1 =>  \44308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR02/\  
  \=44312\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44312\,
                  I0 =>  \CH1302\,
                  I1 =>  \44310\,
                  I2 =>  \CH1402\,
                  I3 => \&48203\ );

  \=44313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44313\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44314\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44314\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44314\,
                   R => '0',
                   S => SYSRESET );

  \=44314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44314\,
                  I0 =>  \44313\,
                  I1 =>  \44315\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44315\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44315\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44315\,
                   R => SYSRESET,
                   S => '0' );

  \=44315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44315\,
                  I0 =>  \44314\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44316\,
                  I0 =>  \44441\,
                  I1 =>  \44314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB03\   
  \=44317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44317\,
                  I0 =>  \44314\,
                  I1 =>  \44314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR03/\  
  \=44318\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44318\,
                  I0 =>  \CH1303\,
                  I1 =>  \44316\,
                  I2 =>  \CH1403\,
                  I3 => \&48205\ );

  \=44319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44319\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44320\,
                   R => '0',
                   S => SYSRESET );

  \=44320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44320\,
                  I0 =>  \44319\,
                  I1 =>  \44321\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44321\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44321\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44321\,
                   R => SYSRESET,
                   S => '0' );

  \=44321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44321\,
                  I0 =>  \44320\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44322\,
                  I0 =>  \44441\,
                  I1 =>  \44320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB04\   
  \=44323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44323\,
                  I0 =>  \44320\,
                  I1 =>  \44320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR04/\  
  \=44324\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44324\,
                  I0 =>  \CH1304\,
                  I1 =>  \44322\,
                  I2 =>  \CH1404\,
                  I3 => \&48207\ );

  \=44325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44325\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44326\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44326\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44326\,
                   R => '0',
                   S => SYSRESET );

  \=44326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44326\,
                  I0 =>  \44325\,
                  I1 =>  \44327\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44327\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44327\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44327\,
                   R => SYSRESET,
                   S => '0' );

  \=44327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44327\,
                  I0 =>  \44326\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44328\,
                  I0 =>  \44441\,
                  I1 =>  \44326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB05\   
  \=44329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44329\,
                  I0 =>  \44326\,
                  I1 =>  \44326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR05/\  
  \=44330\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44330\,
                  I0 =>  \CH1305\,
                  I1 =>  \44328\,
                  I2 =>  \CH1405\,
                  I3 => \&48209\ );

  \=44331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44331\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44332\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44332\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44332\,
                   R => '0',
                   S => SYSRESET );

  \=44332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44332\,
                  I0 =>  \44331\,
                  I1 =>  \44333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44333\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44333\,
                   R => SYSRESET,
                   S => '0' );

  \=44333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44333\,
                  I0 =>  \44332\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44334\,
                  I0 =>  \44441\,
                  I1 =>  \44332\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB06\   
  \=44335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44335\,
                  I0 =>  \44332\,
                  I1 =>  \44332\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR06/\  
  \=44336\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44336\,
                  I0 =>  \CH1306\,
                  I1 =>  \44334\,
                  I2 =>  \CH1406\,
                  I3 => \&48212\ );

  \=44337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44337\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44338\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44338\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44338\,
                   R => '0',
                   S => SYSRESET );

  \=44338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44338\,
                  I0 =>  \44337\,
                  I1 =>  \44339\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44339\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44339\,
                   R => SYSRESET,
                   S => '0' );

  \=44339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44339\,
                  I0 =>  \44338\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44340\,
                  I0 =>  \44441\,
                  I1 =>  \44338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB07\   
  \=44341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44341\,
                  I0 =>  \44338\,
                  I1 =>  \44338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR07/\  
  \=44342\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44342\,
                  I0 =>  \CH1307\,
                  I1 =>  \44340\,
                  I2 =>  \CH1407\,
                  I3 => \&48214\ );

  \=44343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44343\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44344\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44344\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44344\,
                   R => '0',
                   S => SYSRESET );

  \=44344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44344\,
                  I0 =>  \44343\,
                  I1 =>  \44345\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44345\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44345\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44345\,
                   R => SYSRESET,
                   S => '0' );

  \=44345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44345\,
                  I0 =>  \44344\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44346\,
                  I0 =>  \44441\,
                  I1 =>  \44344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB08\   
  \=44347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44347\,
                  I0 =>  \44344\,
                  I1 =>  \44344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR08/\  
  \=44348\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44348\,
                  I0 =>  \CH1308\,
                  I1 =>  \44346\,
                  I2 =>  \CH1408\,
                  I3 => \&48216\ );

  \=44349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44349\,
                  I0 =>  \CHWL09/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44350\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44350\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44350\,
                   R => '0',
                   S => SYSRESET );

  \=44350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44350\,
                  I0 =>  \44349\,
                  I1 =>  \44351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44351\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44351\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44351\,
                   R => SYSRESET,
                   S => '0' );

  \=44351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44351\,
                  I0 =>  \44350\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44352\,
                  I0 =>  \44441\,
                  I1 =>  \44350\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB09\   
  \=44353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44353\,
                  I0 =>  \44350\,
                  I1 =>  \44350\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR09/\  
  \=44354\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44354\,
                  I0 =>  \CH1309\,
                  I1 =>  \44352\,
                  I2 =>  \CH1409\,
                  I3 => \&48438\ );

  \=44355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44355\,
                  I0 =>  \CHWL10/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44356\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44356\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44356\,
                   R => '0',
                   S => SYSRESET );

  \=44356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44356\,
                  I0 =>  \44355\,
                  I1 =>  \44357\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44357\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44357\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44357\,
                   R => SYSRESET,
                   S => '0' );

  \=44357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44357\,
                  I0 =>  \44356\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44358\,
                  I0 =>  \44441\,
                  I1 =>  \44356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB10\   
  \=44359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44359\,
                  I0 =>  \44356\,
                  I1 =>  \44356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR10/\  
  \=44360\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44360\,
                  I0 =>  \CH1310\,
                  I1 =>  \44358\,
                  I2 =>  \CH1410\,
                  I3 => \&48456\ );

  \=44401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44401\,
                  I0 =>  \CHWL11/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44402\,
                   R => '0',
                   S => SYSRESET );

  \=44402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44402\,
                  I0 =>  \44401\,
                  I1 =>  \44403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44403\,
                   R => SYSRESET,
                   S => '0' );

  \=44403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44403\,
                  I0 =>  \44402\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44404\,
                  I0 =>  \44441\,
                  I1 =>  \44402\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RLYB11\   
  \=44405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44405\,
                  I0 =>  \44402\,
                  I1 =>  \44402\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR11/\  
  \=44406\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44406\,
                  I0 =>  \CH1311\,
                  I1 =>  \44404\,
                  I2 =>  \CH1411\,
                  I3 => \&45435\ );

  \=44407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44407\,
                  I0 =>  \CHWL12/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44408\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44408\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44408\,
                   R => '0',
                   S => SYSRESET );

  \=44408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44408\,
                  I0 =>  \44407\,
                  I1 =>  \44409\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44409\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44409\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44409\,
                   R => SYSRESET,
                   S => '0' );

  \=44409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44409\,
                  I0 =>  \44408\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44410\,
                  I0 =>  \44441\,
                  I1 =>  \44408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RYWD12\   
  \=44411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44411\,
                  I0 =>  \44408\,
                  I1 =>  \44408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR12/\  
  \=44412\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44412\,
                  I0 =>  \CH3312\,
                  I1 =>  \44410\,
                  I2 =>  \CH1412\,
                  I3 => \&45438\ );

  \=44413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44413\,
                  I0 =>  \CHWL13/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44414\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44414\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44414\,
                   R => '0',
                   S => SYSRESET );

  \=44414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44414\,
                  I0 =>  \44413\,
                  I1 =>  \44415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44415\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44415\,
                   R => SYSRESET,
                   S => '0' );

  \=44415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44415\,
                  I0 =>  \44414\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44416\,
                  I0 =>  \44441\,
                  I1 =>  \44414\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RYWD13\   
  \=44417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44417\,
                  I0 =>  \44414\,
                  I1 =>  \44414\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR13/\  
  \=44418\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44418\,
                  I0 =>  \CH1213\,
                  I1 =>  \44416\,
                  I2 =>  \CH1413\,
                  I3 => \&44461\ );

  \=44419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44419\,
                  I0 =>  \CHWL14/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44420\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44420\,
                   R => '0',
                   S => SYSRESET );

  \=44420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44420\,
                  I0 =>  \44419\,
                  I1 =>  \44421\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44421\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44421\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44421\,
                   R => SYSRESET,
                   S => '0' );

  \=44421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44421\,
                  I0 =>  \44420\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44422\,
                  I0 =>  \44441\,
                  I1 =>  \44420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RYWD14\   
  \=44423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44423\,
                  I0 =>  \44420\,
                  I1 =>  \44420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR14/\  
  \=44424\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44424\,
                  I0 =>  \CH1214\,
                  I1 =>  \44422\,
                  I2 =>  \CH1414\,
                  I3 => \&45443\ );

  \=44425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44425\,
                  I0 =>  \CHWL16/\,
                  I1 =>  \44432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44426\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \44426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44426\,
                   R => '0',
                   S => SYSRESET );

  \=44426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44426\,
                  I0 =>  \44425\,
                  I1 =>  \44427\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:44427\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \44427\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$44427\,
                   R => SYSRESET,
                   S => '0' );

  \=44427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$44427\,
                  I0 =>  \44426\,
                  I1 =>  \44437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44428\,
                  I0 =>  \44441\,
                  I1 =>  \44426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RYWD16\   
  \=44429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44429\,
                  I0 =>  \44426\,
                  I1 =>  \44426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR16/\  
  \=44430\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44430\,
                  I0 =>  \CH1316\,
                  I1 =>  \44428\,
                  I2 =>  \CH1416\,
                  I3 => \&45445\ );

  \=44431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44431\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XT1/\,
                  I2 =>  \XB0/\,
                  I3 =>  '0' );

  -- Alias \WCH10/\   
  \=44432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44432\,
                  I0 =>  \44431\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44435\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XB0/\,
                  I2 =>  \XT1/\,
                  I3 =>  '0' );

  \=44436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44436\,
                  I0 =>  \44435\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH10\    
  \=44437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44437\,
                  I0 =>  \44436\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44440\,
                  I0 =>  \XB0/\,
                  I1 =>  \XT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH10/\   
  \=44441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44441\,
                  I0 =>  \44440\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44444\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XT1/\,
                  I2 =>  \XB1/\,
                  I3 =>  '0' );

  -- Alias \WCH11/\   
  \=44445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44445\,
                  I0 =>  \44444\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44448\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XB1/\,
                  I2 =>  \XT1/\,
                  I3 =>  '0' );

  \=44449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44449\,
                  I0 =>  \GOJAM\,
                  I1 =>  \44448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH11\    
  \=44450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44450\,
                  I0 =>  \44449\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=44453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44453\,
                  I0 =>  \XB1/\,
                  I1 =>  \XT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH11/\   
  \=44454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44454\,
                  I0 =>  \44453\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR13/\  
  \=44461\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&44461\,
                  I0 =>  \CH1113\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&45441\ );

  -- Alias \XBC\      
  \=44462\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \44462\,
                  I0 =>  \S01\,
                  I1 =>  \S02\,
                  I2 =>  \S03\,
                  I3 =>  '0' );

  -- ****************************
  -- ***                      ***
  -- ***  A18/1 - INOUT III.  ***
  -- ***                      ***
  -- ****************************

  \:45101\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45101\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45101\,
                   R => '0',
                   S => SYSRESET );

  \=45101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45101\,
                  I0 =>  \MKEY1\,
                  I1 =>  \45102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45102\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45102\,
                   R => SYSRESET,
                   S => '0' );

  \=45102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45102\,
                  I0 =>  \45101\,
                  I1 =>  \45123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1501\   
  \=45103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45103\,
                  I0 =>  \45124\,
                  I1 =>  \45101\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45104\,
                  I0 =>  \45101\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45105\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45105\,
                   R => '0',
                   S => SYSRESET );

  \=45105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45105\,
                  I0 =>  \MKEY2\,
                  I1 =>  \45106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45106\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45106\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45106\,
                   R => SYSRESET,
                   S => '0' );

  \=45106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45106\,
                  I0 =>  \45105\,
                  I1 =>  \45123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1502\   
  \=45107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45107\,
                  I0 =>  \45124\,
                  I1 =>  \45105\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45108\,
                  I0 =>  \45105\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45109\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45109\,
                   R => '0',
                   S => SYSRESET );

  \=45109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45109\,
                  I0 =>  \MKEY3\,
                  I1 =>  \45110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45110\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45110\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45110\,
                   R => SYSRESET,
                   S => '0' );

  \=45110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45110\,
                  I0 =>  \45109\,
                  I1 =>  \45123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1503\   
  \=45111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45111\,
                  I0 =>  \45124\,
                  I1 =>  \45109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45112\,
                  I0 =>  \45109\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45113\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45113\,
                   R => '0',
                   S => SYSRESET );

  \=45113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45113\,
                  I0 =>  \MKEY4\,
                  I1 =>  \45114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45114\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45114\,
                   R => SYSRESET,
                   S => '0' );

  \=45114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45114\,
                  I0 =>  \45113\,
                  I1 =>  \45123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1504\   
  \=45115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45115\,
                  I0 =>  \45124\,
                  I1 =>  \45113\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45116\,
                  I0 =>  \45113\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45117\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45117\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45117\,
                   R => '0',
                   S => SYSRESET );

  \=45117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45117\,
                  I0 =>  \MKEY5\,
                  I1 =>  \45118\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45118\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45118\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45118\,
                   R => SYSRESET,
                   S => '0' );

  \=45118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45118\,
                  I0 =>  \45117\,
                  I1 =>  \45123\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1505\   
  \=45119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45119\,
                  I0 =>  \45124\,
                  I1 =>  \45117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45120\,
                  I0 =>  \45117\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45121\,
                  I0 =>  \MAINRS\,
                  I1 =>  \MAINRS\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45122\,
                  I0 =>  \XT1/\,
                  I1 =>  \XB5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45123\,
                  I0 =>  \45121\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH15/\   
  \=45124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45124\,
                  I0 =>  \45122\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45126\    
  \=45125\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45125\,
                  I0 =>  \45104\,
                  I1 =>  \45108\,
                  I2 =>  \45112\,
                  I3 =>  '0' );

  \=45126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45126\,
                  I0 =>  \45116\,
                  I1 =>  \45120\,
                  I2 =>  '0',
                  I3 => \&45125\ );

  \=45127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45127\,
                  I0 =>  \F09A/\,
                  I1 =>  \45126\,
                  I2 =>  \45135\,
                  I3 => \&45132\ );

  -- Alias \TPOR/\    
  \=45128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45128\,
                  I0 =>  \T05\,
                  I1 =>  \T11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45129\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45129\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45129\,
                   R => '0',
                   S => SYSRESET );

  \=45129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45129\,
                  I0 =>  \45127\,
                  I1 =>  \45130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45130\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45130\,
                   R => SYSRESET,
                   S => '0' );

  \=45130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45130\,
                  I0 =>  \45129\,
                  I1 =>  \45126\,
                  I2 =>  \F09D\,
                  I3 =>  '0' );

  -- Alias \KYRPT1\   
  \=45131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45131\,
                  I0 =>  \45128\,
                  I1 =>  \45129\,
                  I2 =>  \F09B/\,
                  I3 =>  '0' );

  -- Alias \45127\    
  \=45132\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45132\,
                  I0 =>  \45123\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45133\,
                  I0 =>  \45126\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45134\,
                  I0 =>  \45133\,
                  I1 =>  \45121\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45135\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45135\,
                   R => SYSRESET,
                   S => '0' );

  \=45135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45135\,
                  I0 =>  \45134\,
                  I1 =>  \45136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45136\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45136\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45136\,
                   R => '0',
                   S => SYSRESET );

  \=45136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45136\,
                  I0 =>  \45135\,
                  I1 =>  \45131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45137\,
                  I0 =>  \WCH13/\,
                  I1 =>  \CHWL11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45138\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45138\,
                   R => '0',
                   S => SYSRESET );

  \=45138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45138\,
                  I0 =>  \45137\,
                  I1 =>  \45139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45139\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45139\,
                   R => SYSRESET,
                   S => '0' );

  \=45139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45139\,
                  I0 =>  \45138\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1311\   
  \=45140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45140\,
                  I0 =>  \45138\,
                  I1 =>  \RCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45141\,
                  I0 =>  \SBYBUT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45142\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45142\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45142\,
                   R => '0',
                   S => SYSRESET );

  \=45142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45142\,
                  I0 =>  \45147\,
                  I1 =>  \45146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45143\,
                  I0 =>  \F17A/\,
                  I1 =>  \45141\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45144\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45144\,
                   R => SYSRESET,
                   S => '0' );

  \=45144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45144\,
                  I0 =>  \45145\,
                  I1 =>  \45141\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45145\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45145\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45145\,
                   R => '0',
                   S => SYSRESET );

  \=45145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45145\,
                  I0 =>  \45143\,
                  I1 =>  \45144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45146\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45146\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45146\,
                   R => SYSRESET,
                   S => '0' );

  \=45146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45146\,
                  I0 =>  \45142\,
                  I1 =>  \45141\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45147\,
                  I0 =>  \F17B/\,
                  I1 =>  \45145\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBY\      
  \=45148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45148\,
                  I0 =>  \45153\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45149\,
                  I0 =>  \45142\,
                  I1 =>  \STOP\,
                  I2 =>  \45138\,
                  I3 =>  '0' );

  \:45150\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45150\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45150\,
                   R => '0',
                   S => SYSRESET );

  \=45150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45150\,
                  I0 =>  \45149\,
                  I1 =>  \45151\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45151\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45151\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45151\,
                   R => SYSRESET,
                   S => '0' );

  \=45151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45151\,
                  I0 =>  \45150\,
                  I1 =>  \45142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45152\,
                  I0 =>  \45151\,
                  I1 =>  \45142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STNDBY/\  
  \=45153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45153\,
                  I0 =>  \45155\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45154\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45154\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45154\,
                   R => '0',
                   S => SYSRESET );

  \=45154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45154\,
                  I0 =>  \45151\,
                  I1 =>  \45155\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STNDBY\   
  \:45155\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45155\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45155\,
                   R => SYSRESET,
                   S => '0' );

  \=45155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45155\,
                  I0 =>  \45154\,
                  I1 =>  \45152\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45156\,
                  I0 =>  \45155\,
                  I1 =>  \ALTEST\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SBYLIT\   
  \=45157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45157\,
                  I0 =>  \45156\,
                  I1 =>  \45156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F17A/\    
  \=45159\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45159\,
                  I0 =>  \F17A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45250\    
  \=45160\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45160\,
                  I0 =>  \45234\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45201\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45201\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45201\,
                   R => '0',
                   S => SYSRESET );

  \=45201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45201\,
                  I0 =>  \NKEY1\,
                  I1 =>  \45202\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45202\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45202\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45202\,
                   R => SYSRESET,
                   S => '0' );

  \=45202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45202\,
                  I0 =>  \45201\,
                  I1 =>  \45223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1601\   
  \=45203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45203\,
                  I0 =>  \45236\,
                  I1 =>  \45201\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45204\,
                  I0 =>  \45201\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45205\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45205\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45205\,
                   R => '0',
                   S => SYSRESET );

  \=45205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45205\,
                  I0 =>  \NKEY2\,
                  I1 =>  \45206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45206\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45206\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45206\,
                   R => SYSRESET,
                   S => '0' );

  \=45206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45206\,
                  I0 =>  \45205\,
                  I1 =>  \45223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1602\   
  \=45207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45207\,
                  I0 =>  \45236\,
                  I1 =>  \45205\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45208\,
                  I0 =>  \45205\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45209\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45209\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45209\,
                   R => '0',
                   S => SYSRESET );

  \=45209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45209\,
                  I0 =>  \NKEY3\,
                  I1 =>  \45210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45210\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45210\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45210\,
                   R => SYSRESET,
                   S => '0' );

  \=45210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45210\,
                  I0 =>  \45209\,
                  I1 =>  \45223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1603\   
  \=45211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45211\,
                  I0 =>  \45236\,
                  I1 =>  \45209\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45212\,
                  I0 =>  \45209\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45213\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45213\,
                   R => '0',
                   S => SYSRESET );

  \=45213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45213\,
                  I0 =>  \NKEY4\,
                  I1 =>  \45214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45214\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45214\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45214\,
                   R => SYSRESET,
                   S => '0' );

  \=45214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45214\,
                  I0 =>  \45213\,
                  I1 =>  \45223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1604\   
  \=45215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45215\,
                  I0 =>  \45236\,
                  I1 =>  \45213\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45216\,
                  I0 =>  \45213\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45217\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45217\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45217\,
                   R => '0',
                   S => SYSRESET );

  \=45217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45217\,
                  I0 =>  \NKEY5\,
                  I1 =>  \45218\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45218\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45218\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45218\,
                   R => SYSRESET,
                   S => '0' );

  \=45218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45218\,
                  I0 =>  \45217\,
                  I1 =>  \45223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1605\   
  \=45219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45219\,
                  I0 =>  \45236\,
                  I1 =>  \45217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45220\,
                  I0 =>  \45217\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45221\,
                  I0 =>  \NAVRST\,
                  I1 =>  \NAVRST\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45222\,
                  I0 =>  \CAURST\,
                  I1 =>  \W1110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45223\,
                  I0 =>  \45221\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ERRST\    
  \=45224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45224\,
                  I0 =>  \45222\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45225\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45225\,
                   R => '0',
                   S => SYSRESET );

  \=45225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45225\,
                  I0 =>  \MARK\,
                  I1 =>  \45226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45226\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45226\,
                   R => SYSRESET,
                   S => '0' );

  \=45226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45226\,
                  I0 =>  \45225\,
                  I1 =>  \45234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1606\   
  \=45227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45227\,
                  I0 =>  \45236\,
                  I1 =>  \45225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45228\,
                  I0 =>  \45225\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45229\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45229\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45229\,
                   R => '0',
                   S => SYSRESET );

  \=45229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45229\,
                  I0 =>  \MRKREJ\,
                  I1 =>  \45230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45230\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45230\,
                   R => SYSRESET,
                   S => '0' );

  \=45230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45230\,
                  I0 =>  \45229\,
                  I1 =>  \45234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1607\   
  \=45231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45231\,
                  I0 =>  \45236\,
                  I1 =>  \45229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45232\,
                  I0 =>  \45229\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45233\,
                  I0 =>  \MRKRST\,
                  I1 =>  \MRKRST\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45234\,
                  I0 =>  \45233\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45235\,
                  I0 =>  \XT1/\,
                  I1 =>  \XB6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH16/\   
  \=45236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45236\,
                  I0 =>  \45235\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45239\    
  \=45238\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45238\,
                  I0 =>  \45204\,
                  I1 =>  \45208\,
                  I2 =>  \45212\,
                  I3 =>  '0' );

  \=45239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45239\,
                  I0 =>  \45216\,
                  I1 =>  \45220\,
                  I2 =>  '0',
                  I3 => \&45238\ );

  \=45240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45240\,
                  I0 =>  \F09A/\,
                  I1 =>  \45239\,
                  I2 =>  \45247\,
                  I3 => \&45243\ );

  \:45241\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45241\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45241\,
                   R => '0',
                   S => SYSRESET );

  \=45241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45241\,
                  I0 =>  \45240\,
                  I1 =>  \45242\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45242\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45242\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45242\,
                   R => SYSRESET,
                   S => '0' );

  \=45242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45242\,
                  I0 =>  \45241\,
                  I1 =>  \45239\,
                  I2 =>  \F09D\,
                  I3 =>  '0' );

  -- Alias \45240\    
  \=45243\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45243\,
                  I0 =>  \45223\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \KYRPT2\   
  \=45244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45244\,
                  I0 =>  \F09B/\,
                  I1 =>  \45241\,
                  I2 =>  \TPOR/\,
                  I3 =>  '0' );

  \=45245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45245\,
                  I0 =>  \45239\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45246\,
                  I0 =>  \45245\,
                  I1 =>  \45221\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45247\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45247\,
                   R => SYSRESET,
                   S => '0' );

  \=45247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45247\,
                  I0 =>  \45246\,
                  I1 =>  \45248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45248\,
                   R => '0',
                   S => SYSRESET );

  \=45248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45248\,
                  I0 =>  \45247\,
                  I1 =>  \45244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45249\,
                  I0 =>  \45228\,
                  I1 =>  \45232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45250\,
                  I0 =>  \F09A/\,
                  I1 =>  \45249\,
                  I2 =>  \45257\,
                  I3 => \&45160\ );

  \:45251\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45251\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45251\,
                   R => '0',
                   S => SYSRESET );

  \=45251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45251\,
                  I0 =>  \45250\,
                  I1 =>  \45252\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45252\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45252\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45252\,
                   R => SYSRESET,
                   S => '0' );

  \=45252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45252\,
                  I0 =>  \45251\,
                  I1 =>  \45249\,
                  I2 =>  \F09D\,
                  I3 =>  '0' );

  -- Alias \MKRPT\    
  \=45254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45254\,
                  I0 =>  \TPOR/\,
                  I1 =>  \45251\,
                  I2 =>  \F09B/\,
                  I3 =>  '0' );

  \=45255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45255\,
                  I0 =>  \45249\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45256\,
                  I0 =>  \45255\,
                  I1 =>  \45233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45257\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45257\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45257\,
                   R => SYSRESET,
                   S => '0' );

  \=45257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45257\,
                  I0 =>  \45256\,
                  I1 =>  \45258\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45258\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45258\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45258\,
                   R => '0',
                   S => SYSRESET );

  \=45258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45258\,
                  I0 =>  \45257\,
                  I1 =>  \45254\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F17B/\    
  \=45261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45261\,
                  I0 =>  \F17B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TEMPIN/\  
  \=45262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45262\,
                  I0 =>  \TEMPIN\,
                  I1 =>  \TEMPIN\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************
  -- ***                      ***
  -- ***  A18/2 - INOUT III.  ***
  -- ***                      ***
  -- ****************************

  \=45301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45301\,
                  I0 =>  \CHWL04/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45302\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45302\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45302\,
                   R => '0',
                   S => SYSRESET );

  \=45302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45302\,
                  I0 =>  \45301\,
                  I1 =>  \45303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45303\,
                   R => SYSRESET,
                   S => '0' );

  \=45303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45303\,
                  I0 =>  \45302\,
                  I1 =>  \CCH13\,
                  I2 =>  \45342\,
                  I3 =>  '0' );

  -- Alias \CH1304\   
  \=45304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45304\,
                  I0 =>  \RCH13/\,
                  I1 =>  \45302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45305\,
                  I0 =>  \45303\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45306\,
                  I0 =>  \CHWL03/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45307\,
                   R => '0',
                   S => SYSRESET );

  \=45307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45307\,
                  I0 =>  \45306\,
                  I1 =>  \45308\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45308\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45308\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45308\,
                   R => SYSRESET,
                   S => '0' );

  \=45308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45308\,
                  I0 =>  \45307\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1303\   
  \=45309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45309\,
                  I0 =>  \RCH13/\,
                  I1 =>  \45307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45310\,
                  I0 =>  \45307\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45311\,
                  I0 =>  \45308\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45312\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45313\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45313\,
                   R => '0',
                   S => SYSRESET );

  \=45313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45313\,
                  I0 =>  \45312\,
                  I1 =>  \45314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45314\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45314\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45314\,
                   R => SYSRESET,
                   S => '0' );

  \=45314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45314\,
                  I0 =>  \45313\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1302\   
  \=45315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45315\,
                  I0 =>  \45313\,
                  I1 =>  \RCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45316\,
                  I0 =>  \WCH13/\,
                  I1 =>  \CHWL01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45317\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45317\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45317\,
                   R => '0',
                   S => SYSRESET );

  \=45317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45317\,
                  I0 =>  \45316\,
                  I1 =>  \45318\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45318\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45318\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45318\,
                   R => SYSRESET,
                   S => '0' );

  \=45318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45318\,
                  I0 =>  \45317\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1301\   
  \=45319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45319\,
                  I0 =>  \RCH13/\,
                  I1 =>  \45317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45320\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45320\,
                   R => '0',
                   S => SYSRESET );

  \=45320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45320\,
                  I0 =>  \45404\,
                  I1 =>  \45321\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45321\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45321\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45321\,
                   R => SYSRESET,
                   S => '0' );

  \=45321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45321\,
                  I0 =>  \45320\,
                  I1 =>  \45434\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=45322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45322\,
                  I0 =>  \45310\,
                  I1 =>  \45320\,
                  I2 =>  \F5BSB2/\,
                  I3 =>  '0' );

  \=45323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45323\,
                  I0 =>  \F5BSB2/\,
                  I1 =>  \45320\,
                  I2 =>  \45311\,
                  I3 =>  '0' );

  \=45324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45324\,
                  I0 =>  \45322\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45325\,
                  I0 =>  \45323\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45326\,
                  I0 =>  \45434\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45327\,
                  I0 =>  \45326\,
                  I1 =>  \GTSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RRRANG\   
  \=45328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45328\,
                  I0 =>  \45314\,
                  I1 =>  \45317\,
                  I2 =>  \45324\,
                  I3 =>  '0' );

  -- Alias \RRRARA\   
  \=45329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45329\,
                  I0 =>  \45324\,
                  I1 =>  \45318\,
                  I2 =>  \45313\,
                  I3 =>  '0' );

  -- Alias \LRXVEL\   
  \=45330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45330\,
                  I0 =>  \45318\,
                  I1 =>  \45314\,
                  I2 =>  \45325\,
                  I3 =>  '0' );

  -- Alias \LRYVEL\   
  \=45331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45331\,
                  I0 =>  \45325\,
                  I1 =>  \45317\,
                  I2 =>  \45314\,
                  I3 =>  '0' );

  -- Alias \LRZVEL\   
  \=45332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45332\,
                  I0 =>  \45325\,
                  I1 =>  \45313\,
                  I2 =>  \45318\,
                  I3 =>  '0' );

  -- Alias \LRRANG\   
  \=45333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45333\,
                  I0 =>  \45325\,
                  I1 =>  \45313\,
                  I2 =>  \45317\,
                  I3 =>  '0' );

  \=45334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45334\,
                  I0 =>  \45318\,
                  I1 =>  \45314\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45335\,
                  I0 =>  \45334\,
                  I1 =>  \45310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45336\,
                  I0 =>  \45335\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45337\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45337\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45337\,
                   R => '0',
                   S => SYSRESET );

  \=45337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45337\,
                  I0 =>  \45327\,
                  I1 =>  \45338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45338\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45338\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45338\,
                   R => SYSRESET,
                   S => '0' );

  \=45338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45338\,
                  I0 =>  \45337\,
                  I1 =>  \45342\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=45339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45339\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \45337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45340\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45340\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45340\,
                   R => '0',
                   S => SYSRESET );

  \=45340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45340\,
                  I0 =>  \45339\,
                  I1 =>  \45341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45341\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45341\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45341\,
                   R => SYSRESET,
                   S => '0' );

  \=45341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45341\,
                  I0 =>  \45340\,
                  I1 =>  \GOJAM\,
                  I2 =>  \F09B\,
                  I3 =>  '0' );

  -- Alias \RADRPT\   
  \=45342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45342\,
                  I0 =>  \45340\,
                  I1 =>  \45340\,
                  I2 =>  \TPORA/\,
                  I3 => \&45343\ );

  -- Alias \45342\    
  \=45343\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45343\,
                  I0 =>  \TPORA/\,
                  I1 =>  \GTRST/\,
                  I2 =>  \GTRST/\,
                  I3 =>  '0' );

  \=45344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45344\,
                  I0 =>  \45339\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RRSYNC\   
  \=45345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45345\,
                  I0 =>  \45336\,
                  I1 =>  \45344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \LRSYNC\   
  \=45346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45346\,
                  I0 =>  \45344\,
                  I1 =>  \45311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45347\,
                  I0 =>  \RRIN1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45348\,
                  I0 =>  \45336\,
                  I1 =>  \45347\,
                  I2 =>  \45305\,
                  I3 =>  '0' );

  \=45349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45349\,
                  I0 =>  \RRIN0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45350\,
                  I0 =>  \45336\,
                  I1 =>  \45349\,
                  I2 =>  \45305\,
                  I3 =>  '0' );

  \=45351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45351\,
                  I0 =>  \45348\,
                  I1 =>  \45354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RNRADP\   
  \=45352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45352\,
                  I0 =>  \45351\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45353\,
                  I0 =>  \LRIN1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45354\,
                  I0 =>  \45311\,
                  I1 =>  \45353\,
                  I2 =>  \45305\,
                  I3 =>  '0' );

  \=45355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45355\,
                  I0 =>  \LRIN0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45356\,
                  I0 =>  \45311\,
                  I1 =>  \45355\,
                  I2 =>  \45305\,
                  I3 =>  '0' );

  \=45357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45357\,
                  I0 =>  \45350\,
                  I1 =>  \45356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RNRADM\   
  \=45358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45358\,
                  I0 =>  \45357\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TPORA/\   
  \=45359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45359\,
                  I0 =>  \HERB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \HERB\     
  \=45360\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45360\,
                  I0 =>  \TPOR/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F10AS0\   
  \=45401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45401\,
                  I0 =>  \F10A/\,
                  I1 =>  \SB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45402\,
                   R => '0',
                   S => SYSRESET );

  \=45402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45402\,
                  I0 =>  \45401\,
                  I1 =>  \45403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45403\,
                   R => SYSRESET,
                   S => '0' );

  \=45403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45403\,
                  I0 =>  \45402\,
                  I1 =>  \45302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45404\,
                  I0 =>  \F10A/\,
                  I1 =>  \45402\,
                  I2 =>  \SB2/\,
                  I3 =>  '0' );

  \:45405\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45405\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45405\,
                   R => SYSRESET,
                   S => '0' );

  \=45405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45405\,
                  I0 =>  \45410\,
                  I1 =>  \45342\,
                  I2 =>  \45407\,
                  I3 =>  '0' );

  -- Alias \45407\    
  \=45406\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45406\,
                  I0 =>  \45405\,
                  I1 =>  \45342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45407\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45407\,
                   R => SYSRESET,
                   S => '0' );

  \=45407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45407\,
                  I0 =>  \45404\,
                  I1 =>  \45408\,
                  I2 =>  '0',
                  I3 => \&45406\ );

  \:45408\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45408\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45408\,
                   R => '0',
                   S => SYSRESET );

  \=45408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45408\,
                  I0 =>  \45407\,
                  I1 =>  \45404\,
                  I2 =>  \45409\,
                  I3 =>  '0' );

  \:45409\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45409\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45409\,
                   R => SYSRESET,
                   S => '0' );

  \=45409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45409\,
                  I0 =>  \45408\,
                  I1 =>  \45411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45410\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45410\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45410\,
                   R => '0',
                   S => SYSRESET );

  \=45410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45410\,
                  I0 =>  \45407\,
                  I1 =>  \45411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45411\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45411\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45411\,
                   R => SYSRESET,
                   S => '0' );

  \=45411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45411\,
                  I0 =>  \45410\,
                  I1 =>  \45408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45412\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45412\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45412\,
                   R => SYSRESET,
                   S => '0' );

  \=45412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45412\,
                  I0 =>  \45417\,
                  I1 =>  \45414\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45414\    
  \=45413\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45413\,
                  I0 =>  \45412\,
                  I1 =>  \45342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45414\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45414\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45414\,
                   R => SYSRESET,
                   S => '0' );

  \=45414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45414\,
                  I0 =>  \45405\,
                  I1 =>  \45415\,
                  I2 =>  '0',
                  I3 => \&45413\ );

  \:45415\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45415\,
                   R => '0',
                   S => SYSRESET );

  \=45415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45415\,
                  I0 =>  \45414\,
                  I1 =>  \45405\,
                  I2 =>  \45416\,
                  I3 =>  '0' );

  \:45416\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45416\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45416\,
                   R => SYSRESET,
                   S => '0' );

  \=45416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45416\,
                  I0 =>  \45415\,
                  I1 =>  \45418\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45417\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45417\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45417\,
                   R => '0',
                   S => SYSRESET );

  \=45417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45417\,
                  I0 =>  \45414\,
                  I1 =>  \45418\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45418\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45418\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45418\,
                   R => SYSRESET,
                   S => '0' );

  \=45418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45418\,
                  I0 =>  \45417\,
                  I1 =>  \45415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45419\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45419\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45419\,
                   R => SYSRESET,
                   S => '0' );

  \=45419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45419\,
                  I0 =>  \45424\,
                  I1 =>  \45421\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45421\    
  \=45420\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45420\,
                  I0 =>  \45419\,
                  I1 =>  \45342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45421\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45421\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45421\,
                   R => SYSRESET,
                   S => '0' );

  \=45421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45421\,
                  I0 =>  \45412\,
                  I1 =>  \45422\,
                  I2 =>  '0',
                  I3 => \&45420\ );

  \:45422\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45422\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45422\,
                   R => '0',
                   S => SYSRESET );

  \=45422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45422\,
                  I0 =>  \45421\,
                  I1 =>  \45412\,
                  I2 =>  \45423\,
                  I3 =>  '0' );

  \:45423\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45423\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45423\,
                   R => SYSRESET,
                   S => '0' );

  \=45423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45423\,
                  I0 =>  \45422\,
                  I1 =>  \45425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45424\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45424\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45424\,
                   R => '0',
                   S => SYSRESET );

  \=45424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45424\,
                  I0 =>  \45421\,
                  I1 =>  \45425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45425\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45425\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45425\,
                   R => SYSRESET,
                   S => '0' );

  \=45425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45425\,
                  I0 =>  \45424\,
                  I1 =>  \45422\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45426\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45426\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45426\,
                   R => SYSRESET,
                   S => '0' );

  \=45426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45426\,
                  I0 =>  \45431\,
                  I1 =>  \45428\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45428\    
  \=45427\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45427\,
                  I0 =>  \45426\,
                  I1 =>  \45342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45428\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45428\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45428\,
                   R => SYSRESET,
                   S => '0' );

  \=45428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45428\,
                  I0 =>  \45419\,
                  I1 =>  \45429\,
                  I2 =>  '0',
                  I3 => \&45427\ );

  \:45429\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45429\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45429\,
                   R => '0',
                   S => SYSRESET );

  \=45429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45429\,
                  I0 =>  \45428\,
                  I1 =>  \45419\,
                  I2 =>  \45430\,
                  I3 =>  '0' );

  \:45430\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45430\,
                   R => SYSRESET,
                   S => '0' );

  \=45430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45430\,
                  I0 =>  \45429\,
                  I1 =>  \45432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45431\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45431\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45431\,
                   R => '0',
                   S => SYSRESET );

  \=45431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45431\,
                  I0 =>  \45428\,
                  I1 =>  \45432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45432\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45432\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45432\,
                   R => SYSRESET,
                   S => '0' );

  \=45432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45432\,
                  I0 =>  \45431\,
                  I1 =>  \45429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \45434\    
  \=45433\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45433\,
                  I0 =>  \45431\,
                  I1 =>  \45425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CNTOF9\   
  \=45434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45434\,
                  I0 =>  \45418\,
                  I1 =>  \F10A\,
                  I2 =>  \45410\,
                  I3 => \&45433\ );

  -- Alias \CHOR11/\  
  \=45435\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45435\,
                  I0 =>  \CHAT11\,
                  I1 =>  \CHBT11\,
                  I2 =>  \CH1111\,
                  I3 => \&45436\ );

  -- Alias \CHOR11/\  
  \=45436\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45436\,
                  I0 =>  \CH3311\,
                  I1 =>  \CH1211\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH11\     
  \=45437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45437\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR12/\  
  \=45438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45438\,
                  I0 =>  \CHAT12\,
                  I1 =>  \CHBT12\,
                  I2 =>  '0',
                  I3 => \&45439\ );

  -- Alias \CHOR12/\  
  \=45439\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45439\,
                  I0 =>  \CH1212\,
                  I1 =>  \CH1112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH12\     
  \=45440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45440\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR13/\  
  \=45441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45441\,
                  I0 =>  \CHAT13\,
                  I1 =>  \CHBT13\,
                  I2 =>  \CH3313\,
                  I3 =>  '0' );

  -- Alias \CH13\     
  \=45442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45442\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR14/\  
  \=45443\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45443\,
                  I0 =>  \CHAT14\,
                  I1 =>  \CHBT14\,
                  I2 =>  \CH3314\,
                  I3 => \&45458\ );

  -- Alias \CH14\     
  \=45444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45444\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR16/\  
  \=45445\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45445\,
                  I0 =>  \CH1116\,
                  I1 =>  \CH1216\,
                  I2 =>  \CH3316\,
                  I3 =>  '0' );

  -- Alias \CH16\     
  \=45446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45446\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45447\,
                  I0 =>  \DKEND\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \END\      
  \=45448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45448\,
                  I0 =>  \45447\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DLKRPT\   
  \:45449\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45449\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45449\,
                   R => SYSRESET,
                   S => '0' );

  \=45449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45449\,
                  I0 =>  \45447\,
                  I1 =>  \45450\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45450\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45450\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45450\,
                   R => SYSRESET,
                   S => '0' );

  \=45450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45450\,
                  I0 =>  \45449\,
                  I1 =>  \45451\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45451\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45451\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45451\,
                   R => '0',
                   S => SYSRESET );

  \=45451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45451\,
                  I0 =>  \45449\,
                  I1 =>  \45452\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45452\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45452\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45452\,
                   R => SYSRESET,
                   S => '0' );

  \=45452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45452\,
                  I0 =>  \45451\,
                  I1 =>  \F10A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=45453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45453\,
                  I0 =>  \45447\,
                  I1 =>  \45449\,
                  I2 =>  \45451\,
                  I3 =>  '0' );

  \:45454\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \45454\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45454\,
                   R => '0',
                   S => SYSRESET );

  \=45454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45454\,
                  I0 =>  \45453\,
                  I1 =>  \45455\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:45455\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \45455\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$45455\,
                   R => SYSRESET,
                   S => '0' );

  \=45455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$45455\,
                  I0 =>  \45454\,
                  I1 =>  \CCH33\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3312\   
  \=45456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \45456\,
                  I0 =>  \45455\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR14/\  
  \=45458\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&45458\,
                  I0 =>  \CH1114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ***************************
  -- ***                     ***
  -- ***  A19/1 - INOUT IV.  ***
  -- ***                     ***
  -- ***************************

  \=46101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46101\,
                  I0 =>  \SHINC/\,
                  I1 =>  \T06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SH3MS/\   
  \:46102\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46102\,
                   R => '0',
                   S => SYSRESET );

  \=46102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46102\,
                  I0 =>  \46101\,
                  I1 =>  \46103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46103\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46103\,
                   R => SYSRESET,
                   S => '0' );

  \=46103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46103\,
                  I0 =>  \46102\,
                  I1 =>  \CSG\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46104\,
                  I0 =>  \CA6/\,
                  I1 =>  \CXB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46105\,
                  I0 =>  \46104\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46106\,
                  I0 =>  \BR1\,
                  I1 =>  \46102\,
                  I2 =>  \46105\,
                  I3 =>  '0' );

  \=46107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46107\,
                  I0 =>  \46102\,
                  I1 =>  \46105\,
                  I2 =>  \BR1/\,
                  I3 =>  '0' );

  \=46108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46108\,
                  I0 =>  \46106\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALT0\     
  \=46109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46109\,
                  I0 =>  \46108\,
                  I1 =>  \46115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALT1\     
  \=46110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46110\,
                  I0 =>  \46115\,
                  I1 =>  \46122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALRT0\    
  \=46111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46111\,
                  I0 =>  \46108\,
                  I1 =>  \46114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALRT1\    
  \=46112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46112\,
                  I0 =>  \46122\,
                  I1 =>  \46114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46113\,
                  I0 =>  \CHWL02/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46114\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46114\,
                   R => '0',
                   S => SYSRESET );

  \=46114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46114\,
                  I0 =>  \46113\,
                  I1 =>  \46115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46115\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46115\,
                   R => SYSRESET,
                   S => '0' );

  \=46115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46115\,
                  I0 =>  \46114\,
                  I1 =>  \CCH14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1402\   
  \=46116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46116\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46117\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46118\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46118\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46118\,
                   R => '0',
                   S => SYSRESET );

  \=46118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46118\,
                  I0 =>  \46117\,
                  I1 =>  \46119\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46119\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46119\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46119\,
                   R => SYSRESET,
                   S => '0' );

  \=46119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46119\,
                  I0 =>  \46118\,
                  I1 =>  \CCH14\,
                  I2 =>  \46128\,
                  I3 =>  '0' );

  -- Alias \CH1403\   
  \=46120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46120\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46121\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46121\,
                  I0 =>  \46119\,
                  I1 =>  \46128\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46122\,
                  I0 =>  \46107\,
                  I1 =>  \46126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46123\,
                  I0 =>  \46118\,
                  I1 =>  \GTSET/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46124\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46124\,
                   R => '0',
                   S => SYSRESET );

  \=46124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46124\,
                  I0 =>  \46123\,
                  I1 =>  \46125\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46125\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46125\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46125\,
                   R => SYSRESET,
                   S => '0' );

  \=46125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46125\,
                  I0 =>  \46124\,
                  I1 =>  \GOJAM\,
                  I2 =>  \GTONE\,
                  I3 =>  '0' );

  \=46126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46126\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46127\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46127\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46127\,
                   R => '0',
                   S => SYSRESET );

  \=46127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46127\,
                  I0 =>  \46126\,
                  I1 =>  \46128\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46128\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46128\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46128\,
                   R => SYSRESET,
                   S => '0' );

  \=46128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46128\,
                  I0 =>  \46127\,
                  I1 =>  \GTSET\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \ALTM\     
  \=46129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46129\,
                  I0 =>  \F5ASB0/\,
                  I1 =>  \46127\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46130\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46130\,
                   R => '0',
                   S => SYSRESET );

  \=46130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46130\,
                  I0 =>  \46128\,
                  I1 =>  \46131\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46131\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46131\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46131\,
                   R => SYSRESET,
                   S => '0' );

  \=46131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46131\,
                  I0 =>  \46130\,
                  I1 =>  \GTONE\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALTSNC\   
  \=46132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46132\,
                  I0 =>  \46133\,
                  I1 =>  \46133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46133\,
                  I0 =>  \46131\,
                  I1 =>  \46128\,
                  I2 =>  \46125\,
                  I3 =>  '0' );

  \=46134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46134\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46135\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46135\,
                   R => '0',
                   S => SYSRESET );

  \=46135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46135\,
                  I0 =>  \46134\,
                  I1 =>  \46136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46136\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46136\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46136\,
                   R => SYSRESET,
                   S => '0' );

  \=46136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46136\,
                  I0 =>  \46135\,
                  I1 =>  \CCH14\,
                  I2 =>  \46142\,
                  I3 =>  '0' );

  \=46137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46137\,
                  I0 =>  \GTSET/\,
                  I1 =>  \46135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46138\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46138\,
                   R => '0',
                   S => SYSRESET );

  \=46138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46138\,
                  I0 =>  \46137\,
                  I1 =>  \46139\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46139\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46139\,
                   R => SYSRESET,
                   S => '0' );

  \=46139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46139\,
                  I0 =>  \46138\,
                  I1 =>  \GTONE\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=46140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46140\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46141\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46141\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46141\,
                   R => '0',
                   S => SYSRESET );

  \=46141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46141\,
                  I0 =>  \46140\,
                  I1 =>  \46142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46142\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46142\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46142\,
                   R => SYSRESET,
                   S => '0' );

  \=46142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46142\,
                  I0 =>  \46141\,
                  I1 =>  \GTSET\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \OTLNKM\   
  \=46143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46143\,
                  I0 =>  \F5ASB0/\,
                  I1 =>  \46141\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46144\,
                  I0 =>  \46136\,
                  I1 =>  \46142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1401\   
  \=46145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46145\,
                  I0 =>  \46144\,
                  I1 =>  \RCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46146\,
                  I0 =>  \BR1/\,
                  I1 =>  \SH3MS/\,
                  I2 =>  \46151\,
                  I3 =>  '0' );

  -- Alias \OTLNK0\   
  \=46147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46147\,
                  I0 =>  \46151\,
                  I1 =>  \SH3MS/\,
                  I2 =>  \BR1\,
                  I3 =>  '0' );

  \=46148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46148\,
                  I0 =>  \46140\,
                  I1 =>  \46146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OTLNK1\   
  \=46149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46149\,
                  I0 =>  \46148\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46150\,
                  I0 =>  \CA5/\,
                  I1 =>  \CXB7/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46151\,
                  I0 =>  \46150\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5ASB0\   
  \=46152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46152\,
                  I0 =>  \SB0/\,
                  I1 =>  \F05A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5ASB0/\  
  \=46153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46153\,
                  I0 =>  \46152\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5ASB2\   
  \=46154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46154\,
                  I0 =>  \SB2/\,
                  I1 =>  \F05A/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5ASB2/\  
  \=46155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46155\,
                  I0 =>  \46154\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5BSB2\   
  \=46156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46156\,
                  I0 =>  \SB2/\,
                  I1 =>  \F05B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F5BSB2/\  
  \=46157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46157\,
                  I0 =>  \46156\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46158\,
                  I0 =>  \CA5/\,
                  I1 =>  \XB5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46159\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46159\,
                  I0 =>  \46158\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T2P\      
  \=46160\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46160\,
                  I0 =>  \CA2/\,
                  I1 =>  \XB5/\,
                  I2 =>  '0',
                  I3 => \&46261\ );

  \=46201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46201\,
                  I0 =>  \46225\,
                  I1 =>  \UPL0/\,
                  I2 =>  \BLKUPL\,
                  I3 =>  '0' );

  \=46202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46202\,
                  I0 =>  \46201\,
                  I1 =>  \46207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INLNKM\   
  \=46203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46203\,
                  I0 =>  \46202\,
                  I1 =>  \46227\,
                  I2 =>  \46216\,
                  I3 =>  '0' );

  \=46204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46204\,
                  I0 =>  \BLKUPL\,
                  I1 =>  \46225\,
                  I2 =>  \UPL1/\,
                  I3 =>  '0' );

  \=46205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46205\,
                  I0 =>  \46204\,
                  I1 =>  \46208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INLNKP\   
  \=46206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46206\,
                  I0 =>  \46227\,
                  I1 =>  \46205\,
                  I2 =>  \46216\,
                  I3 =>  '0' );

  \=46207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46207\,
                  I0 =>  \XLNK0/\,
                  I1 =>  \46224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46208\,
                  I0 =>  \XLNK1/\,
                  I1 =>  \46224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \46210\    
  \=46209\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&46209\,
                  I0 =>  \46201\,
                  I1 =>  \46204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46210\,
                  I0 =>  \46208\,
                  I1 =>  \46207\,
                  I2 =>  '0',
                  I3 => \&46209\ );

  \=46211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46211\,
                  I0 =>  \46210\,
                  I1 =>  \46217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH33\    
  \=46212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46212\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XT3/\,
                  I2 =>  \XB3/\,
                  I3 =>  '0' );

  \:46213\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46213\,
                   R => '0',
                   S => SYSRESET );

  \=46213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46213\,
                  I0 =>  \46211\,
                  I1 =>  \46214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46214\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46214\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46214\,
                   R => SYSRESET,
                   S => '0' );

  \=46214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46214\,
                  I0 =>  \46213\,
                  I1 =>  \46212\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  -- Alias \CH3311\   
  \=46215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46215\,
                  I0 =>  \46214\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46216\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46216\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46216\,
                   R => SYSRESET,
                   S => '0' );

  \=46216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46216\,
                  I0 =>  \46217\,
                  I1 =>  \F04A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46217\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46217\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46217\,
                   R => '0',
                   S => SYSRESET );

  \=46217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46217\,
                  I0 =>  \46219\,
                  I1 =>  \46216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46218\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46218\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46218\,
                   R => SYSRESET,
                   S => '0' );

  \=46218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46218\,
                  I0 =>  \46219\,
                  I1 =>  \46217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46219\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46219\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46219\,
                   R => SYSRESET,
                   S => '0' );

  \=46219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46219\,
                  I0 =>  \46220\,
                  I1 =>  \46218\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C45R/\    
  \=46220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46220\,
                  I0 =>  \C45R\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH3310\   
  \=46221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46221\,
                  I0 =>  \BLKUPL\,
                  I1 =>  \RCH33/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46222\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46223\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46224\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46224\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46224\,
                   R => '0',
                   S => SYSRESET );

  \=46224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46224\,
                  I0 =>  \46222\,
                  I1 =>  \46225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46225\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46225\,
                   R => SYSRESET,
                   S => '0' );

  \=46225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46225\,
                  I0 =>  \46224\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46226\,
                   R => '0',
                   S => SYSRESET );

  \=46226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46226\,
                  I0 =>  \46223\,
                  I1 =>  \46227\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46227\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46227\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46227\,
                   R => SYSRESET,
                   S => '0' );

  \=46227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46227\,
                  I0 =>  \46226\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1305\   
  \=46228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46228\,
                  I0 =>  \46224\,
                  I1 =>  \RCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1306\   
  \=46229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46229\,
                  I0 =>  \46226\,
                  I1 =>  \RCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46230\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46231\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46231\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46231\,
                   R => '0',
                   S => SYSRESET );

  \=46231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46231\,
                  I0 =>  \46230\,
                  I1 =>  \46232\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46232\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46232\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46232\,
                   R => SYSRESET,
                   S => '0' );

  \=46232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46232\,
                  I0 =>  \46231\,
                  I1 =>  \CCH14\,
                  I2 =>  \46242\,
                  I3 =>  '0' );

  -- Alias \CH1404\   
  \=46233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46233\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \THRSTD\   
  \=46234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46234\,
                  I0 =>  \46231\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46235\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46236\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46236\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46236\,
                   R => '0',
                   S => SYSRESET );

  \=46236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46236\,
                  I0 =>  \46235\,
                  I1 =>  \46237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46237\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46237\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46237\,
                   R => SYSRESET,
                   S => '0' );

  \=46237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46237\,
                  I0 =>  \46236\,
                  I1 =>  \46259\,
                  I2 =>  \CCH14\,
                  I3 =>  '0' );

  -- Alias \CH1405\   
  \=46238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46238\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EMSD\     
  \=46239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46239\,
                  I0 =>  \46236\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46240\,
                  I0 =>  \POUT/\,
                  I1 =>  \46159\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46241\,
                  I0 =>  \46159\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46242\,
                  I0 =>  \46159\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46243\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46243\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46243\,
                   R => '0',
                   S => SYSRESET );

  \=46243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46243\,
                  I0 =>  \46240\,
                  I1 =>  \46244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46244\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46244\,
                   R => SYSRESET,
                   S => '0' );

  \=46244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46244\,
                  I0 =>  \46243\,
                  I1 =>  \46231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46245\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46245\,
                   R => '0',
                   S => SYSRESET );

  \=46245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46245\,
                  I0 =>  \46241\,
                  I1 =>  \46246\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46246\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46246\,
                   R => SYSRESET,
                   S => '0' );

  \=46246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46246\,
                  I0 =>  \46245\,
                  I1 =>  \46231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \THRST+\   
  \=46247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46247\,
                  I0 =>  \46243\,
                  I1 =>  \F5ASB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \THRST-\   
  \=46248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46248\,
                  I0 =>  \F5ASB0/\,
                  I1 =>  \46245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46249\,
                  I0 =>  \CA5/\,
                  I1 =>  \XB6/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46250\,
                  I0 =>  \46249\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46251\,
                  I0 =>  \46250\,
                  I1 =>  \POUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46252\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46252\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46252\,
                   R => '0',
                   S => SYSRESET );

  \=46252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46252\,
                  I0 =>  \46251\,
                  I1 =>  \46253\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46253\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46253\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46253\,
                   R => SYSRESET,
                   S => '0' );

  \=46253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46253\,
                  I0 =>  \46252\,
                  I1 =>  \46236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EMS+\     
  \=46254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46254\,
                  I0 =>  \46252\,
                  I1 =>  \F5ASB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46255\,
                  I0 =>  \46250\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46256\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46256\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46256\,
                   R => '0',
                   S => SYSRESET );

  \=46256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46256\,
                  I0 =>  \46255\,
                  I1 =>  \46257\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46257\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46257\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46257\,
                   R => SYSRESET,
                   S => '0' );

  \=46257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46257\,
                  I0 =>  \46256\,
                  I1 =>  \46236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \EMS-\     
  \=46258\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46258\,
                  I0 =>  \46256\,
                  I1 =>  \F5ASB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46259\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46259\,
                  I0 =>  \46250\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \46160\    
  \=46261\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&46261\,
                  I0 =>  \WOVR/\,
                  I1 =>  \OVF/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ***************************
  -- ***                     ***
  -- ***  A19/2 - INOUT IV.  ***
  -- ***                     ***
  -- ***************************

  -- Alias \UPRUPT\   
  \=46303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46303\,
                  I0 =>  \BR1/\,
                  I1 =>  \C45R/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \UPL0/\    
  \=46304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46304\,
                  I0 =>  \UPL0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \UPL1/\    
  \=46305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46305\,
                  I0 =>  \UPL1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XLNK0/\   
  \=46306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46306\,
                  I0 =>  \XLNK0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \XLNK1/\   
  \=46307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46307\,
                  I0 =>  \XLNK1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BLKUPL\   
  \=46308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46308\,
                  I0 =>  \BLKUPL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F10B/\    
  \=46309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46309\,
                  I0 =>  \F10B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T1P\      
  \=46310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46310\,
                  I0 =>  \CNTRSB/\,
                  I1 =>  \46309\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T3P\      
  \=46311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46311\,
                  I0 =>  \46309\,
                  I1 =>  \CNTRSB/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F09B/\    
  \=46312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46312\,
                  I0 =>  \F09B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T4P\      
  \=46313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46313\,
                  I0 =>  \FS10\,
                  I1 =>  \46312\,
                  I2 =>  \CNTRSB/\,
                  I3 =>  '0' );

  -- Alias \F10A/\    
  \=46314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46314\,
                  I0 =>  \F10A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T5P\      
  \=46315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46315\,
                  I0 =>  \46314\,
                  I1 =>  \CNTRSB/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F06B/\    
  \=46316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46316\,
                  I0 =>  \F06B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T6P\      
  \=46317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46317\,
                  I0 =>  \CNTRSB/\,
                  I1 =>  \46316\,
                  I2 =>  \T6ON/\,
                  I3 =>  '0' );

  \=46318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46318\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46319\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46319\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46319\,
                   R => '0',
                   S => SYSRESET );

  \=46319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46319\,
                  I0 =>  \46318\,
                  I1 =>  \46320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46320\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46320\,
                   R => SYSRESET,
                   S => '0' );

  \=46320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46320\,
                  I0 =>  \46319\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1308\   
  \=46321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46321\,
                  I0 =>  \RCH13/\,
                  I1 =>  \46319\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46322\,
                  I0 =>  \46320\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46323\,
                  I0 =>  \WCH13/\,
                  I1 =>  \CHWL09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46324\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46324\,
                   R => '0',
                   S => SYSRESET );

  \=46324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46324\,
                  I0 =>  \46323\,
                  I1 =>  \46325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46325\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46325\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46325\,
                   R => SYSRESET,
                   S => '0' );

  \=46325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46325\,
                  I0 =>  \46324\,
                  I1 =>  \CCH13\,
                  I2 =>  \46330\,
                  I3 =>  '0' );

  -- Alias \CH1309\   
  \=46326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46326\,
                  I0 =>  \RCH13/\,
                  I1 =>  \46324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46327\,
                  I0 =>  \46324\,
                  I1 =>  \F07D/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46328\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46328\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46328\,
                   R => '0',
                   S => SYSRESET );

  \=46328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46328\,
                  I0 =>  \46327\,
                  I1 =>  \46329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46329\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46329\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46329\,
                   R => SYSRESET,
                   S => '0' );

  \=46329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46329\,
                  I0 =>  \46328\,
                  I1 =>  \F07B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RHCGO\    
  \=46330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46330\,
                  I0 =>  \SB2/\,
                  I1 =>  \46328\,
                  I2 =>  \F07C/\,
                  I3 =>  '0' );

  \=46331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46331\,
                  I0 =>  \46329\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46332\,
                  I0 =>  \SIGNX\,
                  I1 =>  \F7CSB1/\,
                  I2 =>  \46331\,
                  I3 =>  '0' );

  \:46333\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46333\,
                   R => '0',
                   S => SYSRESET );

  \=46333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46333\,
                  I0 =>  \46332\,
                  I1 =>  \46334\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46334\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46334\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46334\,
                   R => SYSRESET,
                   S => '0' );

  \=46334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46334\,
                  I0 =>  \46333\,
                  I1 =>  \46351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46335\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46333\,
                  I2 =>  \GATEX/\,
                  I3 =>  '0' );

  \=46336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46336\,
                  I0 =>  \GATEX/\,
                  I1 =>  \46334\,
                  I2 =>  \F5ASB2/\,
                  I3 =>  '0' );

  \=46337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46337\,
                  I0 =>  \BMGXP\,
                  I1 =>  \46335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46338\,
                  I0 =>  \46336\,
                  I1 =>  \BMGXM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGXP\   
  \=46339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46339\,
                  I0 =>  \46322\,
                  I1 =>  \46337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGXM\   
  \=46340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46340\,
                  I0 =>  \46322\,
                  I1 =>  \46338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46341\,
                  I0 =>  \SIGNY\,
                  I1 =>  \F7CSB1/\,
                  I2 =>  \46331\,
                  I3 =>  '0' );

  \:46342\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46342\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46342\,
                   R => '0',
                   S => SYSRESET );

  \=46342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46342\,
                  I0 =>  \46341\,
                  I1 =>  \46343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46343\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46343\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46343\,
                   R => SYSRESET,
                   S => '0' );

  \=46343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46343\,
                  I0 =>  \46342\,
                  I1 =>  \46351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46344\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46342\,
                  I2 =>  \GATEY/\,
                  I3 =>  '0' );

  \=46345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46345\,
                  I0 =>  \GATEY/\,
                  I1 =>  \46343\,
                  I2 =>  \F5ASB2/\,
                  I3 =>  '0' );

  \=46346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46346\,
                  I0 =>  \BMGYP\,
                  I1 =>  \46344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46347\,
                  I0 =>  \46345\,
                  I1 =>  \BMGYM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGYP\   
  \=46348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46348\,
                  I0 =>  \46322\,
                  I1 =>  \46346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGYM\   
  \=46349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46349\,
                  I0 =>  \46322\,
                  I1 =>  \46347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46350\,
                  I0 =>  \SIGNZ\,
                  I1 =>  \F7CSB1/\,
                  I2 =>  \46331\,
                  I3 =>  '0' );

  \=46351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46351\,
                  I0 =>  \46331\,
                  I1 =>  \F07C/\,
                  I2 =>  \SB0/\,
                  I3 =>  '0' );

  \:46352\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46352\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46352\,
                   R => '0',
                   S => SYSRESET );

  \=46352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46352\,
                  I0 =>  \46350\,
                  I1 =>  \46353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46353\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46353\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46353\,
                   R => SYSRESET,
                   S => '0' );

  \=46353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46353\,
                  I0 =>  \46352\,
                  I1 =>  \46351\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46354\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46352\,
                  I2 =>  \GATEZ/\,
                  I3 =>  '0' );

  \=46355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46355\,
                  I0 =>  \GATEZ/\,
                  I1 =>  \46353\,
                  I2 =>  \F5ASB2/\,
                  I3 =>  '0' );

  \=46356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46356\,
                  I0 =>  \BMGZP\,
                  I1 =>  \46354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46357\,
                  I0 =>  \46355\,
                  I1 =>  \BMGZM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGZP\   
  \=46358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46358\,
                  I0 =>  \46322\,
                  I1 =>  \46356\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BMAGZM\   
  \=46359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46359\,
                  I0 =>  \46322\,
                  I1 =>  \46357\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46401\,
                  I0 =>  \CHWL10/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46402\,
                   R => '0',
                   S => SYSRESET );

  \=46402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46402\,
                  I0 =>  \46401\,
                  I1 =>  \46403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46403\,
                   R => SYSRESET,
                   S => '0' );

  \=46403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46403\,
                  I0 =>  \46402\,
                  I1 =>  \46439\,
                  I2 =>  \CCH14\,
                  I3 =>  '0' );

  -- Alias \CH1410\   
  \=46404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46404\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46402\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYROD\    
  \=46405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46405\,
                  I0 =>  \46402\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46406\,
                  I0 =>  \CHWL09/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46407\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46407\,
                   R => '0',
                   S => SYSRESET );

  \=46407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46407\,
                  I0 =>  \46406\,
                  I1 =>  \46408\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46408\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46408\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46408\,
                   R => SYSRESET,
                   S => '0' );

  \=46408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46408\,
                  I0 =>  \46407\,
                  I1 =>  \CCH14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1409\   
  \=46409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46409\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46410\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46411\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46411\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46411\,
                   R => '0',
                   S => SYSRESET );

  \=46411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46411\,
                  I0 =>  \46410\,
                  I1 =>  \46412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46412\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46412\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46412\,
                   R => SYSRESET,
                   S => '0' );

  \=46412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46412\,
                  I0 =>  \46411\,
                  I1 =>  \CCH14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1408\   
  \=46413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46413\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46414\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46415\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46415\,
                   R => '0',
                   S => SYSRESET );

  \=46415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46415\,
                  I0 =>  \46414\,
                  I1 =>  \46416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46416\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46416\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46416\,
                   R => SYSRESET,
                   S => '0' );

  \=46416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46416\,
                  I0 =>  \46415\,
                  I1 =>  \CCH14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1407\   
  \=46417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46417\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46418\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46419\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46419\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46419\,
                   R => '0',
                   S => SYSRESET );

  \=46419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46419\,
                  I0 =>  \46418\,
                  I1 =>  \46420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46420\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46420\,
                   R => SYSRESET,
                   S => '0' );

  \=46420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46420\,
                  I0 =>  \46419\,
                  I1 =>  \CCH14\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1406\   
  \=46421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46421\,
                  I0 =>  \RCH14/\,
                  I1 =>  \46419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46422\,
                  I0 =>  \SB1/\,
                  I1 =>  \46412\,
                  I2 =>  \46415\,
                  I3 =>  '0' );

  \=46423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46423\,
                  I0 =>  \46422\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYXP\     
  \=46424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46424\,
                  I0 =>  \46408\,
                  I1 =>  \46423\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYXM\     
  \=46425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46425\,
                  I0 =>  \46423\,
                  I1 =>  \46407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYYP\     
  \=46426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46426\,
                  I0 =>  \46408\,
                  I1 =>  \46429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYYM\     
  \=46427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46427\,
                  I0 =>  \46429\,
                  I1 =>  \46407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46428\,
                  I0 =>  \SB1/\,
                  I1 =>  \46416\,
                  I2 =>  \46411\,
                  I3 =>  '0' );

  \=46429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46429\,
                  I0 =>  \46428\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46430\,
                  I0 =>  \SB1/\,
                  I1 =>  \46411\,
                  I2 =>  \46415\,
                  I3 =>  '0' );

  \=46431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46431\,
                  I0 =>  \46430\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYZP\     
  \=46432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46432\,
                  I0 =>  \46408\,
                  I1 =>  \46431\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYZM\     
  \=46433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46433\,
                  I0 =>  \46431\,
                  I1 =>  \46407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYENAB\   
  \=46434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46434\,
                  I0 =>  \SB1/\,
                  I1 =>  \46419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46435\,
                  I0 =>  \CA4/\,
                  I1 =>  \XB7/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46436\,
                  I0 =>  \46435\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46437\,
                  I0 =>  \POUT/\,
                  I1 =>  \46436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46438\,
                  I0 =>  \46436\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46439\,
                  I0 =>  \46436\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:46440\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46440\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46440\,
                   R => '0',
                   S => SYSRESET );

  \=46440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46440\,
                  I0 =>  \46441\,
                  I1 =>  \46437\,
                  I2 =>  \46438\,
                  I3 =>  '0' );

  \:46441\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46441\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46441\,
                   R => SYSRESET,
                   S => '0' );

  \=46441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46441\,
                  I0 =>  \46402\,
                  I1 =>  \46440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYRSET\   
  \=46442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46442\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GYRRST\   
  \=46443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46443\,
                  I0 =>  \F5ASB2/\,
                  I1 =>  \46441\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46444\,
                  I0 =>  \CHWL09/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1109/\  
  \:46445\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46445\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46445\,
                   R => '0',
                   S => SYSRESET );

  \=46445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46445\,
                  I0 =>  \46444\,
                  I1 =>  \46446\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1109\   
  \:46446\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46446\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46446\,
                   R => SYSRESET,
                   S => '0' );

  \=46446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46446\,
                  I0 =>  \46445\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1109\   
  \=46447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46447\,
                  I0 =>  \RCH11/\,
                  I1 =>  \46445\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \W1110\    
  \=46448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46448\,
                  I0 =>  \CHWL10/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1110/\  
  \:46449\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46449\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46449\,
                   R => '0',
                   S => SYSRESET );

  \=46449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46449\,
                  I0 =>  \46448\,
                  I1 =>  \46450\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1110\   
  \:46450\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46450\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46450\,
                   R => SYSRESET,
                   S => '0' );

  \=46450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46450\,
                  I0 =>  \46449\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1110\   
  \=46451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46451\,
                  I0 =>  \RCH11/\,
                  I1 =>  \46449\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46452\,
                  I0 =>  \CHWL11/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1111/\  
  \:46453\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46453\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46453\,
                   R => '0',
                   S => SYSRESET );

  \=46453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46453\,
                  I0 =>  \46452\,
                  I1 =>  \46454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1111\   
  \:46454\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46454\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46454\,
                   R => SYSRESET,
                   S => '0' );

  \=46454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46454\,
                  I0 =>  \46453\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1111\   
  \=46455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46455\,
                  I0 =>  \RCH11/\,
                  I1 =>  \46453\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=46456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46456\,
                  I0 =>  \CHWL12/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1112/\  
  \:46457\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \46457\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46457\,
                   R => '0',
                   S => SYSRESET );

  \=46457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46457\,
                  I0 =>  \46456\,
                  I1 =>  \46458\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FF1112\   
  \:46458\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \46458\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$46458\,
                   R => SYSRESET,
                   S => '0' );

  \=46458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$46458\,
                  I0 =>  \46457\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1112\   
  \=46459\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \46459\,
                  I0 =>  \RCH11/\,
                  I1 =>  \46457\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *********************************
  -- ***                           ***
  -- ***  A20/1 - COUNTER CELL I.  ***
  -- ***                           ***
  -- *********************************

  \=31101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31101\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31102\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31102\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31102\,
                   R => '0',
                   S => SYSRESET );

  \=31102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31102\,
                  I0 =>  \CDUXP\,
                  I1 =>  \31103\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31103\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31103\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31103\,
                   R => SYSRESET,
                   S => '0' );

  \=31103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31103\,
                  I0 =>  \31102\,
                  I1 =>  \31112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31104\,
                  I0 =>  \31103\,
                  I1 =>  \31110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31105\,
                  I0 =>  \31101\,
                  I1 =>  \31104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31106\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31106\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31106\,
                   R => '0',
                   S => SYSRESET );

  \=31106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31106\,
                  I0 =>  \31105\,
                  I1 =>  \31107\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31107\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31107\,
                   R => SYSRESET,
                   S => '0' );

  \=31107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31107\,
                  I0 =>  \31106\,
                  I1 =>  \31112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C32A\     
  \=31108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31108\,
                  I0 =>  \CG22\,
                  I1 =>  \31106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31109\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31109\,
                   R => '0',
                   S => SYSRESET );

  \=31109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31109\,
                  I0 =>  \CDUXM\,
                  I1 =>  \31110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31110\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31110\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31110\,
                   R => SYSRESET,
                   S => '0' );

  \=31110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31110\,
                  I0 =>  \31109\,
                  I1 =>  \31112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31111\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C32R\     
  \=31112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31112\,
                  I0 =>  \31111\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  -- Alias \C32P\     
  \=31113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31113\,
                  I0 =>  \31102\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  -- Alias \C32M\     
  \=31114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31114\,
                  I0 =>  \31109\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  \:31115\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31115\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31115\,
                   R => '0',
                   S => SYSRESET );

  \=31115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31115\,
                  I0 =>  \CDUYP\,
                  I1 =>  \31116\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31116\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31116\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31116\,
                   R => SYSRESET,
                   S => '0' );

  \=31116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31116\,
                  I0 =>  \31115\,
                  I1 =>  \31126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31117\,
                  I0 =>  \31116\,
                  I1 =>  \31125\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31118\,
                  I0 =>  \31101\,
                  I1 =>  \31117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31119\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31119\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31119\,
                   R => '0',
                   S => SYSRESET );

  \=31119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31119\,
                  I0 =>  \31118\,
                  I1 =>  \31120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31120\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31120\,
                   R => SYSRESET,
                   S => '0' );

  \=31120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31120\,
                  I0 =>  \31119\,
                  I1 =>  \31126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C33A\     
  \=31121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31121\,
                  I0 =>  \CG22\,
                  I1 =>  \31107\,
                  I2 =>  \31119\,
                  I3 =>  '0' );

  \=31122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31122\,
                  I0 =>  \CG22\,
                  I1 =>  \31120\,
                  I2 =>  \31107\,
                  I3 =>  '0' );

  -- Alias \CG11\     
  \=31123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31123\,
                  I0 =>  \31122\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31124\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31124\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31124\,
                   R => '0',
                   S => SYSRESET );

  \=31124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31124\,
                  I0 =>  \CDUYM\,
                  I1 =>  \31125\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31125\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31125\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31125\,
                   R => SYSRESET,
                   S => '0' );

  \=31125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31125\,
                  I0 =>  \31124\,
                  I1 =>  \31126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C33R\     
  \=31126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31126\,
                  I0 =>  \31111\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  -- Alias \C33P\     
  \=31127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31127\,
                  I0 =>  \31115\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  -- Alias \C33M\     
  \=31128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31128\,
                  I0 =>  \31124\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  \:31129\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31129\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31129\,
                   R => '0',
                   S => SYSRESET );

  \=31129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31129\,
                  I0 =>  \T2P\,
                  I1 =>  \31130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31130\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31130\,
                   R => SYSRESET,
                   S => '0' );

  \=31130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31130\,
                  I0 =>  \31129\,
                  I1 =>  \31135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31131\,
                  I0 =>  \31101\,
                  I1 =>  \31129\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31132\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31132\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31132\,
                   R => '0',
                   S => SYSRESET );

  \=31132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31132\,
                  I0 =>  \31131\,
                  I1 =>  \31133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31133\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31133\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31133\,
                   R => SYSRESET,
                   S => '0' );

  \=31133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31133\,
                  I0 =>  \31132\,
                  I1 =>  \31135\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C24A\     
  \=31134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31134\,
                  I0 =>  \31132\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C24R\     
  \=31135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31135\,
                  I0 =>  \31111\,
                  I1 =>  \CA2/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  \:31136\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31136\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31136\,
                   R => '0',
                   S => SYSRESET );

  \=31136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31136\,
                  I0 =>  \T1P\,
                  I1 =>  \31137\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31137\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31137\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31137\,
                   R => SYSRESET,
                   S => '0' );

  \=31137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31137\,
                  I0 =>  \31136\,
                  I1 =>  \31142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31138\,
                  I0 =>  \31101\,
                  I1 =>  \31136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31139\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31139\,
                   R => '0',
                   S => SYSRESET );

  \=31139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31139\,
                  I0 =>  \31138\,
                  I1 =>  \31140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31140\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31140\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31140\,
                   R => SYSRESET,
                   S => '0' );

  \=31140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31140\,
                  I0 =>  \31139\,
                  I1 =>  \31142\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C25A\     
  \=31141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31141\,
                  I0 =>  '0',
                  I1 =>  \31139\,
                  I2 =>  \31133\,
                  I3 =>  '0' );

  -- Alias \C25R\     
  \=31142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31142\,
                  I0 =>  \31111\,
                  I1 =>  \CA2/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  \:31143\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31143\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31143\,
                   R => '0',
                   S => SYSRESET );

  \=31143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31143\,
                  I0 =>  \T3P\,
                  I1 =>  \31144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31144\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31144\,
                   R => SYSRESET,
                   S => '0' );

  \=31144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31144\,
                  I0 =>  \31143\,
                  I1 =>  \31153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31145\,
                  I0 =>  \31101\,
                  I1 =>  \31143\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31146\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31146\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31146\,
                   R => '0',
                   S => SYSRESET );

  \=31146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31146\,
                  I0 =>  \31145\,
                  I1 =>  \31147\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31147\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31147\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31147\,
                   R => SYSRESET,
                   S => '0' );

  \=31147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31147\,
                  I0 =>  \31146\,
                  I1 =>  \31153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \31149\    
  \=31148\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31148\,
                  I0 =>  '0',
                  I1 =>  \31133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C26A\     
  \=31149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31149\,
                  I0 =>  \31140\,
                  I1 =>  \31146\,
                  I2 =>  '0',
                  I3 => \&31148\ );

  \=31150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31150\,
                  I0 =>  '0',
                  I1 =>  \31133\,
                  I2 =>  '0',
                  I3 => \&31151\ );

  -- Alias \31150\    
  \=31151\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31151\,
                  I0 =>  \31140\,
                  I1 =>  \31147\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CG21\     
  \=31152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31152\,
                  I0 =>  \31150\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C26R\     
  \=31153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31153\,
                  I0 =>  \31111\,
                  I1 =>  \CA2/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  -- Alias \CA3/\     
  \=31154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31154\,
                  I0 =>  \OCTAD3\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CXB7/\    
  \=31158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31158\,
                  I0 =>  \XB7\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31201\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31202\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31202\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31202\,
                   R => '0',
                   S => SYSRESET );

  \=31202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31202\,
                  I0 =>  \CDUZP\,
                  I1 =>  \31203\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31203\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31203\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31203\,
                   R => SYSRESET,
                   S => '0' );

  \=31203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31203\,
                  I0 =>  \31202\,
                  I1 =>  \31212\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31204\,
                  I0 =>  \31203\,
                  I1 =>  \31210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31205\,
                  I0 =>  \31201\,
                  I1 =>  \31204\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31206\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31206\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31206\,
                   R => '0',
                   S => SYSRESET );

  \=31206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31206\,
                  I0 =>  \31205\,
                  I1 =>  \31207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31207\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31207\,
                   R => SYSRESET,
                   S => '0' );

  \=31207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31207\,
                  I0 =>  \31206\,
                  I1 =>  \31212\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C34A\     
  \=31208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31208\,
                  I0 =>  \CG11\,
                  I1 =>  \31206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31209\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31209\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31209\,
                   R => '0',
                   S => SYSRESET );

  \=31209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31209\,
                  I0 =>  \CDUZM\,
                  I1 =>  \31210\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31210\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31210\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31210\,
                   R => SYSRESET,
                   S => '0' );

  \=31210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31210\,
                  I0 =>  \31209\,
                  I1 =>  \31212\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31211\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C34R\     
  \=31212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31212\,
                  I0 =>  \31211\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  -- Alias \C34P\     
  \=31213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31213\,
                  I0 =>  \31202\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  -- Alias \C34M\     
  \=31214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31214\,
                  I0 =>  \31209\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  \:31215\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31215\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31215\,
                   R => '0',
                   S => SYSRESET );

  \=31215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31215\,
                  I0 =>  \TRNP\,
                  I1 =>  \31216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31216\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31216\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31216\,
                   R => SYSRESET,
                   S => '0' );

  \=31216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31216\,
                  I0 =>  \31215\,
                  I1 =>  \31226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31217\,
                  I0 =>  \31216\,
                  I1 =>  \31225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31218\,
                  I0 =>  \31201\,
                  I1 =>  \31217\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31219\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31219\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31219\,
                   R => '0',
                   S => SYSRESET );

  \=31219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31219\,
                  I0 =>  \31218\,
                  I1 =>  \31220\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31220\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31220\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31220\,
                   R => SYSRESET,
                   S => '0' );

  \=31220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31220\,
                  I0 =>  \31219\,
                  I1 =>  \31226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C35A\     
  \=31221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31221\,
                  I0 =>  \CG11\,
                  I1 =>  \31207\,
                  I2 =>  \31219\,
                  I3 =>  '0' );

  \=31222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31222\,
                  I0 =>  \CG11\,
                  I1 =>  \31220\,
                  I2 =>  \31207\,
                  I3 =>  '0' );

  -- Alias \CG12\     
  \=31223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31223\,
                  I0 =>  \31222\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31224\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31224\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31224\,
                   R => '0',
                   S => SYSRESET );

  \=31224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31224\,
                  I0 =>  \TRNM\,
                  I1 =>  \31225\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31225\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31225\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31225\,
                   R => SYSRESET,
                   S => '0' );

  \=31225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31225\,
                  I0 =>  \31224\,
                  I1 =>  \31226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C35R\     
  \=31226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31226\,
                  I0 =>  \31211\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  -- Alias \C35P\     
  \=31227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31227\,
                  I0 =>  \31215\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  -- Alias \C35M\     
  \=31228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31228\,
                  I0 =>  \31224\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  \:31229\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31229\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31229\,
                   R => '0',
                   S => SYSRESET );

  \=31229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31229\,
                  I0 =>  \T4P\,
                  I1 =>  \31230\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31230\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31230\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31230\,
                   R => SYSRESET,
                   S => '0' );

  \=31230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31230\,
                  I0 =>  \31229\,
                  I1 =>  \31235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31231\,
                  I0 =>  \31201\,
                  I1 =>  \31229\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31232\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31232\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31232\,
                   R => '0',
                   S => SYSRESET );

  \=31232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31232\,
                  I0 =>  \31231\,
                  I1 =>  \31233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31233\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31233\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31233\,
                   R => SYSRESET,
                   S => '0' );

  \=31233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31233\,
                  I0 =>  \31232\,
                  I1 =>  \31235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C27A\     
  \=31234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31234\,
                  I0 =>  \31232\,
                  I1 =>  \CG21\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C27R\     
  \=31235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31235\,
                  I0 =>  \31211\,
                  I1 =>  \CA2/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  \:31236\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31236\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31236\,
                   R => '0',
                   S => SYSRESET );

  \=31236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31236\,
                  I0 =>  \T5P\,
                  I1 =>  \31237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31237\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31237\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31237\,
                   R => SYSRESET,
                   S => '0' );

  \=31237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31237\,
                  I0 =>  \31236\,
                  I1 =>  \31242\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31238\,
                  I0 =>  \31201\,
                  I1 =>  \31236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31239\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31239\,
                   R => '0',
                   S => SYSRESET );

  \=31239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31239\,
                  I0 =>  \31238\,
                  I1 =>  \31240\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31240\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31240\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31240\,
                   R => SYSRESET,
                   S => '0' );

  \=31240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31240\,
                  I0 =>  \31239\,
                  I1 =>  \31242\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C30A\     
  \=31241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31241\,
                  I0 =>  \CG21\,
                  I1 =>  \31239\,
                  I2 =>  \31233\,
                  I3 =>  '0' );

  -- Alias \C30R\     
  \=31242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31242\,
                  I0 =>  \31211\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  \:31243\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31243\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31243\,
                   R => '0',
                   S => SYSRESET );

  \=31243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31243\,
                  I0 =>  \T6P\,
                  I1 =>  \31244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31244\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31244\,
                   R => SYSRESET,
                   S => '0' );

  \=31244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31244\,
                  I0 =>  \31243\,
                  I1 =>  \31253\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31245\,
                  I0 =>  \31201\,
                  I1 =>  \31243\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31246\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31246\,
                   R => '0',
                   S => SYSRESET );

  \=31246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31246\,
                  I0 =>  \31245\,
                  I1 =>  \31247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31247\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31247\,
                   R => SYSRESET,
                   S => '0' );

  \=31247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31247\,
                  I0 =>  \31246\,
                  I1 =>  \31253\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \31249\    
  \=31248\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31248\,
                  I0 =>  \CG21\,
                  I1 =>  \31233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C31A\     
  \=31249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31249\,
                  I0 =>  \31240\,
                  I1 =>  \31246\,
                  I2 =>  '0',
                  I3 => \&31248\ );

  \=31250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31250\,
                  I0 =>  \CG21\,
                  I1 =>  \31233\,
                  I2 =>  '0',
                  I3 => \&31251\ );

  -- Alias \31250\    
  \=31251\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31251\,
                  I0 =>  \31240\,
                  I1 =>  \31247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CG22\     
  \=31252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31252\,
                  I0 =>  \31250\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C31R\     
  \=31253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31253\,
                  I0 =>  \31211\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB1/\,
                  I3 =>  '0' );

  -- Alias \CXB2/\    
  \=31256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31256\,
                  I0 =>  \XB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- *********************************
  -- ***                           ***
  -- ***  A20/2 - COUNTER CELL I.  ***
  -- ***                           ***
  -- *********************************

  \=31301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31301\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31302\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31302\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31302\,
                   R => '0',
                   S => SYSRESET );

  \=31302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31302\,
                  I0 =>  \SHAFTP\,
                  I1 =>  \31303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31303\,
                   R => SYSRESET,
                   S => '0' );

  \=31303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31303\,
                  I0 =>  \31302\,
                  I1 =>  \31312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31304\,
                  I0 =>  \31303\,
                  I1 =>  \31310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31305\,
                  I0 =>  \31301\,
                  I1 =>  \31304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31306\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31306\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31306\,
                   R => '0',
                   S => SYSRESET );

  \=31306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31306\,
                  I0 =>  \31305\,
                  I1 =>  \31307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31307\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31307\,
                   R => SYSRESET,
                   S => '0' );

  \=31307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31307\,
                  I0 =>  \31306\,
                  I1 =>  \31312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C36A\     
  \=31308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31308\,
                  I0 =>  \CG12\,
                  I1 =>  \31306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31309\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31309\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31309\,
                   R => '0',
                   S => SYSRESET );

  \=31309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31309\,
                  I0 =>  \SHAFTM\,
                  I1 =>  \31310\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31310\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31310\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31310\,
                   R => SYSRESET,
                   S => '0' );

  \=31310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31310\,
                  I0 =>  \31309\,
                  I1 =>  \31312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31311\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C36R\     
  \=31312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31312\,
                  I0 =>  \31311\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  -- Alias \C36P\     
  \=31313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31313\,
                  I0 =>  \31302\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  -- Alias \C36M\     
  \=31314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31314\,
                  I0 =>  \31309\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  \:31315\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31315\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31315\,
                   R => '0',
                   S => SYSRESET );

  \=31315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31315\,
                  I0 =>  \PIPXP\,
                  I1 =>  \31316\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31316\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31316\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31316\,
                   R => SYSRESET,
                   S => '0' );

  \=31316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31316\,
                  I0 =>  \31315\,
                  I1 =>  \31326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31317\,
                  I0 =>  \31316\,
                  I1 =>  \31325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31318\,
                  I0 =>  \31301\,
                  I1 =>  \31317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31319\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31319\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31319\,
                   R => '0',
                   S => SYSRESET );

  \=31319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31319\,
                  I0 =>  \31318\,
                  I1 =>  \31320\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31320\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31320\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31320\,
                   R => SYSRESET,
                   S => '0' );

  \=31320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31320\,
                  I0 =>  \31319\,
                  I1 =>  \31326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C37A\     
  \=31321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31321\,
                  I0 =>  \CG12\,
                  I1 =>  \31307\,
                  I2 =>  \31319\,
                  I3 =>  '0' );

  \=31322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31322\,
                  I0 =>  \CG12\,
                  I1 =>  \31320\,
                  I2 =>  \31307\,
                  I3 =>  '0' );

  -- Alias \CG14\     
  \=31323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31323\,
                  I0 =>  \31322\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31324\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31324\,
                   R => '0',
                   S => SYSRESET );

  \=31324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31324\,
                  I0 =>  \PIPXM\,
                  I1 =>  \31325\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31325\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31325\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31325\,
                   R => SYSRESET,
                   S => '0' );

  \=31325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31325\,
                  I0 =>  \31324\,
                  I1 =>  \31326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C37R\     
  \=31326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31326\,
                  I0 =>  \31311\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  -- Alias \C37P\     
  \=31327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31327\,
                  I0 =>  \31315\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  -- Alias \C37M\     
  \=31328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31328\,
                  I0 =>  \31324\,
                  I1 =>  \CA3/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  \:31329\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31329\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31329\,
                   R => '0',
                   S => SYSRESET );

  \=31329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31329\,
                  I0 =>  \CDUXD\,
                  I1 =>  \31330\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31330\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31330\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31330\,
                   R => SYSRESET,
                   S => '0' );

  \=31330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31330\,
                  I0 =>  \31329\,
                  I1 =>  \31335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31331\,
                  I0 =>  \31301\,
                  I1 =>  \31329\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31332\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31332\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31332\,
                   R => '0',
                   S => SYSRESET );

  \=31332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31332\,
                  I0 =>  \31331\,
                  I1 =>  \31333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31333\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31333\,
                   R => SYSRESET,
                   S => '0' );

  \=31333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31333\,
                  I0 =>  \31332\,
                  I1 =>  \31335\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C50A\     
  \=31334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31334\,
                  I0 =>  \31332\,
                  I1 =>  \CG26\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C50R\     
  \=31335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31335\,
                  I0 =>  \31311\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  \:31336\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31336\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31336\,
                   R => '0',
                   S => SYSRESET );

  \=31336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31336\,
                  I0 =>  \CDUYD\,
                  I1 =>  \31337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31337\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31337\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31337\,
                   R => SYSRESET,
                   S => '0' );

  \=31337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31337\,
                  I0 =>  \31336\,
                  I1 =>  \31342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31338\,
                  I0 =>  \31301\,
                  I1 =>  \31336\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31339\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31339\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31339\,
                   R => '0',
                   S => SYSRESET );

  \=31339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31339\,
                  I0 =>  \31338\,
                  I1 =>  \31340\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31340\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31340\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31340\,
                   R => SYSRESET,
                   S => '0' );

  \=31340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31340\,
                  I0 =>  \31339\,
                  I1 =>  \31342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C51A\     
  \=31341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31341\,
                  I0 =>  \CG26\,
                  I1 =>  \31339\,
                  I2 =>  \31333\,
                  I3 =>  '0' );

  -- Alias \C51R\     
  \=31342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31342\,
                  I0 =>  \31311\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB1/\,
                  I3 =>  '0' );

  \:31343\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31343\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31343\,
                   R => '0',
                   S => SYSRESET );

  \=31343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31343\,
                  I0 =>  \CDUZD\,
                  I1 =>  \31344\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31344\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31344\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31344\,
                   R => SYSRESET,
                   S => '0' );

  \=31344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31344\,
                  I0 =>  \31343\,
                  I1 =>  \31353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31345\,
                  I0 =>  \31301\,
                  I1 =>  \31343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31346\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31346\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31346\,
                   R => '0',
                   S => SYSRESET );

  \=31346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31346\,
                  I0 =>  \31345\,
                  I1 =>  \31347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31347\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31347\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31347\,
                   R => SYSRESET,
                   S => '0' );

  \=31347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31347\,
                  I0 =>  \31346\,
                  I1 =>  \31353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \31349\    
  \=31348\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31348\,
                  I0 =>  \CG26\,
                  I1 =>  \31333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C52A\     
  \=31349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31349\,
                  I0 =>  \31340\,
                  I1 =>  \31346\,
                  I2 =>  '0',
                  I3 => \&31348\ );

  \=31350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31350\,
                  I0 =>  \CG26\,
                  I1 =>  \31333\,
                  I2 =>  '0',
                  I3 => \&31351\ );

  -- Alias \31350\    
  \=31351\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31351\,
                  I0 =>  \31340\,
                  I1 =>  \31347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CG24\     
  \=31352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31352\,
                  I0 =>  \31350\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C52R\     
  \=31353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31353\,
                  I0 =>  \31311\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  -- Alias \CA4/\     
  \=31354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31354\,
                  I0 =>  \OCTAD4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CXB3/\    
  \=31356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31356\,
                  I0 =>  \XB3\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CA2/\     
  \=31358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31358\,
                  I0 =>  \OCTAD2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31401\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31402\,
                   R => '0',
                   S => SYSRESET );

  \=31402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31402\,
                  I0 =>  \PIPYP\,
                  I1 =>  \31403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31403\,
                   R => SYSRESET,
                   S => '0' );

  \=31403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31403\,
                  I0 =>  \31402\,
                  I1 =>  \31412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31404\,
                  I0 =>  \31403\,
                  I1 =>  \31410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31405\,
                  I0 =>  \31401\,
                  I1 =>  \31404\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31406\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31406\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31406\,
                   R => '0',
                   S => SYSRESET );

  \=31406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31406\,
                  I0 =>  \31405\,
                  I1 =>  \31407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31407\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31407\,
                   R => SYSRESET,
                   S => '0' );

  \=31407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31407\,
                  I0 =>  \31406\,
                  I1 =>  \31412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C40A\     
  \=31408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31408\,
                  I0 =>  \CG14\,
                  I1 =>  \31406\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31409\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31409\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31409\,
                   R => '0',
                   S => SYSRESET );

  \=31409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31409\,
                  I0 =>  \PIPYM\,
                  I1 =>  \31410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31410\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31410\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31410\,
                   R => SYSRESET,
                   S => '0' );

  \=31410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31410\,
                  I0 =>  \31409\,
                  I1 =>  \31412\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31411\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C40R\     
  \=31412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31412\,
                  I0 =>  \31411\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  -- Alias \C40P\     
  \=31413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31413\,
                  I0 =>  \31402\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  -- Alias \C40M\     
  \=31414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31414\,
                  I0 =>  \31409\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  \:31415\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31415\,
                   R => '0',
                   S => SYSRESET );

  \=31415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31415\,
                  I0 =>  \PIPZP\,
                  I1 =>  \31416\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31416\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31416\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31416\,
                   R => SYSRESET,
                   S => '0' );

  \=31416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31416\,
                  I0 =>  \31415\,
                  I1 =>  \31426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31417\,
                  I0 =>  \31416\,
                  I1 =>  \31425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31418\,
                  I0 =>  \31401\,
                  I1 =>  \31417\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31419\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31419\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31419\,
                   R => '0',
                   S => SYSRESET );

  \=31419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31419\,
                  I0 =>  \31418\,
                  I1 =>  \31420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31420\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31420\,
                   R => SYSRESET,
                   S => '0' );

  \=31420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31420\,
                  I0 =>  \31419\,
                  I1 =>  \31426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C41A\     
  \=31421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31421\,
                  I0 =>  \CG14\,
                  I1 =>  \31407\,
                  I2 =>  \31419\,
                  I3 =>  '0' );

  \=31422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31422\,
                  I0 =>  \CG14\,
                  I1 =>  \31420\,
                  I2 =>  \31407\,
                  I3 =>  '0' );

  -- Alias \CG13\     
  \=31423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31423\,
                  I0 =>  \31422\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31424\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31424\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31424\,
                   R => '0',
                   S => SYSRESET );

  \=31424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31424\,
                  I0 =>  \PIPZM\,
                  I1 =>  \31425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31425\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31425\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31425\,
                   R => SYSRESET,
                   S => '0' );

  \=31425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31425\,
                  I0 =>  \31424\,
                  I1 =>  \31426\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C41R\     
  \=31426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31426\,
                  I0 =>  \31411\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB1/\,
                  I3 =>  '0' );

  -- Alias \C41P\     
  \=31427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31427\,
                  I0 =>  \31415\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB1/\,
                  I3 =>  '0' );

  -- Alias \C41M\     
  \=31428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31428\,
                  I0 =>  \31424\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB1/\,
                  I3 =>  '0' );

  \:31429\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31429\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31429\,
                   R => '0',
                   S => SYSRESET );

  \=31429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31429\,
                  I0 =>  \TRUND\,
                  I1 =>  \31430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31430\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31430\,
                   R => SYSRESET,
                   S => '0' );

  \=31430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31430\,
                  I0 =>  \31429\,
                  I1 =>  \31435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31431\,
                  I0 =>  \31401\,
                  I1 =>  \31429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31432\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31432\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31432\,
                   R => '0',
                   S => SYSRESET );

  \=31432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31432\,
                  I0 =>  \31431\,
                  I1 =>  \31433\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31433\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31433\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31433\,
                   R => SYSRESET,
                   S => '0' );

  \=31433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31433\,
                  I0 =>  \31432\,
                  I1 =>  \31435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C53A\     
  \=31434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31434\,
                  I0 =>  \31432\,
                  I1 =>  \CG24\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C53R\     
  \=31435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31435\,
                  I0 =>  \31411\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  \:31436\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31436\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31436\,
                   R => '0',
                   S => SYSRESET );

  \=31436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31436\,
                  I0 =>  \SHAFTD\,
                  I1 =>  \31437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31437\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31437\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31437\,
                   R => SYSRESET,
                   S => '0' );

  \=31437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31437\,
                  I0 =>  \31436\,
                  I1 =>  \31442\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31438\,
                  I0 =>  \31401\,
                  I1 =>  \31436\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31439\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31439\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31439\,
                   R => '0',
                   S => SYSRESET );

  \=31439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31439\,
                  I0 =>  \31438\,
                  I1 =>  \31440\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31440\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31440\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31440\,
                   R => SYSRESET,
                   S => '0' );

  \=31440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31440\,
                  I0 =>  \31439\,
                  I1 =>  \31442\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C54A\     
  \=31441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31441\,
                  I0 =>  \CG24\,
                  I1 =>  \31439\,
                  I2 =>  \31433\,
                  I3 =>  '0' );

  -- Alias \C54R\     
  \=31442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31442\,
                  I0 =>  \31411\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  \:31443\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31443\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31443\,
                   R => '0',
                   S => SYSRESET );

  \=31443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31443\,
                  I0 =>  \THRSTD\,
                  I1 =>  \31444\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31444\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31444\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31444\,
                   R => SYSRESET,
                   S => '0' );

  \=31444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31444\,
                  I0 =>  \31443\,
                  I1 =>  \31453\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=31445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31445\,
                  I0 =>  \31401\,
                  I1 =>  \31443\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31446\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \31446\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31446\,
                   R => '0',
                   S => SYSRESET );

  \=31446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31446\,
                  I0 =>  \31445\,
                  I1 =>  \31447\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:31447\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \31447\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$31447\,
                   R => SYSRESET,
                   S => '0' );

  \=31447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$31447\,
                  I0 =>  \31446\,
                  I1 =>  \31453\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \31449\    
  \=31448\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31448\,
                  I0 =>  \CG24\,
                  I1 =>  \31433\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C55A\     
  \=31449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31449\,
                  I0 =>  \31440\,
                  I1 =>  \31446\,
                  I2 =>  '0',
                  I3 => \&31448\ );

  \=31450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31450\,
                  I0 =>  \CG24\,
                  I1 =>  \31433\,
                  I2 =>  '0',
                  I3 => \&31451\ );

  -- Alias \31450\    
  \=31451\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&31451\,
                  I0 =>  \31440\,
                  I1 =>  \31447\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CG23\     
  \=31452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31452\,
                  I0 =>  \31450\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C55R\     
  \=31453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31453\,
                  I0 =>  \31411\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  -- Alias \CXB4/\    
  \=31456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31456\,
                  I0 =>  \XB4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CA6/\     
  \=31458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \31458\,
                  I0 =>  \OCTAD6\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- **********************************
  -- ***                            ***
  -- ***  A21/1 - COUNTER CELL II.  ***
  -- ***                            ***
  -- **********************************

  -- Alias \32021\    
  \=32001\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32001\,
                  I0 =>  \C25A\,
                  I1 =>  \C27A\,
                  I2 =>  \C31A\,
                  I3 => \&32011\ );

  -- Alias \32022\    
  \=32002\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32002\,
                  I0 =>  \C26A\,
                  I1 =>  \C27A\,
                  I2 =>  \C32A\,
                  I3 => \&32012\ );

  -- Alias \32033\    
  \=32003\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32003\,
                  I0 =>  \C24A\,
                  I1 =>  \C25A\,
                  I2 =>  \C26A\,
                  I3 => \&32013\ );

  -- Alias \32014\    
  \=32004\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32004\,
                  I0 =>  \C30A\,
                  I1 =>  \C31A\,
                  I2 =>  \C32A\,
                  I3 => \&32024\ );

  -- Alias \32015\    
  \=32005\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32005\,
                  I0 =>  \C24A\,
                  I1 =>  \C25A\,
                  I2 =>  \C26A\,
                  I3 =>  '0' );

  -- Alias \32016\    
  \=32006\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32006\,
                  I0 =>  \C40A\,
                  I1 =>  \C41A\,
                  I2 =>  \C42A\,
                  I3 => \&32026\ );

  \=32007\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32007\,
                  I0 =>  \32064\,
                  I1 =>  \32050\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CAD4\     
  \=32008\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32008\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32007\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32021\    
  \=32011\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32011\,
                  I0 =>  \C33A\,
                  I1 =>  \C35A\,
                  I2 =>  \C37A\,
                  I3 => \&32031\ );

  -- Alias \32022\    
  \=32012\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32012\,
                  I0 =>  \C33A\,
                  I1 =>  \C36A\,
                  I2 =>  \C37A\,
                  I3 => \&32032\ );

  -- Alias \32033\    
  \=32013\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32013\,
                  I0 =>  \C27A\,
                  I1 =>  \C34A\,
                  I2 =>  \C35A\,
                  I3 => \&32023\ );

  -- Alias \32004K?\  
  \=32014\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32014\,
                  I0 =>  \C33A\,
                  I1 =>  \C34A\,
                  I2 =>  \C35A\,
                  I3 => \&32004\ );

  \=32015\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32015\,
                  I0 =>  \C27A\,
                  I1 =>  \32064\,
                  I2 =>  \C60A\,
                  I3 => \&32005\ );

  \=32016\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32016\,
                  I0 =>  \C43A\,
                  I1 =>  \C44A\,
                  I2 =>  \C45A\,
                  I3 => \&32006\ );

  \=32021\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32021\,
                  I0 =>  \C41A\,
                  I1 =>  \C43A\,
                  I2 =>  \C45A\,
                  I3 => \&32001\ );

  \=32022\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32022\,
                  I0 =>  \C42A\,
                  I1 =>  \C43A\,
                  I2 =>  \C46A\,
                  I3 => \&32002\ );

  -- Alias \32033\    
  \=32023\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32023\,
                  I0 =>  \C36A\,
                  I1 =>  \C37A\,
                  I2 =>  \C44A\,
                  I3 => \&32043\ );

  -- Alias \32014\    
  \=32024\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32024\,
                  I0 =>  \C36A\,
                  I1 =>  \C37A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32016\    
  \=32026\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32026\,
                  I0 =>  \C46A\,
                  I1 =>  \C47A\,
                  I2 =>  \32050\,
                  I3 => \&32036\ );

  -- Alias \32021\    
  \=32031\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32031\,
                  I0 =>  \C47A\,
                  I1 =>  \C51A\,
                  I2 =>  \C53A\,
                  I3 => \&32041\ );

  -- Alias \32022\    
  \=32032\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32032\,
                  I0 =>  \C47A\,
                  I1 =>  \C52A\,
                  I2 =>  \C53A\,
                  I3 => \&32042\ );

  \=32033\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32033\,
                  I0 =>  \C45A\,
                  I1 =>  \C46A\,
                  I2 =>  \C47A\,
                  I3 => \&32003\ );

  -- Alias \32044\    
  \=32034\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32034\,
                  I0 =>  \C50A\,
                  I1 =>  \C51A\,
                  I2 =>  \C52A\,
                  I3 => \&32054\ );

  -- Alias \CAD5\     
  \=32035\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32035\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32015\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32016\    
  \=32036\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32036\,
                  I0 =>  \C60A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32021\    
  \=32041\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32041\,
                  I0 =>  \C55A\,
                  I1 =>  \C57A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32022\    
  \=32042\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32042\,
                  I0 =>  \C56A\,
                  I1 =>  \C57A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32033\    
  \=32043\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32043\,
                  I0 =>  \C54A\,
                  I1 =>  \C55A\,
                  I2 =>  \C56A\,
                  I3 => \&32053\ );

  \=32044\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32044\,
                  I0 =>  \C53A\,
                  I1 =>  \C54A\,
                  I2 =>  \C55A\,
                  I3 => \&32034\ );

  -- Alias \DINC/\    
  \=32045\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32045\,
                  I0 =>  \DINC\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CAD6\     
  \=32046\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32046\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32016\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DINC\     
  \=32047\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32047\,
                  I0 =>  \32048\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DINCNC/\  
  \:32048\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32048\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32048\,
                   R => '0',
                   S => SYSRESET );

  \=32048\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32048\,
                  I0 =>  \32049\,
                  I1 =>  \32047\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32049\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32049\,
                  I0 =>  \INCSET/\,
                  I1 =>  \32068\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \50SUM\    
  \=32050\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32050\,
                  I0 =>  \32044\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CAD1\     
  \=32051\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32051\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32021\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CAD2\     
  \=32052\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32052\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32022\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32033\    
  \=32053\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32053\,
                  I0 =>  \C57A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32044\    
  \=32054\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32054\,
                  I0 =>  \C56A\,
                  I1 =>  \C57A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32056\    
  \=32055\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32055\,
                  I0 =>  \C45M\,
                  I1 =>  \C46M\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32056\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32056\,
                  I0 =>  \C57A\,
                  I1 =>  \C60A\,
                  I2 =>  '0',
                  I3 => \&32055\ );

  \=32058\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32058\,
                  I0 =>  \INCSET/\,
                  I1 =>  \32056\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHINC/\   
  \:32059\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32059\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32059\,
                   R => '0',
                   S => SYSRESET );

  \=32059\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32059\,
                  I0 =>  \32058\,
                  I1 =>  \32060\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHINC\    
  \=32060\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32060\,
                  I0 =>  \32059\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32061\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32061\,
                  I0 =>  \C45P\,
                  I1 =>  \C46P\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32062\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32062\,
                  I0 =>  \INCSET/\,
                  I1 =>  \32061\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CAD3\     
  \=32063\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32063\,
                  I0 =>  \RSCT/\,
                  I1 =>  \32033\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \30SUM\    
  \=32064\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32064\,
                  I0 =>  \32004K?\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHANC/\   
  \:32065\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32065\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32065\,
                   R => '0',
                   S => SYSRESET );

  \=32065\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32065\,
                  I0 =>  \32062\,
                  I1 =>  \32066\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHANC\    
  \=32066\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32066\,
                  I0 =>  \32065\,
                  I1 =>  \T12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32068\    
  \=32067\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32067\,
                  I0 =>  \C31A\,
                  I1 =>  \C47A\,
                  I2 =>  \C50A\,
                  I3 => \&32069\ );

  \=32068\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32068\,
                  I0 =>  \C51A\,
                  I1 =>  \C52A\,
                  I2 =>  \C53A\,
                  I3 => \&32067\ );

  -- Alias \32068\    
  \=32069\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32069\,
                  I0 =>  \C54A\,
                  I1 =>  \C55A\,
                  I2 =>  \C56A\,
                  I3 =>  '0' );

  -- **********************************
  -- ***                            ***
  -- ***  A21/2 - COUNTER CELL II.  ***
  -- ***                            ***
  -- **********************************

  -- Alias \32202\    
  \=32201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32201\,
                  I0 =>  \T12/\,
                  I1 =>  \PHS4/\,
                  I2 =>  \NISQL/\,
                  I3 =>  '0' );

  \=32202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32202\,
                  I0 =>  \GNHNC\,
                  I1 =>  \PSEUDO\,
                  I2 =>  '0',
                  I3 => \&32201\ );

  \=32203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32203\,
                  I0 =>  \32202\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32204\,
                  I0 =>  \MLOAD\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32205\,
                  I0 =>  \32203\,
                  I1 =>  \32204\,
                  I2 =>  \32238\,
                  I3 =>  '0' );

  \:32206\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32206\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32206\,
                   R => '0',
                   S => SYSRESET );

  \=32206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32206\,
                  I0 =>  \32205\,
                  I1 =>  \32207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32207\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32207\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32207\,
                   R => SYSRESET,
                   S => '0' );

  \=32207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32207\,
                  I0 =>  \32206\,
                  I1 =>  \GOJAM\,
                  I2 =>  \32218\,
                  I3 =>  '0' );

  -- Alias \STORE1\   
  \=32208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32208\,
                  I0 =>  \ST1/\,
                  I1 =>  \32206\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STORE1/\  
  \=32209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32209\,
                  I0 =>  \32208\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \STFET1/\  
  \=32210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32210\,
                  I0 =>  \32208\,
                  I1 =>  \32216\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32211\,
                  I0 =>  \MREAD\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32212\,
                  I0 =>  \32203\,
                  I1 =>  \32211\,
                  I2 =>  \32238\,
                  I3 =>  '0' );

  \:32213\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32213\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32213\,
                   R => '0',
                   S => SYSRESET );

  \=32213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32213\,
                  I0 =>  \32212\,
                  I1 =>  \32214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32214\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32214\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32214\,
                   R => SYSRESET,
                   S => '0' );

  \=32214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32214\,
                  I0 =>  \32213\,
                  I1 =>  \GOJAM\,
                  I2 =>  \32218\,
                  I3 =>  '0' );

  -- Alias \MON/\     
  \=32215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32215\,
                  I0 =>  \32207\,
                  I1 =>  \32214\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FETCH1\   
  \=32216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32216\,
                  I0 =>  \ST1/\,
                  I1 =>  \32213\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FETCH0\   
  \=32217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32217\,
                  I0 =>  \ST0/\,
                  I1 =>  \32215\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32218\,
                  I0 =>  \32215\,
                  I1 =>  \32234\,
                  I2 =>  \ST1/\,
                  I3 =>  '0' );

  -- Alias \FETCH0/\  
  \=32219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32219\,
                  I0 =>  \32217\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32220\,
                  I0 =>  \MLDCH\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32221\,
                  I0 =>  \32203\,
                  I1 =>  \32220\,
                  I2 =>  \32238\,
                  I3 =>  '0' );

  \:32222\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32222\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32222\,
                   R => '0',
                   S => SYSRESET );

  \=32222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32222\,
                  I0 =>  \32221\,
                  I1 =>  \32223\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INOTLD\   
  \:32223\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32223\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32223\,
                   R => SYSRESET,
                   S => '0' );

  \=32223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32223\,
                  I0 =>  \32222\,
                  I1 =>  \32233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32224\,
                  I0 =>  \MRDCH\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32225\,
                  I0 =>  \32203\,
                  I1 =>  \32224\,
                  I2 =>  \32238\,
                  I3 =>  '0' );

  \:32226\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32226\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32226\,
                   R => '0',
                   S => SYSRESET );

  \=32226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32226\,
                  I0 =>  \32225\,
                  I1 =>  \32227\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INOTRD\   
  \:32227\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32227\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32227\,
                   R => SYSRESET,
                   S => '0' );

  \=32227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32227\,
                  I0 =>  \32226\,
                  I1 =>  \32233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32228\,
                  I0 =>  \32207\,
                  I1 =>  \32214\,
                  I2 =>  '0',
                  I3 => \&32229\ );

  -- Alias \32228\    
  \=32229\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32229\,
                  I0 =>  \32223\,
                  I1 =>  \32227\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MREQIN\   
  \=32230\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32230\,
                  I0 =>  \32228\,
                  I1 =>  \32228\,
                  I2 =>  \32228\,
                  I3 =>  '0' );

  -- Alias \MON+CH\   
  \=32231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32231\,
                  I0 =>  \32228\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32232\,
                  I0 =>  \32259\,
                  I1 =>  \T11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32233\,
                  I0 =>  \T12/\,
                  I1 =>  \CT\,
                  I2 =>  \PHS2/\,
                  I3 =>  '0' );

  \=32234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32234\,
                  I0 =>  \32233\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32236\    
  \=32235\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32235\,
                  I0 =>  \MRDCH\,
                  I1 =>  \MLDCH\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32236\,
                  I0 =>  \MREAD\,
                  I1 =>  \MLOAD\,
                  I2 =>  '0',
                  I3 => \&32235\ );

  \=32237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32237\,
                  I0 =>  \PHS2/\,
                  I1 =>  \32236\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32238\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32238\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32238\,
                   R => '0',
                   S => SYSRESET );

  \=32238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32238\,
                  I0 =>  \32237\,
                  I1 =>  \32239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32239\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32239\,
                   R => SYSRESET,
                   S => '0' );

  \=32239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32239\,
                  I0 =>  \32238\,
                  I1 =>  \GOJAM\,
                  I2 =>  \32232\,
                  I3 =>  '0' );

  -- Alias \32241\    
  \=32240\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32240\,
                  I0 =>  \32203\,
                  I1 =>  \MNHNC\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32241\,
                  I0 =>  \32239\,
                  I1 =>  \CTROR/\,
                  I2 =>  '0',
                  I3 => \&32240\ );

  \=32242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32242\,
                  I0 =>  \CTROR/\,
                  I1 =>  \32239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32243\,
                  I0 =>  \32242\,
                  I1 =>  \T12/\,
                  I2 =>  \PHS3/\,
                  I3 =>  '0' );

  \:32244\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32244\,
                   R => '0',
                   S => SYSRESET );

  \=32244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32244\,
                  I0 =>  \32241\,
                  I1 =>  \32245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32245\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32245\,
                   R => SYSRESET,
                   S => '0' );

  \=32245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32245\,
                  I0 =>  \32244\,
                  I1 =>  \32243\,
                  I2 =>  \GOJAM\,
                  I3 =>  '0' );

  \=32246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32246\,
                  I0 =>  \T02/\,
                  I1 =>  \32244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INCSET/\  
  \=32247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32247\,
                  I0 =>  \32246\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INKL/\    
  \=32249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32249\,
                  I0 =>  \32245\,
                  I1 =>  \32245\,
                  I2 =>  '0',
                  I3 => \&32250\ );

  -- Alias \32249\    
  \=32250\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32250\,
                  I0 =>  \32231\,
                  I1 =>  \32231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INKL\     
  \=32251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32251\,
                  I0 =>  \32249\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MINKL\    
  \=32253\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32253\,
                  I0 =>  \32249\,
                  I1 =>  \32249\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSSB\     
  \=32254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32254\,
                  I0 =>  \32244\,
                  I1 =>  \T07/\,
                  I2 =>  \PHS3/\,
                  I3 =>  '0' );

  -- Alias \BKTF/\    
  \=32255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32255\,
                  I0 =>  \T10/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHINC/\   
  \=32256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32256\,
                  I0 =>  \INOTLD\,
                  I1 =>  \INOTRD\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \INKBT1\   
  \=32257\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32257\,
                  I0 =>  \STD2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SCAS17\   
  \=32258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32258\,
                  I0 =>  \FS17\,
                  I1 =>  \DOSCAL\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32259\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32259\,
                  I0 =>  \32216\,
                  I1 =>  \32208\,
                  I2 =>  \CHINC\,
                  I3 =>  '0' );

  -- **********************************
  -- ***                            ***
  -- ***  A21/3 - COUNTER CELL II.  ***
  -- ***                            ***
  -- **********************************

  \=32501\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32501\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32502\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32502\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32502\,
                   R => '0',
                   S => SYSRESET );

  \=32502\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32502\,
                  I0 =>  \BMAGXP\,
                  I1 =>  \32503\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32503\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32503\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32503\,
                   R => SYSRESET,
                   S => '0' );

  \=32503\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32503\,
                  I0 =>  \32502\,
                  I1 =>  \32512\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32504\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32504\,
                  I0 =>  \32503\,
                  I1 =>  \32510\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32505\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32505\,
                  I0 =>  \32501\,
                  I1 =>  \32504\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32506\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32506\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32506\,
                   R => '0',
                   S => SYSRESET );

  \=32506\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32506\,
                  I0 =>  \32505\,
                  I1 =>  \32507\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32507\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32507\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32507\,
                   R => SYSRESET,
                   S => '0' );

  \=32507\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32507\,
                  I0 =>  \32506\,
                  I1 =>  \32512\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C42A\     
  \=32508\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32508\,
                  I0 =>  \CG13\,
                  I1 =>  \32506\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32509\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32509\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32509\,
                   R => '0',
                   S => SYSRESET );

  \=32509\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32509\,
                  I0 =>  \BMAGXM\,
                  I1 =>  \32510\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32510\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32510\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32510\,
                   R => SYSRESET,
                   S => '0' );

  \=32510\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32510\,
                  I0 =>  \32509\,
                  I1 =>  \32512\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32511\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32511\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C42R\     
  \=32512\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32512\,
                  I0 =>  \32511\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  -- Alias \C42P\     
  \=32513\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32513\,
                  I0 =>  \32502\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  -- Alias \C42M\     
  \=32514\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32514\,
                  I0 =>  \32509\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB2/\,
                  I3 =>  '0' );

  \:32515\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32515\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32515\,
                   R => '0',
                   S => SYSRESET );

  \=32515\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32515\,
                  I0 =>  \BMAGYP\,
                  I1 =>  \32516\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32516\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32516\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32516\,
                   R => SYSRESET,
                   S => '0' );

  \=32516\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32516\,
                  I0 =>  \32515\,
                  I1 =>  \32526\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32517\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32517\,
                  I0 =>  \32516\,
                  I1 =>  \32525\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32518\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32518\,
                  I0 =>  \32501\,
                  I1 =>  \32517\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32519\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32519\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32519\,
                   R => '0',
                   S => SYSRESET );

  \=32519\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32519\,
                  I0 =>  \32518\,
                  I1 =>  \32520\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32520\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32520\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32520\,
                   R => SYSRESET,
                   S => '0' );

  \=32520\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32520\,
                  I0 =>  \32519\,
                  I1 =>  \32526\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C43A\     
  \=32521\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32521\,
                  I0 =>  \CG13\,
                  I1 =>  \32507\,
                  I2 =>  \32519\,
                  I3 =>  '0' );

  \=32522\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32522\,
                  I0 =>  \CG13\,
                  I1 =>  \32520\,
                  I2 =>  \32507\,
                  I3 =>  '0' );

  -- Alias \CG15\     
  \=32523\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32523\,
                  I0 =>  \32522\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32524\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32524\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32524\,
                   R => '0',
                   S => SYSRESET );

  \=32524\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32524\,
                  I0 =>  \BMAGYM\,
                  I1 =>  \32525\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32525\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32525\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32525\,
                   R => SYSRESET,
                   S => '0' );

  \=32525\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32525\,
                  I0 =>  \32524\,
                  I1 =>  \32526\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C43R\     
  \=32526\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32526\,
                  I0 =>  \32511\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  -- Alias \C43P\     
  \=32527\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32527\,
                  I0 =>  \32515\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  -- Alias \C43M\     
  \=32528\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32528\,
                  I0 =>  \32524\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB3/\,
                  I3 =>  '0' );

  \:32529\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32529\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32529\,
                   R => '0',
                   S => SYSRESET );

  \=32529\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32529\,
                  I0 =>  \EMSD\,
                  I1 =>  \32530\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32530\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32530\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32530\,
                   R => SYSRESET,
                   S => '0' );

  \=32530\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32530\,
                  I0 =>  \32529\,
                  I1 =>  \32535\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32531\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32531\,
                  I0 =>  \32501\,
                  I1 =>  \32529\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32532\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32532\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32532\,
                   R => '0',
                   S => SYSRESET );

  \=32532\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32532\,
                  I0 =>  \32531\,
                  I1 =>  \32533\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32533\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32533\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32533\,
                   R => SYSRESET,
                   S => '0' );

  \=32533\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32533\,
                  I0 =>  \32532\,
                  I1 =>  \32535\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C56A\     
  \=32534\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32534\,
                  I0 =>  \32532\,
                  I1 =>  \CG23\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C56R\     
  \=32535\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32535\,
                  I0 =>  \32511\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  \:32536\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32536\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32536\,
                   R => '0',
                   S => SYSRESET );

  \=32536\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32536\,
                  I0 =>  \OTLNKM\,
                  I1 =>  \32537\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32537\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32537\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32537\,
                   R => SYSRESET,
                   S => '0' );

  \=32537\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32537\,
                  I0 =>  \32536\,
                  I1 =>  \32542\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32538\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32538\,
                  I0 =>  \32501\,
                  I1 =>  \32536\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32539\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32539\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32539\,
                   R => '0',
                   S => SYSRESET );

  \=32539\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32539\,
                  I0 =>  \32538\,
                  I1 =>  \32540\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32540\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32540\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32540\,
                   R => SYSRESET,
                   S => '0' );

  \=32540\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32540\,
                  I0 =>  \32539\,
                  I1 =>  \32542\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C57A\     
  \=32541\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32541\,
                  I0 =>  \CG23\,
                  I1 =>  \32539\,
                  I2 =>  \32533\,
                  I3 =>  '0' );

  -- Alias \C57R\     
  \=32542\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32542\,
                  I0 =>  \32511\,
                  I1 =>  \CA5/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  \:32543\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32543\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32543\,
                   R => '0',
                   S => SYSRESET );

  \=32543\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32543\,
                  I0 =>  \ALTM\,
                  I1 =>  \32544\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32544\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32544\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32544\,
                   R => SYSRESET,
                   S => '0' );

  \=32544\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32544\,
                  I0 =>  \32543\,
                  I1 =>  \32553\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32545\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32545\,
                  I0 =>  \32501\,
                  I1 =>  \32543\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32546\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32546\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32546\,
                   R => '0',
                   S => SYSRESET );

  \=32546\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32546\,
                  I0 =>  \32545\,
                  I1 =>  \32547\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32547\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32547\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32547\,
                   R => SYSRESET,
                   S => '0' );

  \=32547\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32547\,
                  I0 =>  \32546\,
                  I1 =>  \32553\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \32549\    
  \=32548\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32548\,
                  I0 =>  \CG23\,
                  I1 =>  \32533\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C60A\     
  \=32549\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32549\,
                  I0 =>  \32540\,
                  I1 =>  \32546\,
                  I2 =>  '0',
                  I3 => \&32548\ );

  -- Alias \CTROR/\   
  \=32550\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32550\,
                  I0 =>  \CG23\,
                  I1 =>  \32533\,
                  I2 =>  '0',
                  I3 => \&32551\ );

  -- Alias \32550\    
  \=32551\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&32551\,
                  I0 =>  \32540\,
                  I1 =>  \32547\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CTROR\    
  \=32552\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32552\,
                  I0 =>  \32550\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C60R\     
  \=32553\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32553\,
                  I0 =>  \32511\,
                  I1 =>  \CA6/\,
                  I2 =>  \CXB0/\,
                  I3 =>  '0' );

  -- Alias \CA5/\     
  \=32554\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32554\,
                  I0 =>  \OCTAD5\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CXB5/\    
  \=32556\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32556\,
                  I0 =>  \XB5\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHINC\    
  \=32558\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32558\,
                  I0 =>  \CHINC/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32601\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32601\,
                  I0 =>  \BKTF/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32602\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32602\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32602\,
                   R => '0',
                   S => SYSRESET );

  \=32602\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32602\,
                  I0 =>  \BMAGZP\,
                  I1 =>  \32603\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32603\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32603\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32603\,
                   R => SYSRESET,
                   S => '0' );

  \=32603\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32603\,
                  I0 =>  \32602\,
                  I1 =>  \32612\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32604\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32604\,
                  I0 =>  \32603\,
                  I1 =>  \32610\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32605\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32605\,
                  I0 =>  \32601\,
                  I1 =>  \32604\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32606\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32606\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32606\,
                   R => '0',
                   S => SYSRESET );

  \=32606\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32606\,
                  I0 =>  \32605\,
                  I1 =>  \32607\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32607\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32607\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32607\,
                   R => SYSRESET,
                   S => '0' );

  \=32607\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32607\,
                  I0 =>  \32606\,
                  I1 =>  \32612\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C44A\     
  \=32608\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32608\,
                  I0 =>  \CG15\,
                  I1 =>  \32606\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32609\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32609\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32609\,
                   R => '0',
                   S => SYSRESET );

  \=32609\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32609\,
                  I0 =>  \BMAGZM\,
                  I1 =>  \32610\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32610\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32610\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32610\,
                   R => SYSRESET,
                   S => '0' );

  \=32610\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32610\,
                  I0 =>  \32609\,
                  I1 =>  \32612\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32611\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32611\,
                  I0 =>  \RSSB\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C44R\     
  \=32612\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32612\,
                  I0 =>  \32611\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  -- Alias \C44P\     
  \=32613\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32613\,
                  I0 =>  \32602\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  -- Alias \C44M\     
  \=32614\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32614\,
                  I0 =>  \32609\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB4/\,
                  I3 =>  '0' );

  \:32615\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32615\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32615\,
                   R => '0',
                   S => SYSRESET );

  \=32615\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32615\,
                  I0 =>  \INLNKP\,
                  I1 =>  \32616\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32616\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32616\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32616\,
                   R => SYSRESET,
                   S => '0' );

  \=32616\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32616\,
                  I0 =>  \32615\,
                  I1 =>  \32626\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32617\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32617\,
                  I0 =>  \32616\,
                  I1 =>  \32625\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32618\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32618\,
                  I0 =>  \32601\,
                  I1 =>  \32617\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32619\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32619\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32619\,
                   R => '0',
                   S => SYSRESET );

  \=32619\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32619\,
                  I0 =>  \32618\,
                  I1 =>  \32620\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32620\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32620\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32620\,
                   R => SYSRESET,
                   S => '0' );

  \=32620\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32620\,
                  I0 =>  \32619\,
                  I1 =>  \32626\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C45A\     
  \=32621\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32621\,
                  I0 =>  \CG15\,
                  I1 =>  \32607\,
                  I2 =>  \32619\,
                  I3 =>  '0' );

  \=32622\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32622\,
                  I0 =>  \CG15\,
                  I1 =>  \32620\,
                  I2 =>  \32607\,
                  I3 =>  '0' );

  -- Alias \CG16\     
  \=32623\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32623\,
                  I0 =>  \32622\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32624\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32624\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32624\,
                   R => '0',
                   S => SYSRESET );

  \=32624\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32624\,
                  I0 =>  \INLNKM\,
                  I1 =>  \32625\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32625\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32625\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32625\,
                   R => SYSRESET,
                   S => '0' );

  \=32625\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32625\,
                  I0 =>  \32624\,
                  I1 =>  \32626\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C45R\     
  \=32626\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32626\,
                  I0 =>  \32611\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  -- Alias \C45P\     
  \=32627\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32627\,
                  I0 =>  \32615\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  -- Alias \C45M\     
  \=32628\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32628\,
                  I0 =>  \32624\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB5/\,
                  I3 =>  '0' );

  \:32629\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32629\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32629\,
                   R => '0',
                   S => SYSRESET );

  \=32629\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32629\,
                  I0 =>  \RNRADP\,
                  I1 =>  \32630\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32630\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32630\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32630\,
                   R => SYSRESET,
                   S => '0' );

  \=32630\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32630\,
                  I0 =>  \32629\,
                  I1 =>  \32635\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32631\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32631\,
                  I0 =>  \32601\,
                  I1 =>  \32638\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32632\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32632\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32632\,
                   R => '0',
                   S => SYSRESET );

  \=32632\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32632\,
                  I0 =>  \32631\,
                  I1 =>  \32633\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32633\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32633\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32633\,
                   R => SYSRESET,
                   S => '0' );

  \=32633\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32633\,
                  I0 =>  \32632\,
                  I1 =>  \32635\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C46A\     
  \=32634\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32634\,
                  I0 =>  \32632\,
                  I1 =>  \CG16\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C46R\     
  \=32635\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32635\,
                  I0 =>  \32611\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  \:32636\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32636\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32636\,
                   R => '0',
                   S => SYSRESET );

  \=32636\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32636\,
                  I0 =>  \RNRADM\,
                  I1 =>  \32637\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32637\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32637\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32637\,
                   R => SYSRESET,
                   S => '0' );

  \=32637\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32637\,
                  I0 =>  \32636\,
                  I1 =>  \32635\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32638\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32638\,
                  I0 =>  \32630\,
                  I1 =>  \32637\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C46P\     
  \=32639\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32639\,
                  I0 =>  \32629\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB6/\,
                  I3 =>  '0' );

  -- Alias \C46M\     
  \=32640\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32640\,
                  I0 =>  \CXB6/\,
                  I1 =>  \CA4/\,
                  I2 =>  \32636\,
                  I3 =>  '0' );

  \:32643\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32643\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32643\,
                   R => '0',
                   S => SYSRESET );

  \=32643\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32643\,
                  I0 =>  \GYROD\,
                  I1 =>  \32644\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32644\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32644\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32644\,
                   R => SYSRESET,
                   S => '0' );

  \=32644\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32644\,
                  I0 =>  \32643\,
                  I1 =>  \32653\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=32645\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32645\,
                  I0 =>  \32601\,
                  I1 =>  \32643\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32646\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \32646\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32646\,
                   R => '0',
                   S => SYSRESET );

  \=32646\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32646\,
                  I0 =>  \32645\,
                  I1 =>  \32647\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:32647\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \32647\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$32647\,
                   R => SYSRESET,
                   S => '0' );

  \=32647\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$32647\,
                  I0 =>  \32646\,
                  I1 =>  \32653\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C47A\     
  \=32649\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32649\,
                  I0 =>  \CG16\,
                  I1 =>  \32646\,
                  I2 =>  \32633\,
                  I3 =>  '0' );

  \=32650\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32650\,
                  I0 =>  \CG16\,
                  I1 =>  \32647\,
                  I2 =>  \32633\,
                  I3 =>  '0' );

  -- Alias \CG26\     
  \=32652\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32652\,
                  I0 =>  \32650\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \C47R\     
  \=32653\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32653\,
                  I0 =>  \32611\,
                  I1 =>  \CA4/\,
                  I2 =>  \CXB7/\,
                  I3 =>  '0' );

  -- Alias \CXB0/\    
  \=32654\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32654\,
                  I0 =>  \XB0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CXB6/\    
  \=32656\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32656\,
                  I0 =>  \XB6\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RQ/\      
  \=32658\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \32658\,
                  I0 =>  \RQ\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- **************************
  -- ***                    ***
  -- ***  A22/1 - INOUT V.  ***
  -- ***                    ***
  -- **************************

  \=47101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47101\,
                  I0 =>  \DKSTRT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DLKCLR\   
  \=47102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47102\,
                  I0 =>  \47101\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47104\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47104\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47104\,
                   R => '0',
                   S => SYSRESET );

  \=47104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47104\,
                  I0 =>  \47105\,
                  I1 =>  \END\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RDOUT/\   
  \:47105\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47105\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47105\,
                   R => SYSRESET,
                   S => '0' );

  \=47105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47105\,
                  I0 =>  \47102\,
                  I1 =>  \47104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ADVCTR\   
  \=47106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47106\,
                  I0 =>  \47105\,
                  I1 =>  \WDORDR\,
                  I2 =>  \BSYNC/\,
                  I3 =>  '0' );

  \=47107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47107\,
                  I0 =>  \47102\,
                  I1 =>  \47106\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47108\,
                  I0 =>  \47107\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \1CNT\     
  \:47109\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47109\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47109\,
                   R => SYSRESET,
                   S => '0' );

  \=47109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47109\,
                  I0 =>  \47113\,
                  I1 =>  \47110\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47110\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47110\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47110\,
                   R => SYSRESET,
                   S => '0' );

  \=47110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47110\,
                  I0 =>  \47109\,
                  I1 =>  \47108\,
                  I2 =>  \47111\,
                  I3 =>  '0' );

  \:47111\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47111\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47111\,
                   R => SYSRESET,
                   S => '0' );

  \=47111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47111\,
                  I0 =>  \47110\,
                  I1 =>  \47108\,
                  I2 =>  \47112\,
                  I3 =>  '0' );

  \:47112\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47112\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47112\,
                   R => '0',
                   S => SYSRESET );

  \=47112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47112\,
                  I0 =>  \47111\,
                  I1 =>  \47114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47113\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47113\,
                   R => '0',
                   S => SYSRESET );

  \=47113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47113\,
                  I0 =>  \47110\,
                  I1 =>  \47114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47114\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47114\,
                   R => SYSRESET,
                   S => '0' );

  \=47114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47114\,
                  I0 =>  \47113\,
                  I1 =>  \47102\,
                  I2 =>  \47111\,
                  I3 =>  '0' );

  -- Alias \DKCTR1/\  
  \=47115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47115\,
                  I0 =>  \47113\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR1\   
  \=47116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47116\,
                  I0 =>  \47114\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47117\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47117\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47117\,
                   R => SYSRESET,
                   S => '0' );

  \=47117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47117\,
                  I0 =>  \47121\,
                  I1 =>  \47118\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47118\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47118\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47118\,
                   R => SYSRESET,
                   S => '0' );

  \=47118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47118\,
                  I0 =>  \47117\,
                  I1 =>  \47112\,
                  I2 =>  \47119\,
                  I3 =>  '0' );

  \:47119\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47119\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47119\,
                   R => SYSRESET,
                   S => '0' );

  \=47119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47119\,
                  I0 =>  \47118\,
                  I1 =>  \47112\,
                  I2 =>  \47120\,
                  I3 =>  '0' );

  \:47120\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47120\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47120\,
                   R => '0',
                   S => SYSRESET );

  \=47120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47120\,
                  I0 =>  \47119\,
                  I1 =>  \47122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47121\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47121\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47121\,
                   R => '0',
                   S => SYSRESET );

  \=47121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47121\,
                  I0 =>  \47118\,
                  I1 =>  \47122\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47122\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47122\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47122\,
                   R => SYSRESET,
                   S => '0' );

  \=47122\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47122\,
                  I0 =>  \47121\,
                  I1 =>  \47102\,
                  I2 =>  \47119\,
                  I3 =>  '0' );

  -- Alias \DKCTR2/\  
  \=47123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47123\,
                  I0 =>  \47121\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR2\   
  \=47124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47124\,
                  I0 =>  \47122\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47125\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47125\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47125\,
                   R => SYSRESET,
                   S => '0' );

  \=47125\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47125\,
                  I0 =>  \47129\,
                  I1 =>  \47126\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47126\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47126\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47126\,
                   R => SYSRESET,
                   S => '0' );

  \=47126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47126\,
                  I0 =>  \47125\,
                  I1 =>  \47120\,
                  I2 =>  \47127\,
                  I3 =>  '0' );

  \:47127\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47127\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47127\,
                   R => SYSRESET,
                   S => '0' );

  \=47127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47127\,
                  I0 =>  \47126\,
                  I1 =>  \47120\,
                  I2 =>  \47128\,
                  I3 =>  '0' );

  \:47128\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47128\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47128\,
                   R => '0',
                   S => SYSRESET );

  \=47128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47128\,
                  I0 =>  \47127\,
                  I1 =>  \47130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47129\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47129\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47129\,
                   R => '0',
                   S => SYSRESET );

  \=47129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47129\,
                  I0 =>  \47126\,
                  I1 =>  \47130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47130\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47130\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47130\,
                   R => SYSRESET,
                   S => '0' );

  \=47130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47130\,
                  I0 =>  \47129\,
                  I1 =>  \47102\,
                  I2 =>  \47127\,
                  I3 =>  '0' );

  -- Alias \DKCTR3/\  
  \=47131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47131\,
                  I0 =>  \47129\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR3\   
  \=47132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47132\,
                  I0 =>  \47130\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47133\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47133\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47133\,
                   R => SYSRESET,
                   S => '0' );

  \=47133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47133\,
                  I0 =>  \47137\,
                  I1 =>  \47134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47134\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47134\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47134\,
                   R => SYSRESET,
                   S => '0' );

  \=47134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47134\,
                  I0 =>  \47133\,
                  I1 =>  \47128\,
                  I2 =>  \47135\,
                  I3 =>  '0' );

  \:47135\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47135\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47135\,
                   R => SYSRESET,
                   S => '0' );

  \=47135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47135\,
                  I0 =>  \47134\,
                  I1 =>  \47128\,
                  I2 =>  \47136\,
                  I3 =>  '0' );

  \:47136\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47136\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47136\,
                   R => '0',
                   S => SYSRESET );

  \=47136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47136\,
                  I0 =>  \47135\,
                  I1 =>  \47138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR4\   
  \:47137\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47137\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47137\,
                   R => '0',
                   S => SYSRESET );

  \=47137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47137\,
                  I0 =>  \47134\,
                  I1 =>  \47138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR4/\  
  \:47138\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47138\,
                   R => SYSRESET,
                   S => '0' );

  \=47138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47138\,
                  I0 =>  \47137\,
                  I1 =>  \47102\,
                  I2 =>  \47135\,
                  I3 =>  '0' );

  -- Alias \16CNT\    
  \:47139\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47139\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47139\,
                   R => SYSRESET,
                   S => '0' );

  \=47139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47139\,
                  I0 =>  \47143\,
                  I1 =>  \47140\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47140\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47140\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47140\,
                   R => SYSRESET,
                   S => '0' );

  \=47140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47140\,
                  I0 =>  \47139\,
                  I1 =>  \47136\,
                  I2 =>  \47141\,
                  I3 =>  '0' );

  \:47141\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47141\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47141\,
                   R => SYSRESET,
                   S => '0' );

  \=47141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47141\,
                  I0 =>  \47140\,
                  I1 =>  \47136\,
                  I2 =>  \47142\,
                  I3 =>  '0' );

  -- Alias \32CNT\    
  \:47142\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47142\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47142\,
                   R => '0',
                   S => SYSRESET );

  \=47142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47142\,
                  I0 =>  \47141\,
                  I1 =>  \47144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR5\   
  \:47143\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47143\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47143\,
                   R => '0',
                   S => SYSRESET );

  \=47143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47143\,
                  I0 =>  \47140\,
                  I1 =>  \47144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKCTR5/\  
  \:47144\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47144\,
                   R => SYSRESET,
                   S => '0' );

  \=47144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47144\,
                  I0 =>  \47143\,
                  I1 =>  \47102\,
                  I2 =>  \47141\,
                  I3 =>  '0' );

  \=47145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47145\,
                  I0 =>  \BSYNC/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47147\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47147\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47147\,
                   R => SYSRESET,
                   S => '0' );

  \=47147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47147\,
                  I0 =>  \47145\,
                  I1 =>  \47150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47148\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47148\,
                   R => SYSRESET,
                   S => '0' );

  \=47148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47148\,
                  I0 =>  \47147\,
                  I1 =>  \47151\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47149\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47149\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47149\,
                   R => SYSRESET,
                   S => '0' );

  \=47149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47149\,
                  I0 =>  \47151\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47150\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47150\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47150\,
                   R => '0',
                   S => SYSRESET );

  \=47150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47150\,
                  I0 =>  \47149\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47151\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47151\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47151\,
                   R => '0',
                   S => SYSRESET );

  \=47151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47151\,
                  I0 =>  \47145\,
                  I1 =>  \47148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47153\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47153\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47153\,
                   R => SYSRESET,
                   S => '0' );

  \=47153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47153\,
                  I0 =>  \DLKCLR\,
                  I1 =>  \47154\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WDORDR\   
  \:47154\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47154\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47154\,
                   R => '0',
                   S => SYSRESET );

  \=47154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47154\,
                  I0 =>  \47153\,
                  I1 =>  \47147\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47155\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47156\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47156\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47156\,
                   R => '0',
                   S => SYSRESET );

  \=47156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47156\,
                  I0 =>  \47157\,
                  I1 =>  \47155\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47157\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47157\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47157\,
                   R => SYSRESET,
                   S => '0' );

  \=47157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47157\,
                  I0 =>  \CCH13\,
                  I1 =>  \47156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1307\   
  \=47158\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47158\,
                  I0 =>  \RCH13/\,
                  I1 =>  \47156\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ORDRBT\   
  \=47159\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47159\,
                  I0 =>  \47156\,
                  I1 =>  \47153\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F12B/\    
  \=47161\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47161\,
                  I0 =>  \F12B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F14H\     
  \=47162\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47162\,
                  I0 =>  \F12B/\,
                  I1 =>  \FS14\,
                  I2 =>  \FS13/\,
                  I3 =>  '0' );

  \=47201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47201\,
                  I0 =>  \XB3/\,
                  I1 =>  \XT1/\,
                  I2 =>  \WCHG/\,
                  I3 =>  '0' );

  -- Alias \WCH13/\   
  \=47202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47202\,
                  I0 =>  \47201\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47205\,
                  I0 =>  \XT1/\,
                  I1 =>  \XB3/\,
                  I2 =>  \CCHG/\,
                  I3 =>  '0' );

  \=47206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47206\,
                  I0 =>  \47205\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH13\    
  \=47207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47207\,
                  I0 =>  \47206\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47210\,
                  I0 =>  \XB3/\,
                  I1 =>  \XT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH13/\   
  \=47211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47211\,
                  I0 =>  \47210\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47214\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XB4/\,
                  I2 =>  \XT1/\,
                  I3 =>  '0' );

  -- Alias \WCH14/\   
  \=47215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47215\,
                  I0 =>  \47214\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47218\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XT1/\,
                  I2 =>  \XB4/\,
                  I3 =>  '0' );

  \=47219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47219\,
                  I0 =>  \GOJAM\,
                  I1 =>  \47218\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH14\    
  \=47220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47220\,
                  I0 =>  \47219\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47223\,
                  I0 =>  \XB4/\,
                  I1 =>  \XT1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH14/\   
  \=47224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47224\,
                  I0 =>  \47223\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BSYNC/\   
  \=47227\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47227\,
                  I0 =>  \DKBSNC\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47228\,
                  I0 =>  \DKCTR1\,
                  I1 =>  \DKCTR3\,
                  I2 =>  \DKCTR2\,
                  I3 =>  '0' );

  -- Alias \LOW0/\    
  \=47229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47229\,
                  I0 =>  \47228\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47230\,
                  I0 =>  \DKCTR1/\,
                  I1 =>  \DKCTR3\,
                  I2 =>  \DKCTR2\,
                  I3 =>  '0' );

  -- Alias \LOW1/\    
  \=47231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47231\,
                  I0 =>  \47230\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47232\,
                  I0 =>  \DKCTR1\,
                  I1 =>  \DKCTR3\,
                  I2 =>  \DKCTR2/\,
                  I3 =>  '0' );

  -- Alias \LOW2/\    
  \=47233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47233\,
                  I0 =>  \47232\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47234\,
                  I0 =>  \DKCTR1/\,
                  I1 =>  \DKCTR3\,
                  I2 =>  \DKCTR2/\,
                  I3 =>  '0' );

  -- Alias \LOW3/\    
  \=47235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47235\,
                  I0 =>  \47234\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47236\,
                  I0 =>  \DKCTR2\,
                  I1 =>  \DKCTR3/\,
                  I2 =>  \DKCTR1\,
                  I3 =>  '0' );

  -- Alias \LOW4/\    
  \=47237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47237\,
                  I0 =>  \47236\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47238\,
                  I0 =>  \DKCTR2\,
                  I1 =>  \DKCTR3/\,
                  I2 =>  \DKCTR1/\,
                  I3 =>  '0' );

  -- Alias \LOW5/\    
  \=47239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47239\,
                  I0 =>  \47238\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47240\,
                  I0 =>  \DKCTR2/\,
                  I1 =>  \DKCTR3/\,
                  I2 =>  \DKCTR1\,
                  I3 =>  '0' );

  -- Alias \LOW6/\    
  \=47241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47241\,
                  I0 =>  \47240\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47242\,
                  I0 =>  \DKCTR2/\,
                  I1 =>  \DKCTR3/\,
                  I2 =>  \DKCTR1/\,
                  I3 =>  '0' );

  -- Alias \LOW7/\    
  \=47243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47243\,
                  I0 =>  \47242\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47244\,
                  I0 =>  \CHWL16/\,
                  I1 =>  \WCH34/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47245\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47246\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47246\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47246\,
                   R => '0',
                   S => SYSRESET );

  \=47246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47246\,
                  I0 =>  \47244\,
                  I1 =>  \47247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47247\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47247\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47247\,
                   R => SYSRESET,
                   S => '0' );

  \=47247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47247\,
                  I0 =>  \47246\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47248\,
                   R => '0',
                   S => SYSRESET );

  \=47248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47248\,
                  I0 =>  \47245\,
                  I1 =>  \47249\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47249\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47249\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47249\,
                   R => SYSRESET,
                   S => '0' );

  \=47249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47249\,
                  I0 =>  \47248\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47250\,
                  I0 =>  \47229\,
                  I1 =>  \47246\,
                  I2 =>  \HIGH0/\,
                  I3 =>  '0' );

  \=47251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47251\,
                  I0 =>  \47231\,
                  I1 =>  \47248\,
                  I2 =>  \HIGH0/\,
                  I3 =>  '0' );

  -- Alias \47253\    
  \=47252\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47252\,
                  I0 =>  \WRD1B1\,
                  I1 =>  \WRD1BP\,
                  I2 =>  \WRD2B3\,
                  I3 => \&47321\ );

  -- Alias \DATA/\    
  \=47253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47253\,
                  I0 =>  \47250\,
                  I1 =>  \WRD2B2\,
                  I2 =>  \47251\,
                  I3 => \&47252\ );

  \=47254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47254\,
                  I0 =>  \47253\,
                  I1 =>  \WDORDR\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKDAT/\   
  \=47255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47255\,
                  I0 =>  \47254\,
                  I1 =>  \ORDRBT\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DKDATA\   
  \=47256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47256\,
                  I0 =>  \47227\,
                  I1 =>  \RDOUT/\,
                  I2 =>  \DKDAT/\,
                  I3 =>  '0' );

  -- Alias \DKDATB\   
  \=47261\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47261\,
                  I0 =>  \47227\,
                  I1 =>  \RDOUT/\,
                  I2 =>  \DKDAT/\,
                  I3 =>  '0' );

  -- Alias \FS13/\    
  \=47262\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47262\,
                  I0 =>  \FS13\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- **************************
  -- ***                    ***
  -- ***  A22/2 - INOUT V.  ***
  -- ***                    ***
  -- **************************

  \=47301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47301\,
                  I0 =>  \WCH34/\,
                  I1 =>  \PC15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47302\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47302\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47302\,
                   R => '0',
                   S => SYSRESET );

  \=47302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47302\,
                  I0 =>  \47301\,
                  I1 =>  \47303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47303\,
                   R => SYSRESET,
                   S => '0' );

  \=47303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47303\,
                  I0 =>  \47302\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WRD1BP\   
  \=47304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47304\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47302\,
                  I2 =>  \LOW7/\,
                  I3 =>  '0' );

  \=47305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47305\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47306\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47306\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47306\,
                   R => '0',
                   S => SYSRESET );

  \=47306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47306\,
                  I0 =>  \47305\,
                  I1 =>  \47307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47307\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47307\,
                   R => SYSRESET,
                   S => '0' );

  \=47307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47307\,
                  I0 =>  \47306\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WRD1B1\   
  \=47308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47308\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47306\,
                  I2 =>  \LOW6/\,
                  I3 =>  '0' );

  \=47309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47309\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47310\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47310\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47310\,
                   R => '0',
                   S => SYSRESET );

  \=47310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47310\,
                  I0 =>  \47309\,
                  I1 =>  \47311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47311\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47311\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47311\,
                   R => SYSRESET,
                   S => '0' );

  \=47311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47311\,
                  I0 =>  \47310\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47312\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47310\,
                  I2 =>  \LOW5/\,
                  I3 =>  '0' );

  \=47313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47313\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47314\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47314\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47314\,
                   R => '0',
                   S => SYSRESET );

  \=47314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47314\,
                  I0 =>  \47313\,
                  I1 =>  \47315\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47315\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47315\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47315\,
                   R => SYSRESET,
                   S => '0' );

  \=47315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47315\,
                  I0 =>  \47314\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47316\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47314\,
                  I2 =>  \LOW2/\,
                  I3 =>  '0' );

  \=47317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47317\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47318\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47318\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47318\,
                   R => '0',
                   S => SYSRESET );

  \=47318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47318\,
                  I0 =>  \47317\,
                  I1 =>  \47319\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47319\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47319\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47319\,
                   R => SYSRESET,
                   S => '0' );

  \=47319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47319\,
                  I0 =>  \47318\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47320\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47318\,
                  I2 =>  \LOW3/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47321\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47321\,
                  I0 =>  \47312\,
                  I1 =>  \47316\,
                  I2 =>  \47320\,
                  I3 => \&47334\ );

  \=47322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47322\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47323\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47323\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47323\,
                   R => '0',
                   S => SYSRESET );

  \=47323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47323\,
                  I0 =>  \47322\,
                  I1 =>  \47324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47324\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47324\,
                   R => SYSRESET,
                   S => '0' );

  \=47324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47324\,
                  I0 =>  \47323\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47325\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47323\,
                  I2 =>  \LOW4/\,
                  I3 =>  '0' );

  \=47326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47326\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47327\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47327\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47327\,
                   R => '0',
                   S => SYSRESET );

  \=47327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47327\,
                  I0 =>  \47326\,
                  I1 =>  \47328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47328\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47328\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47328\,
                   R => SYSRESET,
                   S => '0' );

  \=47328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47328\,
                  I0 =>  \47327\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47329\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47327\,
                  I2 =>  \LOW5/\,
                  I3 =>  '0' );

  \=47330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47330\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47331\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47331\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47331\,
                   R => '0',
                   S => SYSRESET );

  \=47331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47331\,
                  I0 =>  \47330\,
                  I1 =>  \47332\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47332\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47332\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47332\,
                   R => SYSRESET,
                   S => '0' );

  \=47332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47332\,
                  I0 =>  \47331\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47333\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47331\,
                  I2 =>  \LOW6/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47334\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47334\,
                  I0 =>  \47325\,
                  I1 =>  \47329\,
                  I2 =>  \47333\,
                  I3 => \&47343\ );

  \=47335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47335\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47336\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47336\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47336\,
                   R => '0',
                   S => SYSRESET );

  \=47336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47336\,
                  I0 =>  \47335\,
                  I1 =>  \47337\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47337\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47337\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47337\,
                   R => SYSRESET,
                   S => '0' );

  \=47337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47337\,
                  I0 =>  \47336\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47338\,
                  I0 =>  \HIGH0/\,
                  I1 =>  \47336\,
                  I2 =>  \LOW7/\,
                  I3 =>  '0' );

  \=47339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47339\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47340\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47340\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47340\,
                   R => '0',
                   S => SYSRESET );

  \=47340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47340\,
                  I0 =>  \47339\,
                  I1 =>  \47341\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47341\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47341\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47341\,
                   R => SYSRESET,
                   S => '0' );

  \=47341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47341\,
                  I0 =>  \47340\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47342\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47340\,
                  I2 =>  \LOW0/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47343\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47343\,
                  I0 =>  \47338\,
                  I1 =>  \47342\,
                  I2 =>  \47347\,
                  I3 => \&47360\ );

  \=47344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47344\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47345\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47345\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47345\,
                   R => '0',
                   S => SYSRESET );

  \=47345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47345\,
                  I0 =>  \47344\,
                  I1 =>  \47346\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47346\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47346\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47346\,
                   R => SYSRESET,
                   S => '0' );

  \=47346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47346\,
                  I0 =>  \47345\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47347\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47345\,
                  I2 =>  \LOW1/\,
                  I3 =>  '0' );

  \=47348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47348\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47349\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47349\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47349\,
                   R => '0',
                   S => SYSRESET );

  \=47349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47349\,
                  I0 =>  \47348\,
                  I1 =>  \47350\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47350\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47350\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47350\,
                   R => SYSRESET,
                   S => '0' );

  \=47350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47350\,
                  I0 =>  \47349\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47351\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47349\,
                  I2 =>  \LOW2/\,
                  I3 =>  '0' );

  \=47352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47352\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47353\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47353\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47353\,
                   R => '0',
                   S => SYSRESET );

  \=47353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47353\,
                  I0 =>  \47352\,
                  I1 =>  \47354\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47354\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47354\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47354\,
                   R => SYSRESET,
                   S => '0' );

  \=47354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47354\,
                  I0 =>  \47353\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47355\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47353\,
                  I2 =>  \LOW3/\,
                  I3 =>  '0' );

  \=47356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47356\,
                  I0 =>  \WCH34/\,
                  I1 =>  \CHWL03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47357\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47357\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47357\,
                   R => '0',
                   S => SYSRESET );

  \=47357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47357\,
                  I0 =>  \47356\,
                  I1 =>  \47358\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47358\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47358\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47358\,
                   R => SYSRESET,
                   S => '0' );

  \=47358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47358\,
                  I0 =>  \47357\,
                  I1 =>  \CCH34\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47359\,
                  I0 =>  \HIGH1/\,
                  I1 =>  \47357\,
                  I2 =>  \LOW4/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47360\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47360\,
                  I0 =>  \47351\,
                  I1 =>  \47355\,
                  I2 =>  \47359\,
                  I3 => \&47421\ );

  \=47401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47401\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47402\,
                   R => '0',
                   S => SYSRESET );

  \=47402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47402\,
                  I0 =>  \47401\,
                  I1 =>  \47403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47403\,
                   R => SYSRESET,
                   S => '0' );

  \=47403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47403\,
                  I0 =>  \47402\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WRD2B2\   
  \=47404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47404\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47402\,
                  I2 =>  \LOW5/\,
                  I3 =>  '0' );

  \=47405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47405\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47406\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47406\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47406\,
                   R => '0',
                   S => SYSRESET );

  \=47406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47406\,
                  I0 =>  \47405\,
                  I1 =>  \47407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47407\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47407\,
                   R => SYSRESET,
                   S => '0' );

  \=47407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47407\,
                  I0 =>  \47406\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WRD2B3\   
  \=47408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47408\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47406\,
                  I2 =>  \LOW4/\,
                  I3 =>  '0' );

  \=47409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47409\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47410\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47410\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47410\,
                   R => '0',
                   S => SYSRESET );

  \=47410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47410\,
                  I0 =>  \47409\,
                  I1 =>  \47411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47411\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47411\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47411\,
                   R => SYSRESET,
                   S => '0' );

  \=47411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47411\,
                  I0 =>  \47410\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47412\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47410\,
                  I2 =>  \LOW3/\,
                  I3 =>  '0' );

  \=47413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47413\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47414\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47414\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47414\,
                   R => '0',
                   S => SYSRESET );

  \=47414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47414\,
                  I0 =>  \47413\,
                  I1 =>  \47415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47415\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47415\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47415\,
                   R => SYSRESET,
                   S => '0' );

  \=47415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47415\,
                  I0 =>  \47414\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47416\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47414\,
                  I2 =>  \LOW0/\,
                  I3 =>  '0' );

  \=47417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47417\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47418\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47418\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47418\,
                   R => '0',
                   S => SYSRESET );

  \=47418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47418\,
                  I0 =>  \47417\,
                  I1 =>  \47419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47419\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47419\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47419\,
                   R => SYSRESET,
                   S => '0' );

  \=47419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47419\,
                  I0 =>  \47418\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47420\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47418\,
                  I2 =>  \LOW1/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47421\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47421\,
                  I0 =>  \47416\,
                  I1 =>  \47420\,
                  I2 =>  \47425\,
                  I3 => \&47434\ );

  \=47422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47422\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47423\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47423\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47423\,
                   R => '0',
                   S => SYSRESET );

  \=47423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47423\,
                  I0 =>  \47422\,
                  I1 =>  \47424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47424\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47424\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47424\,
                   R => SYSRESET,
                   S => '0' );

  \=47424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47424\,
                  I0 =>  \47423\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47425\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47423\,
                  I2 =>  \LOW2/\,
                  I3 =>  '0' );

  \=47426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47426\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47427\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47427\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47427\,
                   R => '0',
                   S => SYSRESET );

  \=47427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47427\,
                  I0 =>  \47426\,
                  I1 =>  \47428\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47428\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47428\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47428\,
                   R => SYSRESET,
                   S => '0' );

  \=47428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47428\,
                  I0 =>  \47427\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47429\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47427\,
                  I2 =>  \LOW3/\,
                  I3 =>  '0' );

  \=47430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47430\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47431\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47431\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47431\,
                   R => '0',
                   S => SYSRESET );

  \=47431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47431\,
                  I0 =>  \47430\,
                  I1 =>  \47432\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47432\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47432\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47432\,
                   R => SYSRESET,
                   S => '0' );

  \=47432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47432\,
                  I0 =>  \47431\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47433\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47431\,
                  I2 =>  \LOW4/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47434\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47434\,
                  I0 =>  \47429\,
                  I1 =>  \47433\,
                  I2 =>  \47438\,
                  I3 => \&47447\ );

  \=47435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47435\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47436\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47436\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47436\,
                   R => '0',
                   S => SYSRESET );

  \=47436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47436\,
                  I0 =>  \47435\,
                  I1 =>  \47437\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47437\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47437\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47437\,
                   R => SYSRESET,
                   S => '0' );

  \=47437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47437\,
                  I0 =>  \47436\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47438\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47438\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47436\,
                  I2 =>  \LOW5/\,
                  I3 =>  '0' );

  \=47439\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47439\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL09/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47440\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47440\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47440\,
                   R => '0',
                   S => SYSRESET );

  \=47440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47440\,
                  I0 =>  \47439\,
                  I1 =>  \47441\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47441\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47441\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47441\,
                   R => SYSRESET,
                   S => '0' );

  \=47441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47441\,
                  I0 =>  \47440\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47442\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47440\,
                  I2 =>  \LOW6/\,
                  I3 =>  '0' );

  \=47443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47443\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47444\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47444\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47444\,
                   R => '0',
                   S => SYSRESET );

  \=47444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47444\,
                  I0 =>  \47443\,
                  I1 =>  \47445\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47445\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47445\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47445\,
                   R => SYSRESET,
                   S => '0' );

  \=47445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47445\,
                  I0 =>  \47444\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47446\,
                  I0 =>  \HIGH2/\,
                  I1 =>  \47444\,
                  I2 =>  \LOW7/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47447\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47447\,
                  I0 =>  \47442\,
                  I1 =>  \47446\,
                  I2 =>  \47451\,
                  I3 => \&47460\ );

  \=47448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47448\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47449\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47449\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47449\,
                   R => '0',
                   S => SYSRESET );

  \=47449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47449\,
                  I0 =>  \47448\,
                  I1 =>  \47450\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47450\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47450\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47450\,
                   R => SYSRESET,
                   S => '0' );

  \=47450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47450\,
                  I0 =>  \47449\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47451\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47449\,
                  I2 =>  \LOW0/\,
                  I3 =>  '0' );

  \=47452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47452\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47453\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47453\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47453\,
                   R => '0',
                   S => SYSRESET );

  \=47453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47453\,
                  I0 =>  \47452\,
                  I1 =>  \47454\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47454\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47454\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47454\,
                   R => SYSRESET,
                   S => '0' );

  \=47454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47454\,
                  I0 =>  \47453\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47455\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47455\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47453\,
                  I2 =>  \LOW1/\,
                  I3 =>  '0' );

  \=47456\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47456\,
                  I0 =>  \WCH35/\,
                  I1 =>  \CHWL05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47457\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \47457\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47457\,
                   R => '0',
                   S => SYSRESET );

  \=47457\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47457\,
                  I0 =>  \47456\,
                  I1 =>  \47458\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:47458\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \47458\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$47458\,
                   R => SYSRESET,
                   S => '0' );

  \=47458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$47458\,
                  I0 =>  \47457\,
                  I1 =>  \CCH35\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=47459\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \47459\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \47457\,
                  I2 =>  \LOW2/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=47460\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&47460\,
                  I0 =>  \47455\,
                  I1 =>  \47459\,
                  I2 =>  \47412\,
                  I3 => \&48117\ );

  -- ***************************
  -- ***                     ***
  -- ***  A23/1 - INOUT VI.  ***
  -- ***                     ***
  -- ***************************

  -- Alias \48102\    
  \=48101\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48101\,
                  I0 =>  \NOXP\,
                  I1 =>  \NOXM\,
                  I2 =>  \NOYP\,
                  I3 =>  '0' );

  \=48102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48102\,
                  I0 =>  \NOYM\,
                  I1 =>  \NOZP\,
                  I2 =>  \NOZM\,
                  I3 => \&48101\ );

  \=48103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48103\,
                  I0 =>  \F18B/\,
                  I1 =>  \48102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48104\,
                  I0 =>  \MISSX\,
                  I1 =>  \MISSY\,
                  I2 =>  \MISSZ\,
                  I3 =>  '0' );

  \=48105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48105\,
                  I0 =>  \F5ASB0/\,
                  I1 =>  \48104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \48107\    
  \=48106\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48106\,
                  I0 =>  \BOTHZ\,
                  I1 =>  \BOTHY\,
                  I2 =>  \BOTHX\,
                  I3 =>  '0' );

  \:48107\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48107\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48107\,
                   R => '0',
                   S => SYSRESET );

  \=48107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48107\,
                  I0 =>  \48103\,
                  I1 =>  \48105\,
                  I2 =>  \48108\,
                  I3 => \&48106\ );

  -- Alias \PIPAFL\   
  \:48108\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48108\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48108\,
                   R => SYSRESET,
                   S => '0' );

  \=48108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48108\,
                  I0 =>  \48107\,
                  I1 =>  \CCH33\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48109\,
                  I0 =>  \CHWL01/\,
                  I1 =>  \48120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48110\,
                  I0 =>  \PC15/\,
                  I1 =>  \48120\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48111\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48111\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48111\,
                   R => '0',
                   S => SYSRESET );

  \=48111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48111\,
                  I0 =>  \48109\,
                  I1 =>  \48112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48112\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48112\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48112\,
                   R => SYSRESET,
                   S => '0' );

  \=48112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48112\,
                  I0 =>  \48111\,
                  I1 =>  \48124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48113\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48113\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48113\,
                   R => '0',
                   S => SYSRESET );

  \=48113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48113\,
                  I0 =>  \48110\,
                  I1 =>  \48114\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48114\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48114\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48114\,
                   R => SYSRESET,
                   S => '0' );

  \=48114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48114\,
                  I0 =>  \48113\,
                  I1 =>  \48124\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48115\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \48111\,
                  I2 =>  \LOW6/\,
                  I3 =>  '0' );

  \=48116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48116\,
                  I0 =>  \HIGH3/\,
                  I1 =>  \48113\,
                  I2 =>  \LOW7/\,
                  I3 =>  '0' );

  -- Alias \DATA/\    
  \=48117\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48117\,
                  I0 =>  \48115\,
                  I1 =>  \48116\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48118\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48118\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XB5/\,
                  I2 =>  \XT3/\,
                  I3 =>  '0' );

  \=48119\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48119\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB5/\,
                  I2 =>  \CCHG/\,
                  I3 =>  '0' );

  -- Alias \WCH35/\   
  \=48120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48120\,
                  I0 =>  \48118\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48123\,
                  I0 =>  \48119\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH35\    
  \=48124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48124\,
                  I0 =>  \48123\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BOTHX\    
  \=48127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48127\,
                  I0 =>  \48129\,
                  I1 =>  \48130\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48128\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48128\,
                  I0 =>  \F5ASB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48129\,
                  I0 =>  \PIPGX+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48130\,
                  I0 =>  \PIPGX-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48131\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48131\,
                  I0 =>  \48130\,
                  I1 =>  \48148\,
                  I2 =>  \48138\,
                  I3 =>  '0' );

  \=48132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48132\,
                  I0 =>  \48137\,
                  I1 =>  \48148\,
                  I2 =>  \48129\,
                  I3 =>  '0' );

  \:48133\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48133\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48133\,
                   R => '0',
                   S => SYSRESET );

  \=48133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48133\,
                  I0 =>  \48131\,
                  I1 =>  \48134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48134\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48134\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48134\,
                   R => SYSRESET,
                   S => '0' );

  \=48134\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48134\,
                  I0 =>  \48133\,
                  I1 =>  \48132\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48135\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48135\,
                  I0 =>  \48128\,
                  I1 =>  \48133\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48136\,
                  I0 =>  \48128\,
                  I1 =>  \48134\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48137\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48137\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48137\,
                   R => '0',
                   S => SYSRESET );

  \=48137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48137\,
                  I0 =>  \48135\,
                  I1 =>  \48138\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48138\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48138\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48138\,
                   R => SYSRESET,
                   S => '0' );

  \=48138\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48138\,
                  I0 =>  \48137\,
                  I1 =>  \48136\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48139\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48139\,
                  I0 =>  \48138\,
                  I1 =>  \48148\,
                  I2 =>  \48129\,
                  I3 =>  '0' );

  \=48140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48140\,
                  I0 =>  \48137\,
                  I1 =>  \48148\,
                  I2 =>  \48130\,
                  I3 =>  '0' );

  \=48141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48141\,
                  I0 =>  \48138\,
                  I1 =>  \48147\,
                  I2 =>  \48130\,
                  I3 =>  '0' );

  \=48142\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48142\,
                  I0 =>  \48137\,
                  I1 =>  \48147\,
                  I2 =>  \48129\,
                  I3 =>  '0' );

  \:48143\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48143\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48143\,
                   R => '0',
                   S => SYSRESET );

  \=48143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48143\,
                  I0 =>  \48139\,
                  I1 =>  \48140\,
                  I2 =>  \48144\,
                  I3 =>  '0' );

  \:48144\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48144\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48144\,
                   R => SYSRESET,
                   S => '0' );

  \=48144\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48144\,
                  I0 =>  \48143\,
                  I1 =>  \48141\,
                  I2 =>  \48142\,
                  I3 =>  '0' );

  \=48145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48145\,
                  I0 =>  \48128\,
                  I1 =>  \48143\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48146\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48146\,
                  I0 =>  \48128\,
                  I1 =>  \48144\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48147\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48147\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48147\,
                   R => '0',
                   S => SYSRESET );

  \=48147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48147\,
                  I0 =>  \48145\,
                  I1 =>  \48148\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48148\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48148\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48148\,
                   R => SYSRESET,
                   S => '0' );

  \=48148\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48148\,
                  I0 =>  \48147\,
                  I1 =>  \48146\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOXM\     
  \:48149\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48149\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48149\,
                   R => '0',
                   S => SYSRESET );

  \=48149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48149\,
                  I0 =>  \PIPGX-\,
                  I1 =>  \48150\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48150\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48150\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48150\,
                   R => SYSRESET,
                   S => '0' );

  \=48150\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48150\,
                  I0 =>  \48149\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOXP\     
  \:48151\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48151\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48151\,
                   R => '0',
                   S => SYSRESET );

  \=48151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48151\,
                  I0 =>  \PIPGX+\,
                  I1 =>  \48152\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48152\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48152\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48152\,
                   R => SYSRESET,
                   S => '0' );

  \=48152\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48152\,
                  I0 =>  \48151\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MISSX\    
  \:48153\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48153\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48153\,
                   R => '0',
                   S => SYSRESET );

  \=48153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48153\,
                  I0 =>  \PIPGX+\,
                  I1 =>  \PIPGX-\,
                  I2 =>  \48154\,
                  I3 =>  '0' );

  \:48154\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48154\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48154\,
                   R => SYSRESET,
                   S => '0' );

  \=48154\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48154\,
                  I0 =>  \48153\,
                  I1 =>  \F5ASB2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPXP\    
  \=48155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48155\,
                  I0 =>  \48138\,
                  I1 =>  \48129\,
                  I2 =>  \48147\,
                  I3 =>  '0' );

  -- Alias \PIPXM\    
  \=48156\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48156\,
                  I0 =>  \48137\,
                  I1 =>  \48130\,
                  I2 =>  \48147\,
                  I3 =>  '0' );

  -- Alias \F18B/\    
  \=48157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48157\,
                  I0 =>  \F18B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR01/\  
  \=48201\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48201\,
                  I0 =>  \CHAT01\,
                  I1 =>  \CHBT01\,
                  I2 =>  \CH1601\,
                  I3 =>  '0' );

  -- Alias \CH01\     
  \=48202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48202\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR01/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR02/\  
  \=48203\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48203\,
                  I0 =>  \CHAT02\,
                  I1 =>  \CHBT02\,
                  I2 =>  \CH1602\,
                  I3 =>  '0' );

  -- Alias \CH02\     
  \=48204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48204\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR02/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR03/\  
  \=48205\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48205\,
                  I0 =>  \CHAT03\,
                  I1 =>  \CHBT03\,
                  I2 =>  \CH1603\,
                  I3 =>  '0' );

  -- Alias \CH03\     
  \=48206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48206\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR03/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR04/\  
  \=48207\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48207\,
                  I0 =>  \CHAT04\,
                  I1 =>  \CHBT04\,
                  I2 =>  \CH1604\,
                  I3 =>  '0' );

  -- Alias \CH04\     
  \=48208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48208\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR04/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR05/\  
  \=48209\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48209\,
                  I0 =>  \CHAT05\,
                  I1 =>  \CHBT05\,
                  I2 =>  '0',
                  I3 => \&48210\ );

  -- Alias \CHOR05/\  
  \=48210\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48210\,
                  I0 =>  \CH1605\,
                  I1 =>  \CH1505\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH05\     
  \=48211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48211\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR06/\  
  \=48212\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48212\,
                  I0 =>  \CHAT06\,
                  I1 =>  \CHBT06\,
                  I2 =>  \CH1606\,
                  I3 =>  '0' );

  -- Alias \CH06\     
  \=48213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48213\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR06/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR07/\  
  \=48214\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48214\,
                  I0 =>  \CHAT07\,
                  I1 =>  \CHBT07\,
                  I2 =>  \CH1607\,
                  I3 =>  '0' );

  -- Alias \CH07\     
  \=48215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48215\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR07/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR08/\  
  \=48216\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48216\,
                  I0 =>  \CHAT08\,
                  I1 =>  \CHBT08\,
                  I2 =>  '0',
                  I3 => \&48217\ );

  -- Alias \CHOR08/\  
  \=48217\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48217\,
                  I0 =>  \CH1108\,
                  I1 =>  \CH1208\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH08\     
  \=48218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48218\,
                  I0 =>  \RCHG/\,
                  I1 =>  \CHOR08/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48219\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XB4/\,
                  I2 =>  \XT3/\,
                  I3 =>  '0' );

  \=48220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48220\,
                  I0 =>  \XT3/\,
                  I1 =>  \XB4/\,
                  I2 =>  \CCHG/\,
                  I3 =>  '0' );

  -- Alias \WCH34/\   
  \=48221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48221\,
                  I0 =>  \48219\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48224\,
                  I0 =>  \48220\,
                  I1 =>  \GOJAM\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH34\    
  \=48225\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48225\,
                  I0 =>  \48224\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BOTHY\    
  \=48228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48228\,
                  I0 =>  \48230\,
                  I1 =>  \48231\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48229\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48229\,
                  I0 =>  \F5ASB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48230\,
                  I0 =>  \PIPGY+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48231\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48231\,
                  I0 =>  \PIPGY-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48232\,
                  I0 =>  \48231\,
                  I1 =>  \48249\,
                  I2 =>  \48239\,
                  I3 =>  '0' );

  \=48233\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48233\,
                  I0 =>  \48238\,
                  I1 =>  \48249\,
                  I2 =>  \48230\,
                  I3 =>  '0' );

  \:48234\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48234\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48234\,
                   R => '0',
                   S => SYSRESET );

  \=48234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48234\,
                  I0 =>  \48232\,
                  I1 =>  \48235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48235\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48235\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48235\,
                   R => SYSRESET,
                   S => '0' );

  \=48235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48235\,
                  I0 =>  \48234\,
                  I1 =>  \48233\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48236\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48236\,
                  I0 =>  \48229\,
                  I1 =>  \48234\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48237\,
                  I0 =>  \48229\,
                  I1 =>  \48235\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48238\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48238\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48238\,
                   R => '0',
                   S => SYSRESET );

  \=48238\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48238\,
                  I0 =>  \48236\,
                  I1 =>  \48239\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48239\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48239\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48239\,
                   R => SYSRESET,
                   S => '0' );

  \=48239\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48239\,
                  I0 =>  \48238\,
                  I1 =>  \48237\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48240\,
                  I0 =>  \48239\,
                  I1 =>  \48249\,
                  I2 =>  \48230\,
                  I3 =>  '0' );

  \=48241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48241\,
                  I0 =>  \48238\,
                  I1 =>  \48249\,
                  I2 =>  \48231\,
                  I3 =>  '0' );

  \=48242\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48242\,
                  I0 =>  \48239\,
                  I1 =>  \48248\,
                  I2 =>  \48231\,
                  I3 =>  '0' );

  \=48243\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48243\,
                  I0 =>  \48238\,
                  I1 =>  \48248\,
                  I2 =>  \48230\,
                  I3 =>  '0' );

  \:48244\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48244\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48244\,
                   R => '0',
                   S => SYSRESET );

  \=48244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48244\,
                  I0 =>  \48240\,
                  I1 =>  \48241\,
                  I2 =>  \48245\,
                  I3 =>  '0' );

  \:48245\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48245\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48245\,
                   R => SYSRESET,
                   S => '0' );

  \=48245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48245\,
                  I0 =>  \48244\,
                  I1 =>  \48242\,
                  I2 =>  \48243\,
                  I3 =>  '0' );

  \=48246\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48246\,
                  I0 =>  \48229\,
                  I1 =>  \48244\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48247\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48247\,
                  I0 =>  \48229\,
                  I1 =>  \48245\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48248\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48248\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48248\,
                   R => '0',
                   S => SYSRESET );

  \=48248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48248\,
                  I0 =>  \48246\,
                  I1 =>  \48249\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48249\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48249\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48249\,
                   R => SYSRESET,
                   S => '0' );

  \=48249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48249\,
                  I0 =>  \48248\,
                  I1 =>  \48247\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPYP\    
  \=48250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48250\,
                  I0 =>  \48239\,
                  I1 =>  \48248\,
                  I2 =>  \48230\,
                  I3 =>  '0' );

  -- Alias \PIPYM\    
  \=48251\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48251\,
                  I0 =>  \48238\,
                  I1 =>  \48248\,
                  I2 =>  \48231\,
                  I3 =>  '0' );

  -- Alias \NOYM\     
  \:48252\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48252\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48252\,
                   R => '0',
                   S => SYSRESET );

  \=48252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48252\,
                  I0 =>  \PIPGY-\,
                  I1 =>  \48253\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48253\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48253\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48253\,
                   R => SYSRESET,
                   S => '0' );

  \=48253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48253\,
                  I0 =>  \48252\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOYP\     
  \:48254\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48254\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48254\,
                   R => '0',
                   S => SYSRESET );

  \=48254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48254\,
                  I0 =>  \PIPGY+\,
                  I1 =>  \48255\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48255\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48255\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48255\,
                   R => SYSRESET,
                   S => '0' );

  \=48255\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48255\,
                  I0 =>  \48254\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MISSY\    
  \:48256\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48256\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48256\,
                   R => '0',
                   S => SYSRESET );

  \=48256\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48256\,
                  I0 =>  \PIPGY+\,
                  I1 =>  \PIPGY-\,
                  I2 =>  \48257\,
                  I3 =>  '0' );

  \:48257\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48257\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48257\,
                   R => SYSRESET,
                   S => '0' );

  \=48257\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48257\,
                  I0 =>  \48256\,
                  I1 =>  \F5ASB2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T7PHS4\   
  \=48258\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48258\,
                  I0 =>  \FUTEXT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ***************************
  -- ***                     ***
  -- ***  A23/2 - INOUT VI.  ***
  -- ***                     ***
  -- ***************************

  \=48301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48301\,
                  I0 =>  \CHWL16/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48302\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48302\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48302\,
                   R => '0',
                   S => SYSRESET );

  \=48302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48302\,
                  I0 =>  \48301\,
                  I1 =>  \48303\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48303\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48303\,
                   R => SYSRESET,
                   S => '0' );

  \=48303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48303\,
                  I0 =>  \48302\,
                  I1 =>  \CCH14\,
                  I2 =>  \48310\,
                  I3 =>  '0' );

  -- Alias \CH1416\   
  \=48304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48304\,
                  I0 =>  \RCH14/\,
                  I1 =>  \48302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUXD\    
  \=48305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48305\,
                  I0 =>  \48302\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48306\,
                  I0 =>  \XB0/\,
                  I1 =>  \48357\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48307\,
                  I0 =>  \48306\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUXDP\   
  \=48308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48308\,
                  I0 =>  \POUT/\,
                  I1 =>  \48307\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUXDM\   
  \=48309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48309\,
                  I0 =>  \48307\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48310\,
                  I0 =>  \48307\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48311\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48312\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48312\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48312\,
                   R => '0',
                   S => SYSRESET );

  \=48312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48312\,
                  I0 =>  \48311\,
                  I1 =>  \48313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48313\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48313\,
                   R => SYSRESET,
                   S => '0' );

  \=48313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48313\,
                  I0 =>  \48312\,
                  I1 =>  \CCH14\,
                  I2 =>  \48320\,
                  I3 =>  '0' );

  -- Alias \CH1414\   
  \=48314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48314\,
                  I0 =>  \RCH14/\,
                  I1 =>  \48312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUYD\    
  \=48315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48315\,
                  I0 =>  \48312\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48316\,
                  I0 =>  \48357\,
                  I1 =>  \XB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48317\,
                  I0 =>  \48316\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUYDP\   
  \=48318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48318\,
                  I0 =>  \POUT/\,
                  I1 =>  \48317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUYDM\   
  \=48319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48319\,
                  I0 =>  \48317\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48320\,
                  I0 =>  \48317\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48321\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48322\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48322\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48322\,
                   R => '0',
                   S => SYSRESET );

  \=48322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48322\,
                  I0 =>  \48321\,
                  I1 =>  \48324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1413\   
  \=48323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48323\,
                  I0 =>  \RCH14/\,
                  I1 =>  \48322\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48324\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48324\,
                   R => SYSRESET,
                   S => '0' );

  \=48324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48324\,
                  I0 =>  \48322\,
                  I1 =>  \CCH14\,
                  I2 =>  \48330\,
                  I3 =>  '0' );

  -- Alias \CDUZD\    
  \=48325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48325\,
                  I0 =>  \48322\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUZDP\   
  \=48326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48326\,
                  I0 =>  \POUT/\,
                  I1 =>  \48328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48327\,
                  I0 =>  \48357\,
                  I1 =>  \XB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48328\,
                  I0 =>  \48327\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUZDM\   
  \=48329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48329\,
                  I0 =>  \48328\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48330\,
                  I0 =>  \48328\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48331\,
                  I0 =>  \WCH14/\,
                  I1 =>  \CHWL12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48332\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48332\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48332\,
                   R => '0',
                   S => SYSRESET );

  \=48332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48332\,
                  I0 =>  \48331\,
                  I1 =>  \48333\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48333\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48333\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48333\,
                   R => SYSRESET,
                   S => '0' );

  \=48333\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48333\,
                  I0 =>  \48332\,
                  I1 =>  \CCH14\,
                  I2 =>  \48340\,
                  I3 =>  '0' );

  -- Alias \CH1412\   
  \=48334\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48334\,
                  I0 =>  \RCH14/\,
                  I1 =>  \48332\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TRUND\    
  \=48335\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48335\,
                  I0 =>  \48332\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TRNDP\    
  \=48336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48336\,
                  I0 =>  \POUT/\,
                  I1 =>  \48338\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48337\,
                  I0 =>  \48357\,
                  I1 =>  \XB3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48338\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48338\,
                  I0 =>  \48337\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \TRNDM\    
  \=48339\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48339\,
                  I0 =>  \48338\,
                  I1 =>  \MOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48340\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48340\,
                  I0 =>  \48338\,
                  I1 =>  \ZOUT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48341\,
                  I0 =>  \CHWL11/\,
                  I1 =>  \WCH14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48342\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48342\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48342\,
                   R => '0',
                   S => SYSRESET );

  \=48342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48342\,
                  I0 =>  \48341\,
                  I1 =>  \48343\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48343\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48343\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48343\,
                   R => SYSRESET,
                   S => '0' );

  \=48343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48343\,
                  I0 =>  \48342\,
                  I1 =>  \CCH14\,
                  I2 =>  \48350\,
                  I3 =>  '0' );

  -- Alias \CH1411\   
  \=48344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48344\,
                  I0 =>  \RCH14/\,
                  I1 =>  \48342\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHAFTD\   
  \=48345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48345\,
                  I0 =>  \48342\,
                  I1 =>  \F5ASB2/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48346\,
                  I0 =>  \48357\,
                  I1 =>  \XB4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48347\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48347\,
                  I0 =>  \48346\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHFTDP\   
  \=48348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48348\,
                  I0 =>  \48351\,
                  I1 =>  \48347\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SHFTDM\   
  \=48349\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48349\,
                  I0 =>  \48347\,
                  I1 =>  \48353\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48350\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48350\,
                  I0 =>  \48347\,
                  I1 =>  \48355\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \POUT/\    
  \=48351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48351\,
                  I0 =>  \POUT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MOUT/\    
  \=48353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48353\,
                  I0 =>  \MOUT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ZOUT/\    
  \=48355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48355\,
                  I0 =>  \ZOUT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48357\,
                  I0 =>  \OCTAD5\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T7PHS4/\  
  \=48358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48358\,
                  I0 =>  \T7PHS4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T7PHS4\   
  \=48359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48359\,
                  I0 =>  \T07/\,
                  I1 =>  \PHS4/\,
                  I2 =>  '0',
                  I3 => \&48258\ );

  \=48401\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48401\,
                  I0 =>  \CHWL05/\,
                  I1 =>  \48415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48402\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48402\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48402\,
                   R => '0',
                   S => SYSRESET );

  \=48402\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48402\,
                  I0 =>  \48401\,
                  I1 =>  \48403\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \E5\       
  \:48403\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48403\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48403\,
                   R => SYSRESET,
                   S => '0' );

  \=48403\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48403\,
                  I0 =>  \48402\,
                  I1 =>  '0',
                  I2 =>  \48413\,
                  I3 =>  '0' );

  -- Alias \CH0705\   
  \=48404\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48404\,
                  I0 =>  \48417\,
                  I1 =>  \48402\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48405\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48405\,
                  I0 =>  \CHWL06/\,
                  I1 =>  \48415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48406\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48406\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48406\,
                   R => '0',
                   S => SYSRESET );

  \=48406\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48406\,
                  I0 =>  \48405\,
                  I1 =>  \48407\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \E6\       
  \:48407\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48407\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48407\,
                   R => SYSRESET,
                   S => '0' );

  \=48407\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48407\,
                  I0 =>  \48406\,
                  I1 =>  '0',
                  I2 =>  \48413\,
                  I3 =>  '0' );

  -- Alias \CH0706\   
  \=48408\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48408\,
                  I0 =>  \48417\,
                  I1 =>  \48406\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48409\,
                  I0 =>  \CHWL07/\,
                  I1 =>  \48415\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \E7/\      
  \:48410\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48410\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48410\,
                   R => '0',
                   S => SYSRESET );

  \=48410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48410\,
                  I0 =>  \48409\,
                  I1 =>  \48411\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48411\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48411\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48411\,
                   R => SYSRESET,
                   S => '0' );

  \=48411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48411\,
                  I0 =>  \48410\,
                  I1 =>  '0',
                  I2 =>  \48413\,
                  I3 =>  '0' );

  -- Alias \CH0707\   
  \=48412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48412\,
                  I0 =>  \48417\,
                  I1 =>  \48410\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCH07\    
  \=48413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48413\,
                  I0 =>  \CCHG/\,
                  I1 =>  \XB7/\,
                  I2 =>  \XT0/\,
                  I3 =>  '0' );

  \=48414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48414\,
                  I0 =>  \WCHG/\,
                  I1 =>  \XT0/\,
                  I2 =>  \XB7/\,
                  I3 =>  '0' );

  -- Alias \WCH07/\   
  \=48415\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48415\,
                  I0 =>  \48414\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48416\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48416\,
                  I0 =>  \XT0/\,
                  I1 =>  \XB7/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCH07/\   
  \=48417\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48417\,
                  I0 =>  \48416\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48418\,
                  I0 =>  \CHWL08/\,
                  I1 =>  \WCH11/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48419\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48419\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48419\,
                   R => '0',
                   S => SYSRESET );

  \=48419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48419\,
                  I0 =>  \48418\,
                  I1 =>  \48420\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48420\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48420\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48420\,
                   R => SYSRESET,
                   S => '0' );

  \=48420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48420\,
                  I0 =>  \48419\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1108\   
  \=48421\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48421\,
                  I0 =>  \RCH11/\,
                  I1 =>  \48419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1108\   
  \=48422\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48422\,
                  I0 =>  \48419\,
                  I1 =>  \48419\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48423\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48423\,
                  I0 =>  \WCH11/\,
                  I1 =>  \CHWL13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48424\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48424\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48424\,
                   R => '0',
                   S => SYSRESET );

  \=48424\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48424\,
                  I0 =>  \48423\,
                  I1 =>  \48425\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48425\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48425\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48425\,
                   R => SYSRESET,
                   S => '0' );

  \=48425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48425\,
                  I0 =>  \48424\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1113\   
  \=48426\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48426\,
                  I0 =>  \RCH11/\,
                  I1 =>  \48424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1113\   
  \=48427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48427\,
                  I0 =>  \48424\,
                  I1 =>  \48424\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48428\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48428\,
                  I0 =>  \WCH11/\,
                  I1 =>  \CHWL14/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48429\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48429\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48429\,
                   R => '0',
                   S => SYSRESET );

  \=48429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48429\,
                  I0 =>  \48428\,
                  I1 =>  \48430\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48430\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48430\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48430\,
                   R => SYSRESET,
                   S => '0' );

  \=48430\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48430\,
                  I0 =>  \48429\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1114\   
  \=48431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48431\,
                  I0 =>  \RCH11/\,
                  I1 =>  \48429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1114\   
  \=48432\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48432\,
                  I0 =>  \48429\,
                  I1 =>  \48429\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48433\,
                  I0 =>  \WCH11/\,
                  I1 =>  \CHWL16/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48434\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48434\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48434\,
                   R => '0',
                   S => SYSRESET );

  \=48434\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48434\,
                  I0 =>  \48433\,
                  I1 =>  \48435\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48435\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48435\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48435\,
                   R => SYSRESET,
                   S => '0' );

  \=48435\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48435\,
                  I0 =>  \48434\,
                  I1 =>  \CCH11\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1116\   
  \=48436\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48436\,
                  I0 =>  \RCH11/\,
                  I1 =>  \48434\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1116\   
  \=48437\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48437\,
                  I0 =>  \48434\,
                  I1 =>  \48434\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR09/\  
  \=48438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48438\,
                  I0 =>  \CHAT09\,
                  I1 =>  \CHBT09\,
                  I2 =>  '0',
                  I3 => \&48439\ );

  -- Alias \CHOR09/\  
  \=48439\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48439\,
                  I0 =>  \CH1109\,
                  I1 =>  \CH1209\,
                  I2 =>  \CH3209\,
                  I3 =>  '0' );

  -- Alias \CH09\     
  \=48440\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48440\,
                  I0 =>  \CHOR09/\,
                  I1 =>  \RCHG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48441\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48441\,
                  I0 =>  \CHWL16/\,
                  I1 =>  \WCH12/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48442\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48442\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48442\,
                   R => '0',
                   S => SYSRESET );

  \=48442\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48442\,
                  I0 =>  \48441\,
                  I1 =>  \48443\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48443\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48443\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48443\,
                   R => SYSRESET,
                   S => '0' );

  \=48443\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48443\,
                  I0 =>  \48442\,
                  I1 =>  \CCH12\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1216\   
  \=48444\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48444\,
                  I0 =>  \RCH12/\,
                  I1 =>  \48442\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ISSTDC\   
  \=48445\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48445\,
                  I0 =>  \48442\,
                  I1 =>  \48442\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48446\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48446\,
                  I0 =>  \CHWL16/\,
                  I1 =>  \WCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \T6ON/\    
  \:48447\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48447\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48447\,
                   R => '0',
                   S => SYSRESET );

  \=48447\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48447\,
                  I0 =>  \48446\,
                  I1 =>  \48448\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48448\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48448\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48448\,
                   R => SYSRESET,
                   S => '0' );

  \=48448\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48448\,
                  I0 =>  \48447\,
                  I1 =>  \T6RPT\,
                  I2 =>  \CCH13\,
                  I3 =>  '0' );

  -- Alias \CH1316\   
  \=48449\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48449\,
                  I0 =>  \48447\,
                  I1 =>  \RCH13/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=48450\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48450\,
                  I0 =>  \WCH13/\,
                  I1 =>  \CHWL10/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48451\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \48451\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48451\,
                   R => '0',
                   S => SYSRESET );

  \=48451\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48451\,
                  I0 =>  \48450\,
                  I1 =>  \48452\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:48452\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \48452\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$48452\,
                   R => SYSRESET,
                   S => '0' );

  \=48452\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$48452\,
                  I0 =>  \48451\,
                  I1 =>  \CCH13\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CH1310\   
  \=48453\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48453\,
                  I0 =>  \RCH13/\,
                  I1 =>  \48451\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ALTEST\   
  \=48454\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48454\,
                  I0 =>  \48451\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHOR10/\  
  \=48456\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48456\,
                  I0 =>  \CHAT10\,
                  I1 =>  \CHBT10\,
                  I2 =>  '0',
                  I3 => \&48457\ );

  -- Alias \CHOR10/\  
  \=48457\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&48457\,
                  I0 =>  \CH1110\,
                  I1 =>  \CH1210\,
                  I2 =>  \CH3210\,
                  I3 =>  '0' );

  -- Alias \CH10\     
  \=48458\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \48458\,
                  I0 =>  \CHOR10/\,
                  I1 =>  \RCHG/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************
  -- ***                      ***
  -- ***  A24/1 - INOUT VII.  ***
  -- ***                      ***
  -- ****************************

  \=49101\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49101\,
                  I0 =>  \A16/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49102\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49102\,
                  I0 =>  \A15/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49103\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49103\,
                  I0 =>  \49101\,
                  I1 =>  \A15/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49104\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49104\,
                  I0 =>  \A16/\,
                  I1 =>  \49102\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49105\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49105\,
                  I0 =>  \49103\,
                  I1 =>  \49104\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49106\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49106\,
                  I0 =>  \49105\,
                  I1 =>  \NISQ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49107\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49107\,
                  I0 =>  \49103\,
                  I1 =>  \49104\,
                  I2 =>  \NISQ/\,
                  I3 =>  '0' );

  \:49108\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49108\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49108\,
                   R => '0',
                   S => SYSRESET );

  \=49108\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49108\,
                  I0 =>  \49106\,
                  I1 =>  \49109\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OVNHRP\   
  \=49109\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49109\,
                  I0 =>  \49108\,
                  I1 =>  \49107\,
                  I2 =>  \MP3\,
                  I3 =>  '0' );

  \=49110\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49110\,
                  I0 =>  \T02/\,
                  I1 =>  \CA6/\,
                  I2 =>  \XB7/\,
                  I3 =>  '0' );

  \=49111\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49111\,
                  I0 =>  \49110\,
                  I1 =>  \49112\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49112\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49112\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49112\,
                   R => '0',
                   S => SYSRESET );

  \=49112\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49112\,
                  I0 =>  \49111\,
                  I1 =>  \F17B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49113\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49113\,
                  I0 =>  \F17A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WATCHP\   
  \=49114\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49114\,
                  I0 =>  \SB2/\,
                  I1 =>  \49112\,
                  I2 =>  \49113\,
                  I3 =>  '0' );

  \=49115\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49115\,
                  I0 =>  \49113\,
                  I1 =>  \SB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WATCH/\   
  \:49116\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49116\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49116\,
                   R => '0',
                   S => SYSRESET );

  \=49116\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49116\,
                  I0 =>  \49114\,
                  I1 =>  \49117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WATCH\    
  \=49117\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49117\,
                  I0 =>  \49116\,
                  I1 =>  \49115\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWATCH/\  
  \=49118\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49118\,
                  I0 =>  \49117\,
                  I1 =>  \49117\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49120\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49120\,
                  I0 =>  \DKCTR5\,
                  I1 =>  \DKCTR4\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \HIGH0/\   
  \=49121\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49121\,
                  I0 =>  \49120\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49123\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49123\,
                  I0 =>  \DKCTR5\,
                  I1 =>  \DKCTR4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \HIGH1/\   
  \=49124\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49124\,
                  I0 =>  \49123\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49126\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49126\,
                  I0 =>  \DKCTR4\,
                  I1 =>  \DKCTR5/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \HIGH2/\   
  \=49127\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49127\,
                  I0 =>  \49126\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49129\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49129\,
                  I0 =>  \DKCTR5/\,
                  I1 =>  \DKCTR4/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \HIGH3/\   
  \=49130\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49130\,
                  I0 =>  \49129\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49132\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49132\,
                  I0 =>  \RCH/\,
                  I1 =>  \RT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCHG/\    
  \=49133\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49133\,
                  I0 =>  \49132\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49136\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49136\,
                  I0 =>  \WT/\,
                  I1 =>  \WCH/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \WCHG/\    
  \=49137\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49137\,
                  I0 =>  \49136\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49140\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49140\,
                  I0 =>  \WCH/\,
                  I1 =>  \CT/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CCHG/\    
  \=49141\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49141\,
                  I0 =>  \49140\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL01/\  
  \=49143\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49143\,
                  I0 =>  \WL01\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL02/\  
  \=49145\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49145\,
                  I0 =>  \WL02\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL03/\  
  \=49147\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49147\,
                  I0 =>  \WL03\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL04/\  
  \=49149\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49149\,
                  I0 =>  \WL04\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL05/\  
  \=49151\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49151\,
                  I0 =>  \WL05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL06/\  
  \=49153\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49153\,
                  I0 =>  \WL06\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL07/\  
  \=49155\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49155\,
                  I0 =>  \WL07\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL08/\  
  \=49157\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49157\,
                  I0 =>  \WL08\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL09/\  
  \=49159\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49159\,
                  I0 =>  \WL09\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49201\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49201\,
                  I0 =>  \FS04\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49202\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49202\,
                  I0 =>  \F03B/\,
                  I1 =>  \49201\,
                  I2 =>  \FS05\,
                  I3 =>  '0' );

  -- Alias \PIPPLS/\  
  \=49203\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49203\,
                  I0 =>  \49202\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPASW\   
  \=49204\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49204\,
                  I0 =>  \49203\,
                  I1 =>  \49226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS05/\    
  \=49205\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49205\,
                  I0 =>  \FS05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPDAT\   
  \=49206\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49206\,
                  I0 =>  \49203\,
                  I1 =>  \49228\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49207\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49207\,
                  I0 =>  \SB4\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPINT\   
  \=49208\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49208\,
                  I0 =>  \49203\,
                  I1 =>  \49207\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \800SET\   
  \=49209\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49209\,
                  I0 =>  \F07A/\,
                  I1 =>  \49226\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \800RST\   
  \=49210\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49210\,
                  I0 =>  \49226\,
                  I1 =>  \F07B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3200A\    
  \=49211\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49211\,
                  I0 =>  \F05A/\,
                  I1 =>  \49224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3200B\    
  \=49212\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49212\,
                  I0 =>  \F05B/\,
                  I1 =>  \49224\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3200C\    
  \=49213\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49213\,
                  I0 =>  \FS05\,
                  I1 =>  \49224\,
                  I2 =>  \49214\,
                  I3 =>  '0' );

  \=49214\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49214\,
                  I0 =>  \F04B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \3200D\    
  \=49215\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49215\,
                  I0 =>  \49214\,
                  I1 =>  \49224\,
                  I2 =>  \49205\,
                  I3 =>  '0' );

  \=49216\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49216\,
                  I0 =>  \F02B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \12KPPS\   
  \=49217\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49217\,
                  I0 =>  \FS03\,
                  I1 =>  \49216\,
                  I2 =>  \49224\,
                  I3 =>  '0' );

  -- Alias \RRRST\    
  \=49218\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49218\,
                  I0 =>  \F05B/\,
                  I1 =>  \SB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \LRRST\    
  \=49219\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49219\,
                  I0 =>  \F05B/\,
                  I1 =>  \SB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \25KPPS\   
  \=49220\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49220\,
                  I0 =>  \49224\,
                  I1 =>  \FS02\,
                  I2 =>  \49221\,
                  I3 =>  '0' );

  \=49221\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49221\,
                  I0 =>  \F01B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49222\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49222\,
                  I0 =>  \F01A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUCLK\   
  \=49223\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49223\,
                  I0 =>  \49222\,
                  I1 =>  \SB0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB0/\     
  \=49224\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49224\,
                  I0 =>  \SB0\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB1/\     
  \=49226\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49226\,
                  I0 =>  \SB1\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \SB2/\     
  \=49228\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49228\,
                  I0 =>  \SB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F05A/\    
  \=49230\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49230\,
                  I0 =>  \F05A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F05B/\    
  \=49232\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49232\,
                  I0 =>  \F05B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07B/\    
  \=49234\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49234\,
                  I0 =>  \F07B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL10/\  
  \=49235\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49235\,
                  I0 =>  \WL10\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NISQ\     
  \=49237\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49237\,
                  I0 =>  \NISQ/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MNISQ\    
  \=49238\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49238\,
                  I0 =>  \NISQ/\,
                  I1 =>  \NISQ/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MON800\   
  \=49239\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49239\,
                  I0 =>  \FS07A\,
                  I1 =>  \FS07A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49240\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49240\,
                  I0 =>  \XB4/\,
                  I1 =>  \XT0/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCHAT/\   
  \=49241\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49241\,
                  I0 =>  \49240\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49244\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49244\,
                  I0 =>  \XT0/\,
                  I1 =>  \XB3/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RCHBT/\   
  \=49245\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49245\,
                  I0 =>  \49244\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49248\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49248\,
                  I0 =>  \FS07A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ELSNCN\   
  \=49249\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49249\,
                  I0 =>  \49248\,
                  I1 =>  \49248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ELSNCM\   
  \=49250\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49250\,
                  I0 =>  \49248\,
                  I1 =>  \49248\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1110\   
  \=49252\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49252\,
                  I0 =>  \FF1110/\,
                  I1 =>  \FF1110/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1111\   
  \=49253\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49253\,
                  I0 =>  \FF1111/\,
                  I1 =>  \FF1111/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OT1112\   
  \=49254\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49254\,
                  I0 =>  \FF1112/\,
                  I1 =>  \FF1112/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- ****************************
  -- ***                      ***
  -- ***  A24/2 - INOUT VII.  ***
  -- ***                      ***
  -- ****************************

  \=49301\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49301\,
                  I0 =>  \PIPGZ+\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49302\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49302\,
                  I0 =>  \PIPGZ-\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOZM\     
  \:49303\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49303\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49303\,
                   R => '0',
                   S => SYSRESET );

  \=49303\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49303\,
                  I0 =>  \PIPGZ-\,
                  I1 =>  \49304\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49304\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49304\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49304\,
                   R => SYSRESET,
                   S => '0' );

  \=49304\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49304\,
                  I0 =>  \49303\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NOZP\     
  \:49305\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49305\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49305\,
                   R => '0',
                   S => SYSRESET );

  \=49305\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49305\,
                  I0 =>  \PIPGZ+\,
                  I1 =>  \49306\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49306\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49306\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49306\,
                   R => SYSRESET,
                   S => '0' );

  \=49306\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49306\,
                  I0 =>  \49305\,
                  I1 =>  \F18AX\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MISSZ\    
  \:49307\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49307\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49307\,
                   R => '0',
                   S => SYSRESET );

  \=49307\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49307\,
                  I0 =>  \PIPGZ+\,
                  I1 =>  \PIPGZ-\,
                  I2 =>  \49308\,
                  I3 =>  '0' );

  \:49308\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49308\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49308\,
                   R => SYSRESET,
                   S => '0' );

  \=49308\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49308\,
                  I0 =>  \49307\,
                  I1 =>  \F5ASB2\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \BOTHZ\    
  \=49309\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49309\,
                  I0 =>  \49301\,
                  I1 =>  \49302\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49310\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49310\,
                  I0 =>  \49302\,
                  I1 =>  \49328\,
                  I2 =>  \49317\,
                  I3 =>  '0' );

  \=49311\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49311\,
                  I0 =>  \49316\,
                  I1 =>  \49328\,
                  I2 =>  \49301\,
                  I3 =>  '0' );

  \:49312\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49312\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49312\,
                   R => '0',
                   S => SYSRESET );

  \=49312\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49312\,
                  I0 =>  \49310\,
                  I1 =>  \49313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49313\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49313\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49313\,
                   R => SYSRESET,
                   S => '0' );

  \=49313\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49313\,
                  I0 =>  \49312\,
                  I1 =>  \49311\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49314\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49314\,
                  I0 =>  \49318\,
                  I1 =>  \49312\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49315\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49315\,
                  I0 =>  \49318\,
                  I1 =>  \49313\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49316\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49316\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49316\,
                   R => '0',
                   S => SYSRESET );

  \=49316\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49316\,
                  I0 =>  \49314\,
                  I1 =>  \49317\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49317\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49317\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49317\,
                   R => SYSRESET,
                   S => '0' );

  \=49317\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49317\,
                  I0 =>  \49316\,
                  I1 =>  \49315\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49318\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49318\,
                  I0 =>  \F5ASB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49319\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49319\,
                  I0 =>  \49317\,
                  I1 =>  \49328\,
                  I2 =>  \49301\,
                  I3 =>  '0' );

  \=49320\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49320\,
                  I0 =>  \49316\,
                  I1 =>  \49328\,
                  I2 =>  \49302\,
                  I3 =>  '0' );

  \=49321\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49321\,
                  I0 =>  \49317\,
                  I1 =>  \49327\,
                  I2 =>  \49302\,
                  I3 =>  '0' );

  \=49322\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49322\,
                  I0 =>  \49316\,
                  I1 =>  \49327\,
                  I2 =>  \49301\,
                  I3 =>  '0' );

  \:49323\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49323\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49323\,
                   R => '0',
                   S => SYSRESET );

  \=49323\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49323\,
                  I0 =>  \49319\,
                  I1 =>  \49320\,
                  I2 =>  \49324\,
                  I3 =>  '0' );

  \:49324\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49324\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49324\,
                   R => SYSRESET,
                   S => '0' );

  \=49324\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49324\,
                  I0 =>  \49323\,
                  I1 =>  \49321\,
                  I2 =>  \49322\,
                  I3 =>  '0' );

  \=49325\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49325\,
                  I0 =>  \49318\,
                  I1 =>  \49323\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49326\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49326\,
                  I0 =>  \49318\,
                  I1 =>  \49324\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49327\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49327\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49327\,
                   R => '0',
                   S => SYSRESET );

  \=49327\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49327\,
                  I0 =>  \49325\,
                  I1 =>  \49328\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49328\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49328\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49328\,
                   R => SYSRESET,
                   S => '0' );

  \=49328\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49328\,
                  I0 =>  \49327\,
                  I1 =>  \49326\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PIPZP\    
  \=49329\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49329\,
                  I0 =>  \49317\,
                  I1 =>  \49327\,
                  I2 =>  \49301\,
                  I3 =>  '0' );

  -- Alias \PIPZM\    
  \=49330\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49330\,
                  I0 =>  \49316\,
                  I1 =>  \49327\,
                  I2 =>  \49302\,
                  I3 =>  '0' );

  -- Alias \CNTRSB/\  
  \=49331\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49331\,
                  I0 =>  \SB2\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \RSCT/\    
  \=49332\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49332\,
                  I0 =>  \RSCT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWCH\     
  \=49334\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49334\,
                  I0 =>  \WCH/\,
                  I1 =>  \WCH/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRCH\     
  \=49335\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49335\,
                  I0 =>  \RCH/\,
                  I1 =>  \RCH/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \US2SG\    
  \=49336\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49336\,
                  I0 =>  \RUSG/\,
                  I1 =>  \SUMA15/\,
                  I2 =>  \SUMB15/\,
                  I3 =>  '0' );

  -- Alias \U2BBKG/\  
  \=49337\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49337\,
                  I0 =>  \U2BBK\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \OUTCOM\   
  \=49339\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49339\,
                  I0 =>  \FF1109/\,
                  I1 =>  \FF1109/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49341\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49341\,
                  I0 =>  \FS07/\,
                  I1 =>  \FS08/\,
                  I2 =>  \49348\,
                  I3 =>  '0' );

  \=49342\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49342\,
                  I0 =>  \49341\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GTSET\    
  \=49343\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49343\,
                  I0 =>  \FS06/\,
                  I1 =>  \F05B/\,
                  I2 =>  \49342\,
                  I3 =>  '0' );

  -- Alias \GTSET/\   
  \=49344\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49344\,
                  I0 =>  \49343\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \GTRST\    
  \=49345\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49345\,
                  I0 =>  \49342\,
                  I1 =>  \F05B/\,
                  I2 =>  \FS06\,
                  I3 =>  '0' );

  -- Alias \GTONE\    
  \=49346\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49346\,
                  I0 =>  \FS06\,
                  I1 =>  \F05B/\,
                  I2 =>  \FS07A\,
                  I3 => \&49347\ );

  -- Alias \49346\    
  \=49347\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49347\,
                  I0 =>  \FS08\,
                  I1 =>  \FS09\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FS09/\    
  \=49348\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49348\,
                  I0 =>  \FS09\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49351\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49351\,
                  I0 =>  \F08B/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F09D\     
  \=49352\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49352\,
                  I0 =>  \49351\,
                  I1 =>  \49348\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F09A/\    
  \=49353\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49353\,
                  I0 =>  \F09A\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CI\       
  \=49354\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49354\,
                  I0 =>  \CI/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49355\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49355\,
                  I0 =>  \FS07/\,
                  I1 =>  \F06B/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49356\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49356\,
                  I0 =>  \F06B/\,
                  I1 =>  \FS07A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07D/\    
  \=49357\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49357\,
                  I0 =>  \49355\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F07C/\    
  \=49358\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49358\,
                  I0 =>  \49356\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=49359\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49359\,
                  I0 =>  \49358\,
                  I1 =>  \SB1/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F7CSB1/\  
  \=49360\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49360\,
                  I0 =>  \49359\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FLASH\    
  \=49409\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49409\,
                  I0 =>  \FS17\,
                  I1 =>  \FS16\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \FLASH/\   
  \=49410\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49410\,
                  I0 =>  \49409\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \ONE\      
  \=49411\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49411\,
                  I0 =>  '0',
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:49412\    : FDRSE generic map( INIT=>'0' ) port map(
                   Q => \49412\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49412\,
                   R => SYSRESET,
                   S => '0' );

  \=49412\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49412\,
                  I0 =>  \T08\,
                  I1 =>  \49413\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CDUSTB/\  
  \:49413\    : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \49413\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$49413\,
                   R => '0',
                   S => SYSRESET );

  \=49413\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$49413\,
                  I0 =>  \49412\,
                  I1 =>  \T06\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \PHS3/\    
  \=49414\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49414\,
                  I0 =>  \CT\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F04B/\    
  \=49418\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49418\,
                  I0 =>  \F04B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \IC11/\    
  \=49419\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49419\,
                  I0 =>  \IC11\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \F05D\     
  \=49420\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49420\,
                  I0 =>  \49418\,
                  I1 =>  \FS05/\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL11/\  
  \=49425\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49425\,
                  I0 =>  \WL11\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL12/\  
  \=49427\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49427\,
                  I0 =>  \WL12\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL13/\  
  \=49429\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49429\,
                  I0 =>  \WL13\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL14/\  
  \=49431\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49431\,
                  I0 =>  \WL14\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CHWL16/\  
  \=49433\    : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \49433\,
                  I0 =>  \WL16\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \CTPLS/\   
  \=49435\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49435\,
                  I0 =>  \T1P\,
                  I1 =>  \T2P\,
                  I2 =>  \T3P\,
                  I3 => \&49436\ );

  -- Alias \CTPLS/\   
  \=49436\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49436\,
                  I0 =>  \T4P\,
                  I1 =>  \T5P\,
                  I2 =>  \T6P\,
                  I3 => \&49437\ );

  -- Alias \CTPLS/\   
  \=49437\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49437\,
                  I0 =>  \CDUXP\,
                  I1 =>  \CDUXM\,
                  I2 =>  \CDUYP\,
                  I3 => \&49438\ );

  -- Alias \CTPLS/\   
  \=49438\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49438\,
                  I0 =>  \CDUYM\,
                  I1 =>  \CDUZP\,
                  I2 =>  \CDUZM\,
                  I3 => \&49439\ );

  -- Alias \CTPLS/\   
  \=49439\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49439\,
                  I0 =>  \TRNP\,
                  I1 =>  \TRNM\,
                  I2 =>  \SHAFTP\,
                  I3 => \&49440\ );

  -- Alias \CTPLS/\   
  \=49440\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49440\,
                  I0 =>  \SHAFTM\,
                  I1 =>  \PIPXP\,
                  I2 =>  \PIPXM\,
                  I3 => \&49441\ );

  -- Alias \CTPLS/\   
  \=49441\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49441\,
                  I0 =>  \PIPYP\,
                  I1 =>  \PIPYM\,
                  I2 =>  \PIPZP\,
                  I3 => \&49442\ );

  -- Alias \CTPLS/\   
  \=49442\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49442\,
                  I0 =>  \PIPZM\,
                  I1 =>  \BMAGXP\,
                  I2 =>  \BMAGXM\,
                  I3 => \&49443\ );

  -- Alias \CTPLS/\   
  \=49443\    : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&49443\,
                  I0 =>  \BMAGYP\,
                  I1 =>  \BMAGYM\,
                  I2 =>  \BMAGZP\,
                  I3 =>  '0' );

  -- ***********************************
  -- ***                             ***
  -- ***  CH77/1 - RESTART MONITOR.  ***
  -- ***                             ***
  -- ***********************************

  \=1A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \1A\,
                  I0 =>  \MWL01\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=2A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \2A\,
                  I0 =>  \MWL02\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=2B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \2B\,
                  I0 =>  \MWL03\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=3A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \3A\,
                  I0 =>  \MWL04\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=3B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \3B\,
                  I0 =>  \MWL05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=4A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \4A\,
                  I0 =>  \MWL06\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=4B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \4B\,
                  I0 =>  \MT01\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=5A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \5A\,
                  I0 =>  \MWSG\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=6A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \6A\,
                  I0 =>  \MT12\,
                  I1 =>  \6B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:6B\       : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \6B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$6B\,
                   R => '0',
                   S => SYSRESET );

  \=6B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$6B\,
                  I0 =>  \6A\,
                  I1 =>  \1B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=7A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \7A\,
                  I0 =>  \MWCH\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=8A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \8A\,
                  I0 =>  \MRCH\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=1B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \1B\,
                  I0 =>  \1A\,
                  I1 =>  \2A\,
                  I2 =>  \2B\,
                  I3 => \&10A\ );

  -- Alias \1B\       
  \=10A\      : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&10A\,
                  I0 =>  \3A\,
                  I1 =>  \3B\,
                  I2 =>  \4A\,
                  I3 => \&10B\ );

  -- Alias \1B\       
  \=10B\      : LUT4_L generic map( INIT=>X"FFFE" ) port map(
                  LO => \&10B\,
                  I0 =>  \4B\,
                  I1 =>  \5A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=5B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \5B\,
                  I0 =>  \6B\,
                  I1 =>  \7A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=8B\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \8B\,
                  I0 =>  \6B\,
                  I1 =>  \8A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=9A\       : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \9A\,
                  I0 =>  \8B\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=12A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \12A\,
                  I0 =>  \MT05\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=11A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \11A\,
                  I0 =>  \MPAL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=13A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \13A\,
                  I0 =>  \MPAL/\,
                  I1 =>  \12A\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=14A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \14A\,
                  I0 =>  \MTCAL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=15A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \15A\,
                  I0 =>  \MRPTAL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=16A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \16A\,
                  I0 =>  \MWATCH/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=17A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \17A\,
                  I0 =>  \MVFAIL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=18A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \18A\,
                  I0 =>  \MCTRAL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=19A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \19A\,
                  I0 =>  \MSCAFL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \=20A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \20A\,
                  I0 =>  \MSCDBL/\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  \:11B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \11B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$11B\,
                   R => '0',
                   S => SYSRESET );

  \=11B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$11B\,
                  I0 =>  \11A\,
                  I1 =>  \21B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=21B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \21B\,
                  I0 =>  \11B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:13B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \13B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$13B\,
                   R => '0',
                   S => SYSRESET );

  \=13B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$13B\,
                  I0 =>  \13A\,
                  I1 =>  \22B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=22B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \22B\,
                  I0 =>  \13B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:14B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \14B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$14B\,
                   R => '0',
                   S => SYSRESET );

  \=14B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$14B\,
                  I0 =>  \14A\,
                  I1 =>  \23B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=23B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \23B\,
                  I0 =>  \14B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:15B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \15B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$15B\,
                   R => '0',
                   S => SYSRESET );

  \=15B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$15B\,
                  I0 =>  \15A\,
                  I1 =>  \24B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=24B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \24B\,
                  I0 =>  \15B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:16B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \16B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$16B\,
                   R => '0',
                   S => SYSRESET );

  \=16B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$16B\,
                  I0 =>  \16A\,
                  I1 =>  \25B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=25B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \25B\,
                  I0 =>  \16B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:17B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \17B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$17B\,
                   R => '0',
                   S => SYSRESET );

  \=17B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$17B\,
                  I0 =>  \17A\,
                  I1 =>  \26B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=26B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \26B\,
                  I0 =>  \17B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:18B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \18B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$18B\,
                   R => '0',
                   S => SYSRESET );

  \=18B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$18B\,
                  I0 =>  \18A\,
                  I1 =>  \27B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=27B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \27B\,
                  I0 =>  \18B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:19B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \19B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$19B\,
                   R => '0',
                   S => SYSRESET );

  \=19B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$19B\,
                  I0 =>  \19A\,
                  I1 =>  \28B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=28B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \28B\,
                  I0 =>  \19B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \:20B\      : FDRSE generic map( INIT=>'1' ) port map(
                   Q => \20B\,
                   C => SYSCLOCK,
                  CE => '1',
                   D => \$20B\,
                   R => '0',
                   S => SYSRESET );

  \=20B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO => \$20B\,
                  I0 =>  \20A\,
                  I1 =>  \29B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  \=29B\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \29B\,
                  I0 =>  \20B\,
                  I1 =>  \5B\,
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT01\    
  \=21A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \21A\,
                  I0 =>  '0',
                  I1 =>  \11B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT02\    
  \=22A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \22A\,
                  I0 =>  '0',
                  I1 =>  \13B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT03\    
  \=23A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \23A\,
                  I0 =>  '0',
                  I1 =>  \14B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT04\    
  \=24A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \24A\,
                  I0 =>  '0',
                  I1 =>  \15B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT05\    
  \=25A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \25A\,
                  I0 =>  '0',
                  I1 =>  \16B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT06\    
  \=26A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \26A\,
                  I0 =>  '0',
                  I1 =>  \17B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT07\    
  \=27A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \27A\,
                  I0 =>  '0',
                  I1 =>  \18B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT08\    
  \=28A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \28A\,
                  I0 =>  '0',
                  I1 =>  \19B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \MDT09\    
  \=29A\      : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \29A\,
                  I0 =>  '0',
                  I1 =>  \20B\,
                  I2 =>  \9A\,
                  I3 =>  '0' );

  -- Alias \DERHI\    
  \=PULLD01\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD01\,
                  I0 =>  '0',
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DERLO\    
  \=PULLD02\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD02\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT10\    
  \=PULLD03\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD03\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT11\    
  \=PULLD04\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD04\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT12\    
  \=PULLD05\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD05\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT13\    
  \=PULLD06\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD06\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT14\    
  \=PULLD07\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD07\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT15\    
  \=PULLD08\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD08\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MDT16\    
  \=PULLD09\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD09\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MNHSBF\   
  \=PULLD10\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD10\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MNHNC\    
  \=PULLD11\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD11\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MNHRPT\   
  \=PULLD12\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD12\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MTCSAI\   
  \=PULLD13\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD13\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSTRT\    
  \=PULLD14\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD14\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSTP\     
  \=PULLD15\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD15\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MSBSTP\   
  \=PULLD16\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD16\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MRDCH\    
  \=PULLD17\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD17\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MLDCH\    
  \=PULLD18\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD18\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MONPAR\   
  \=PULLD19\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD19\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MONWBK\   
  \=PULLD20\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD20\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MLOAD\    
  \=PULLD21\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD21\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MREAD\    
  \=PULLD22\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD22\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \NHALGA\   
  \=PULLD23\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD23\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DOSCAL\   
  \=PULLD24\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD24\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \DBLTST\   
  \=PULLD25\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD25\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MAMU\     
  \=PULLD26\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLD26\,
                  I0 =>  \DERHI\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 =>  '0' );

  -- Alias \MWL01\    
  \=PULLU01\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU01\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51153\ );

  -- Alias \MWL02\    
  \=PULLU02\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU02\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51253\ );

  -- Alias \MWL03\    
  \=PULLU03\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU03\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51453\ );

  -- Alias \MWL04\    
  \=PULLU04\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU04\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51353\ );

  -- Alias \MWL05\    
  \=PULLU05\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU05\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52153\ );

  -- Alias \MWL06\    
  \=PULLU06\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU06\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52253\ );

  -- Alias \MT01\     
  \=PULLU07\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU07\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37404\ );

  -- Alias \MWSG\     
  \=PULLU08\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU08\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33241\ );

  -- Alias \MT12\     
  \=PULLU09\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU09\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37454\ );

  -- Alias \MWCH\     
  \=PULLU10\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU10\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49334\ );

  -- Alias \MRCH\     
  \=PULLU11\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU11\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49335\ );

  -- Alias \MPAL/\    
  \=PULLU12\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU12\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&34252\ );

  -- Alias \MT05\     
  \=PULLU13\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU13\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37422\ );

  -- Alias \MTCAL/\   
  \=PULLU14\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU14\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41127\ );

  -- Alias \MRPTAL/\  
  \=PULLU15\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU15\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41114\ );

  -- Alias \MWATCH/\  
  \=PULLU16\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU16\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49118\ );

  -- Alias \MVFAIL/\  
  \=PULLU17\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU17\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41207\ );

  -- Alias \MCTRAL/\  
  \=PULLU18\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU18\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41144\ );

  -- Alias \MSCAFL/\  
  \=PULLU19\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU19\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41222\ );

  -- Alias \MSCDBL/\  
  \=PULLU20\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU20\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&34254\ );

  -- Alias \GEM01\    
  \=PULLU21\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU21\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51150\ );

  -- Alias \GEM02\    
  \=PULLU22\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU22\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51250\ );

  -- Alias \GEM03\    
  \=PULLU23\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU23\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51450\ );

  -- Alias \GEM04\    
  \=PULLU24\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU24\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&51350\ );

  -- Alias \GEM05\    
  \=PULLU25\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU25\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52150\ );

  -- Alias \GEM06\    
  \=PULLU26\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU26\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52250\ );

  -- Alias \GEM07\    
  \=PULLU27\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU27\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52450\ );

  -- Alias \GEM08\    
  \=PULLU28\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU28\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52350\ );

  -- Alias \GEM09\    
  \=PULLU29\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU29\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53150\ );

  -- Alias \GEM10\    
  \=PULLU30\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU30\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53250\ );

  -- Alias \GEM11\    
  \=PULLU31\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU31\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53450\ );

  -- Alias \GEM12\    
  \=PULLU32\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU32\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53350\ );

  -- Alias \GEM13\    
  \=PULLU33\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU33\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54150\ );

  -- Alias \GEM14\    
  \=PULLU34\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU34\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54250\ );

  -- Alias \GEM16\    
  \=PULLU35\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU35\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54350\ );

  -- Alias \GEMP\     
  \=PULLU36\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU36\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&34243\ );

  -- Alias \SBE\      
  \=PULLU37\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU37\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42251\ );

  -- Alias \SBF\      
  \=PULLU38\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU38\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42121\ );

  -- Alias \ZID\      
  \=PULLU39\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU39\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42222\ );

  -- Alias \REX\      
  \=PULLU40\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU40\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42237\ );

  -- Alias \REY\      
  \=PULLU41\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU41\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42236\ );

  -- Alias \WEX\      
  \=PULLU42\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU42\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42207\ );

  -- Alias \WEY\      
  \=PULLU43\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU43\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42208\ );

  -- Alias \CLROPE\   
  \=PULLU44\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU44\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52162\ );

  -- Alias \FILTIN\   
  \=PULLU45\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU45\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41216\ );

  -- Alias \HIMOD\    
  \=PULLU46\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU46\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35449\ );

  -- Alias \IHENV\    
  \=PULLU47\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU47\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42108\ );

  -- Alias \IL01\     
  \=PULLU48\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU48\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40226\ );

  -- Alias \IL01/\    
  \=PULLU49\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU49\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40227\ );

  -- Alias \IL02\     
  \=PULLU50\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU50\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40228\ );

  -- Alias \IL02/\    
  \=PULLU51\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU51\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40229\ );

  -- Alias \IL03\     
  \=PULLU52\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU52\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40230\ );

  -- Alias \IL03/\    
  \=PULLU53\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU53\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40231\ );

  -- Alias \IL04\     
  \=PULLU54\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU54\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40232\ );

  -- Alias \IL04/\    
  \=PULLU55\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU55\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40233\ );

  -- Alias \IL05\     
  \=PULLU56\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU56\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40234\ );

  -- Alias \IL05/\    
  \=PULLU57\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU57\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40235\ );

  -- Alias \IL06\     
  \=PULLU58\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU58\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40236\ );

  -- Alias \IL06/\    
  \=PULLU59\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU59\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40237\ );

  -- Alias \IL07\     
  \=PULLU60\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU60\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40238\ );

  -- Alias \IL07/\    
  \=PULLU61\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU61\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40239\ );

  -- Alias \ILP\      
  \=PULLU62\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU62\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42446\ );

  -- Alias \ILP/\     
  \=PULLU63\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU63\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42447\ );

  -- Alias \LOMOD\    
  \=PULLU64\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU64\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35429\ );

  -- Alias \MBR1\     
  \=PULLU65\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU65\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36260\ );

  -- Alias \MBR2\     
  \=PULLU66\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU66\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36262\ );

  -- Alias \MGOJAM\   
  \=PULLU67\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU67\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37251\ );

  -- Alias \MGP/\     
  \=PULLU68\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU68\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&34241\ );

  -- Alias \MIIP\     
  \=PULLU69\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU69\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30112\ );

  -- Alias \MINHL\    
  \=PULLU70\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU70\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30111\ );

  -- Alias \MINKL\    
  \=PULLU71\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU71\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&32253\ );

  -- Alias \MNISQ\    
  \=PULLU72\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU72\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49238\ );

  -- Alias \MON800\   
  \=PULLU73\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU73\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49239\ );

  -- Alias \MONWT\    
  \=PULLU74\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU74\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37136\ );

  -- Alias \MOSCAL/\  
  \=PULLU75\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU75\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41231\ );

  -- Alias \MPIPAL/\  
  \=PULLU76\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU76\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41106\ );

  -- Alias \MRAG\     
  \=PULLU77\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU77\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33326\ );

  -- Alias \MREQIN\   
  \=PULLU78\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU78\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&32230\ );

  -- Alias \MRGG\     
  \=PULLU79\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU79\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33320\ );

  -- Alias \MRLG\     
  \=PULLU80\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU80\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33335\ );

  -- Alias \MRSC\     
  \=PULLU81\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU81\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36459\ );

  -- Alias \MRULOG\   
  \=PULLU82\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU82\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33347\ );

  -- Alias \MSP\      
  \=PULLU83\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU83\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&34244\ );

  -- Alias \MSQ10\    
  \=PULLU84\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU84\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30140\ );

  -- Alias \MSQ11\    
  \=PULLU85\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU85\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30139\ );

  -- Alias \MSQ12\    
  \=PULLU86\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU86\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30138\ );

  -- Alias \MSQ13\    
  \=PULLU87\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU87\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30028\ );

  -- Alias \MSQ14\    
  \=PULLU88\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU88\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30025\ );

  -- Alias \MSQ16\    
  \=PULLU89\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU89\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30022\ );

  -- Alias \MSQEXT\   
  \=PULLU90\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU90\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30123\ );

  -- Alias \MST1\     
  \=PULLU91\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU91\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36116\ );

  -- Alias \MST2\     
  \=PULLU92\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU92\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36125\ );

  -- Alias \MST3\     
  \=PULLU93\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU93\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&36143\ );

  -- Alias \MSTPIT/\  
  \=PULLU94\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU94\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37244\ );

  -- Alias \MT02\     
  \=PULLU95\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU95\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37407\ );

  -- Alias \MT03\     
  \=PULLU96\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU96\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37411\ );

  -- Alias \MT04\     
  \=PULLU97\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU97\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37415\ );

  -- Alias \MT06\     
  \=PULLU98\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU98\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37427\ );

  -- Alias \MT07\     
  \=PULLU99\  : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU99\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37432\ );

  -- Alias \MT08\     
  \=PULLU100\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU100\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37437\ );

  -- Alias \MT09\     
  \=PULLU101\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU101\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37442\ );

  -- Alias \MT10\     
  \=PULLU102\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU102\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37447\ );

  -- Alias \MT11\     
  \=PULLU103\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU103\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37450\ );

  -- Alias \MTCSA/\   
  \=PULLU104\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU104\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30438\ );

  -- Alias \MWAG\     
  \=PULLU105\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU105\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33255\ );

  -- Alias \MWARNF/\  
  \=PULLU106\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU106\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&41223\ );

  -- Alias \MWBBEG\   
  \=PULLU107\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU107\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33315\ );

  -- Alias \MWBG\     
  \=PULLU108\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU108\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33135\ );

  -- Alias \MWEBG\    
  \=PULLU109\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU109\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33303\ );

  -- Alias \MWFBG\    
  \=PULLU110\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU110\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33311\ );

  -- Alias \MWG\      
  \=PULLU111\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU111\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33139\ );

  -- Alias \MWL07\    
  \=PULLU112\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU112\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52453\ );

  -- Alias \MWL08\    
  \=PULLU113\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU113\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52353\ );

  -- Alias \MWL09\    
  \=PULLU114\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU114\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53153\ );

  -- Alias \MWL10\    
  \=PULLU115\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU115\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53253\ );

  -- Alias \MWL11\    
  \=PULLU116\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU116\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53453\ );

  -- Alias \MWL12\    
  \=PULLU117\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU117\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&53353\ );

  -- Alias \MWL13\    
  \=PULLU118\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU118\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54153\ );

  -- Alias \MWL14\    
  \=PULLU119\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU119\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54253\ );

  -- Alias \MWL15\    
  \=PULLU120\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU120\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54453\ );

  -- Alias \MWL16\    
  \=PULLU121\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU121\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&54353\ );

  -- Alias \MWLG\     
  \=PULLU122\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU122\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33218\ );

  -- Alias \MWQG\     
  \=PULLU123\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU123\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33251\ );

  -- Alias \MWYG\     
  \=PULLU124\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU124\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33115\ );

  -- Alias \MWZG\     
  \=PULLU125\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU125\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33207\ );

  -- Alias \OUTCOM\   
  \=PULLU126\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU126\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&49339\ );

  -- Alias \Q2A\      
  \=PULLU127\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU127\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&37138\ );

  -- Alias \RESETA\   
  \=PULLU128\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU128\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42133\ );

  -- Alias \RESETB\   
  \=PULLU129\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU129\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42134\ );

  -- Alias \RESETC\   
  \=PULLU130\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU130\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42139\ );

  -- Alias \RESETD\   
  \=PULLU131\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU131\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42140\ );

  -- Alias \ROPER\    
  \=PULLU132\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU132\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52462\ );

  -- Alias \ROPES\    
  \=PULLU133\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU133\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52463\ );

  -- Alias \ROPET\    
  \=PULLU134\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU134\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&52363\ );

  -- Alias \RSTKX/\   
  \=PULLU135\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU135\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40224\ );

  -- Alias \RSTKY/\   
  \=PULLU136\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU136\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&40225\ );

  -- Alias \SBYREL/\  
  \=PULLU137\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU137\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42457\ );

  -- Alias \SCAS10\   
  \=PULLU138\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU138\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&30059\ );

  -- Alias \SCAS17\   
  \=PULLU139\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU139\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&32258\ );

  -- Alias \SETAB\    
  \=PULLU140\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU140\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42118\ );

  -- Alias \SETCD\    
  \=PULLU141\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU141\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42119\ );

  -- Alias \SETEK\    
  \=PULLU142\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU142\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42230\ );

  -- Alias \STR14\    
  \=PULLU143\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU143\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35421\ );

  -- Alias \STR19\    
  \=PULLU144\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU144\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35412\ );

  -- Alias \STR210\   
  \=PULLU145\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU145\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35409\ );

  -- Alias \STR311\   
  \=PULLU146\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU146\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35406\ );

  -- Alias \STR412\   
  \=PULLU147\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU147\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35403\ );

  -- Alias \STR58\    
  \=PULLU148\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU148\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35436\ );

  -- Alias \STR912\   
  \=PULLU149\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU149\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&35457\ );

  -- Alias \XB0E\     
  \=PULLU151\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU151\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42306\ );

  -- Alias \XB1E\     
  \=PULLU152\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU152\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42311\ );

  -- Alias \XB2E\     
  \=PULLU153\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU153\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42316\ );

  -- Alias \XB3E\     
  \=PULLU154\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU154\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42321\ );

  -- Alias \XB4E\     
  \=PULLU155\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU155\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42326\ );

  -- Alias \XB5E\     
  \=PULLU156\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU156\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42331\ );

  -- Alias \XB6E\     
  \=PULLU157\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU157\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42336\ );

  -- Alias \XB7E\     
  \=PULLU158\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU158\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42341\ );

  -- Alias \XT0E\     
  \=PULLU159\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU159\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42404\ );

  -- Alias \XT1E\     
  \=PULLU160\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU160\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42408\ );

  -- Alias \XT2E\     
  \=PULLU161\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU161\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42412\ );

  -- Alias \XT3E\     
  \=PULLU162\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU162\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42416\ );

  -- Alias \XT4E\     
  \=PULLU163\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU163\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42420\ );

  -- Alias \XT5E\     
  \=PULLU164\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU164\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42424\ );

  -- Alias \XT6E\     
  \=PULLU165\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU165\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42428\ );

  -- Alias \XT7E\     
  \=PULLU166\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU166\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42432\ );

  -- Alias \YB0E\     
  \=PULLU167\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU167\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42345\ );

  -- Alias \YB1E\     
  \=PULLU168\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU168\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42348\ );

  -- Alias \YB2E\     
  \=PULLU169\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU169\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42351\ );

  -- Alias \YB3E\     
  \=PULLU170\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU170\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&42354\ );

  -- Alias \YT0E\     
  \=PULLU171\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU171\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33435\ );

  -- Alias \YT1E\     
  \=PULLU172\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU172\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33438\ );

  -- Alias \YT2E\     
  \=PULLU173\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU173\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33441\ );

  -- Alias \YT3E\     
  \=PULLU174\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU174\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33444\ );

  -- Alias \YT4E\     
  \=PULLU175\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU175\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33447\ );

  -- Alias \YT5E\     
  \=PULLU176\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU176\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33450\ );

  -- Alias \YT6E\     
  \=PULLU177\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU177\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33453\ );

  -- Alias \YT7E\     
  \=PULLU178\ : LUT4_L generic map( INIT=>X"0001" ) port map(
                  LO =>  \PULLU178\,
                  I0 =>  \DERLO\,
                  I1 =>  '0',
                  I2 =>  '0',
                  I3 => \&33456\ );

  -- **************************************
  -- ***                                ***
  -- ***  Real gate alias assignments.  ***
  -- ***                                ***
  -- **************************************

  \CHAT05\    <= \38101\    ; -- A1 /1 - SCALER.
  \F10A\      <= \38102\    ; -- A1 /1 - SCALER.
  \FS10\      <= \38106\    ; -- A1 /1 - SCALER.
  \F10B\      <= \38107\    ; -- A1 /1 - SCALER.
  \CHAT06\    <= \38111\    ; -- A1 /1 - SCALER.
  \F11A\      <= \38112\    ; -- A1 /1 - SCALER.
  \FS11\      <= \38116\    ; -- A1 /1 - SCALER.
  \F11B\      <= \38117\    ; -- A1 /1 - SCALER.
  \CHAT07\    <= \38121\    ; -- A1 /1 - SCALER.
  \F12A\      <= \38122\    ; -- A1 /1 - SCALER.
  \FS12\      <= \38126\    ; -- A1 /1 - SCALER.
  \F12B\      <= \38127\    ; -- A1 /1 - SCALER.
  \CHAT08\    <= \38131\    ; -- A1 /1 - SCALER.
  \F13A\      <= \38132\    ; -- A1 /1 - SCALER.
  \FS13\      <= \38136\    ; -- A1 /1 - SCALER.
  \F13B\      <= \38137\    ; -- A1 /1 - SCALER.
  \CHAT09\    <= \38141\    ; -- A1 /1 - SCALER.
  \F14A\      <= \38142\    ; -- A1 /1 - SCALER.
  \FS14\      <= \38146\    ; -- A1 /1 - SCALER.
  \F14B\      <= \38147\    ; -- A1 /1 - SCALER.
  \CHAT10\    <= \38151\    ; -- A1 /1 - SCALER.
  \F15A\      <= \38152\    ; -- A1 /1 - SCALER.
  \FS15\      <= \38156\    ; -- A1 /1 - SCALER.
  \F15B\      <= \38157\    ; -- A1 /1 - SCALER.
  \CHAT11\    <= \38161\    ; -- A1 /1 - SCALER.
  \F16A\      <= \38162\    ; -- A1 /1 - SCALER.
  \FS16\      <= \38166\    ; -- A1 /1 - SCALER.
  \F16B\      <= \38167\    ; -- A1 /1 - SCALER.
  \CHAT12\    <= \38171\    ; -- A1 /1 - SCALER.
  \F17A\      <= \38172\    ; -- A1 /1 - SCALER.
  \FS17\      <= \38176\    ; -- A1 /1 - SCALER.
  \F17B\      <= \38177\    ; -- A1 /1 - SCALER.
  \FS06/\     <= \38190\    ; -- A1 /1 - SCALER.
  \FS07/\     <= \38191\    ; -- A1 /1 - SCALER.
  \FS02A\     <= \38201\    ; -- A1 /1 - SCALER.
  \F02A\      <= \38202\    ; -- A1 /1 - SCALER.
  \FS02\      <= \38206\    ; -- A1 /1 - SCALER.
  \F02B\      <= \38207\    ; -- A1 /1 - SCALER.
  \FS03A\     <= \38211\    ; -- A1 /1 - SCALER.
  \F03A\      <= \38212\    ; -- A1 /1 - SCALER.
  \FS03\      <= \38216\    ; -- A1 /1 - SCALER.
  \F03B\      <= \38217\    ; -- A1 /1 - SCALER.
  \FS04A\     <= \38221\    ; -- A1 /1 - SCALER.
  \F04A\      <= \38222\    ; -- A1 /1 - SCALER.
  \FS04\      <= \38226\    ; -- A1 /1 - SCALER.
  \F04B\      <= \38227\    ; -- A1 /1 - SCALER.
  \FS05A\     <= \38231\    ; -- A1 /1 - SCALER.
  \F05A\      <= \38232\    ; -- A1 /1 - SCALER.
  \FS05\      <= \38236\    ; -- A1 /1 - SCALER.
  \F05B\      <= \38237\    ; -- A1 /1 - SCALER.
  \CHAT01\    <= \38241\    ; -- A1 /1 - SCALER.
  \F06A\      <= \38242\    ; -- A1 /1 - SCALER.
  \FS06\      <= \38246\    ; -- A1 /1 - SCALER.
  \F06B\      <= \38247\    ; -- A1 /1 - SCALER.
  \CHAT02\    <= \38251\    ; -- A1 /1 - SCALER.
  \F07A\      <= \38252\    ; -- A1 /1 - SCALER.
  \FS07\      <= \38256\    ; -- A1 /1 - SCALER.
  \F07B\      <= \38257\    ; -- A1 /1 - SCALER.
  \CHAT03\    <= \38261\    ; -- A1 /1 - SCALER.
  \F08A\      <= \38262\    ; -- A1 /1 - SCALER.
  \FS08\      <= \38266\    ; -- A1 /1 - SCALER.
  \F08B\      <= \38267\    ; -- A1 /1 - SCALER.
  \CHAT04\    <= \38271\    ; -- A1 /1 - SCALER.
  \F09A\      <= \38272\    ; -- A1 /1 - SCALER.
  \FS09\      <= \38276\    ; -- A1 /1 - SCALER.
  \F09B\      <= \38277\    ; -- A1 /1 - SCALER.
  \FS08/\     <= \38290\    ; -- A1 /1 - SCALER.
  \FS07A\     <= \38291\    ; -- A1 /1 - SCALER.
  \CHAT13\    <= \38301\    ; -- A1 /2 - SCALER.
  \F18A\      <= \38302\    ; -- A1 /2 - SCALER.
  \FS18\      <= \38306\    ; -- A1 /2 - SCALER.
  \F18B\      <= \38307\    ; -- A1 /2 - SCALER.
  \CHAT14\    <= \38311\    ; -- A1 /2 - SCALER.
  \F19A\      <= \38312\    ; -- A1 /2 - SCALER.
  \FS19\      <= \38316\    ; -- A1 /2 - SCALER.
  \F19B\      <= \38317\    ; -- A1 /2 - SCALER.
  \CHBT01\    <= \38321\    ; -- A1 /2 - SCALER.
  \F20A\      <= \38322\    ; -- A1 /2 - SCALER.
  \FS20\      <= \38326\    ; -- A1 /2 - SCALER.
  \F20B\      <= \38327\    ; -- A1 /2 - SCALER.
  \CHBT02\    <= \38331\    ; -- A1 /2 - SCALER.
  \F21A\      <= \38332\    ; -- A1 /2 - SCALER.
  \FS21\      <= \38336\    ; -- A1 /2 - SCALER.
  \F21B\      <= \38337\    ; -- A1 /2 - SCALER.
  \CHBT03\    <= \38341\    ; -- A1 /2 - SCALER.
  \F22A\      <= \38342\    ; -- A1 /2 - SCALER.
  \FS22\      <= \38346\    ; -- A1 /2 - SCALER.
  \F22B\      <= \38347\    ; -- A1 /2 - SCALER.
  \CHBT04\    <= \38351\    ; -- A1 /2 - SCALER.
  \F23A\      <= \38352\    ; -- A1 /2 - SCALER.
  \FS23\      <= \38356\    ; -- A1 /2 - SCALER.
  \F23B\      <= \38357\    ; -- A1 /2 - SCALER.
  \CHBT05\    <= \38361\    ; -- A1 /2 - SCALER.
  \F24A\      <= \38362\    ; -- A1 /2 - SCALER.
  \FS24\      <= \38366\    ; -- A1 /2 - SCALER.
  \F24B\      <= \38367\    ; -- A1 /2 - SCALER.
  \CHBT06\    <= \38371\    ; -- A1 /2 - SCALER.
  \F25A\      <= \38372\    ; -- A1 /2 - SCALER.
  \FS25\      <= \38376\    ; -- A1 /2 - SCALER.
  \F25B\      <= \38377\    ; -- A1 /2 - SCALER.
  \F18AX\     <= \38390\    ; -- A1 /2 - SCALER.
  \F07A/\     <= \38391\    ; -- A1 /2 - SCALER.
  \CHBT07\    <= \38401\    ; -- A1 /2 - SCALER.
  \F26A\      <= \38402\    ; -- A1 /2 - SCALER.
  \FS26\      <= \38406\    ; -- A1 /2 - SCALER.
  \F26B\      <= \38407\    ; -- A1 /2 - SCALER.
  \CHBT08\    <= \38411\    ; -- A1 /2 - SCALER.
  \F27A\      <= \38412\    ; -- A1 /2 - SCALER.
  \FS27\      <= \38416\    ; -- A1 /2 - SCALER.
  \F27B\      <= \38417\    ; -- A1 /2 - SCALER.
  \CHBT09\    <= \38421\    ; -- A1 /2 - SCALER.
  \F28A\      <= \38422\    ; -- A1 /2 - SCALER.
  \FS28\      <= \38426\    ; -- A1 /2 - SCALER.
  \F28B\      <= \38427\    ; -- A1 /2 - SCALER.
  \CHBT10\    <= \38431\    ; -- A1 /2 - SCALER.
  \F29A\      <= \38432\    ; -- A1 /2 - SCALER.
  \FS29\      <= \38436\    ; -- A1 /2 - SCALER.
  \F29B\      <= \38437\    ; -- A1 /2 - SCALER.
  \CHBT11\    <= \38441\    ; -- A1 /2 - SCALER.
  \F30A\      <= \38442\    ; -- A1 /2 - SCALER.
  \FS30\      <= \38446\    ; -- A1 /2 - SCALER.
  \F30B\      <= \38447\    ; -- A1 /2 - SCALER.
  \CHBT12\    <= \38451\    ; -- A1 /2 - SCALER.
  \F31A\      <= \38452\    ; -- A1 /2 - SCALER.
  \FS31\      <= \38456\    ; -- A1 /2 - SCALER.
  \F31B\      <= \38457\    ; -- A1 /2 - SCALER.
  \CHBT13\    <= \38461\    ; -- A1 /2 - SCALER.
  \F32A\      <= \38462\    ; -- A1 /2 - SCALER.
  \FS32\      <= \38466\    ; -- A1 /2 - SCALER.
  \F32B\      <= \38467\    ; -- A1 /2 - SCALER.
  \CHBT14\    <= \38471\    ; -- A1 /2 - SCALER.
  \F33A\      <= \38472\    ; -- A1 /2 - SCALER.
  \FS33\      <= \38476\    ; -- A1 /2 - SCALER.
  \F33B\      <= \38477\    ; -- A1 /2 - SCALER.
  \F18A/\     <= \38490\    ; -- A1 /2 - SCALER.
  \F03B/\     <= \38491\    ; -- A1 /2 - SCALER.
  \PHS2\      <= \37104\    ; -- A2 /1 - TIMER.
  \PHS4\      <= \37108\    ; -- A2 /1 - TIMER.
  \PHS4/\     <= \37109\    ; -- A2 /1 - TIMER.
  \RINGA/\    <= \37115\    ; -- A2 /1 - TIMER.
  \RINGB/\    <= \37119\    ; -- A2 /1 - TIMER.
  \ODDSET/\   <= \37122\    ; -- A2 /1 - TIMER.
  \EVNSET\    <= \37125\    ; -- A2 /1 - TIMER.
  \EVNSET/\   <= \37126\    ; -- A2 /1 - TIMER.
  \RT\        <= \37129\    ; -- A2 /1 - TIMER.
  \WT\        <= \37130\    ; -- A2 /1 - TIMER.
  \WT/\       <= \37131\    ; -- A2 /1 - TIMER.
  \TT/\       <= \37135\    ; -- A2 /1 - TIMER.
  \CLK\       <= \37137\    ; -- A2 /1 - TIMER.
  \CT\        <= \37140\    ; -- A2 /1 - TIMER.
  \CT/\       <= \37142\    ; -- A2 /1 - TIMER.
  \OVFSTB/\   <= \37151\    ; -- A2 /1 - TIMER.
  \PHS2/\     <= \37155\    ; -- A2 /1 - TIMER.
  \P01\       <= \37203\    ; -- A2 /2 - TIMER.
  \P01/\      <= \37204\    ; -- A2 /2 - TIMER.
  \P02\       <= \37207\    ; -- A2 /2 - TIMER.
  \P02/\      <= \37208\    ; -- A2 /2 - TIMER.
  \P03\       <= \37211\    ; -- A2 /2 - TIMER.
  \P03/\      <= \37212\    ; -- A2 /2 - TIMER.
  \P04\       <= \37215\    ; -- A2 /2 - TIMER.
  \P04/\      <= \37216\    ; -- A2 /2 - TIMER.
  \P05\       <= \37219\    ; -- A2 /2 - TIMER.
  \P05/\      <= \37220\    ; -- A2 /2 - TIMER.
  \F01D\      <= \37221\    ; -- A2 /2 - TIMER.
  \F01B\      <= \37222\    ; -- A2 /2 - TIMER.
  \F01A\      <= \37223\    ; -- A2 /2 - TIMER.
  \F01C\      <= \37224\    ; -- A2 /2 - TIMER.
  \FS01/\     <= \37225\    ; -- A2 /2 - TIMER.
  \FS01\      <= \37226\    ; -- A2 /2 - TIMER.
  \GOSET/\    <= \37228\    ; -- A2 /2 - TIMER.
  \STOPA\     <= \37234\    ; -- A2 /2 - TIMER.
  \GOJAM/\    <= \37240\    ; -- A2 /2 - TIMER.
  \STOP/\     <= \37242\    ; -- A2 /2 - TIMER.
  \STOP\      <= \37243\    ; -- A2 /2 - TIMER.
  \GOJAM\     <= \37245\    ; -- A2 /2 - TIMER.
  \SB0\       <= \37255\    ; -- A2 /2 - TIMER.
  \SB1\       <= \37256\    ; -- A2 /2 - TIMER.
  \SB2\       <= \37257\    ; -- A2 /2 - TIMER.
  \SB4\       <= \37258\    ; -- A2 /2 - TIMER.
  \EDSET\     <= \37259\    ; -- A2 /2 - TIMER.
  \T12\       <= \37301\    ; -- A2 /3 - TIMER.
  \T12DC/\    <= \37302\    ; -- A2 /3 - TIMER.
  \T01DC/\    <= \37305\    ; -- A2 /3 - TIMER.
  \T01\       <= \37307\    ; -- A2 /3 - TIMER.
  \T02DC/\    <= \37309\    ; -- A2 /3 - TIMER.
  \T02\       <= \37311\    ; -- A2 /3 - TIMER.
  \T03DC/\    <= \37313\    ; -- A2 /3 - TIMER.
  \T03\       <= \37315\    ; -- A2 /3 - TIMER.
  \T04\       <= \37319\    ; -- A2 /3 - TIMER.
  \T05\       <= \37323\    ; -- A2 /3 - TIMER.
  \T06DC/\    <= \37326\    ; -- A2 /3 - TIMER.
  \T06\       <= \37328\    ; -- A2 /3 - TIMER.
  \T07DC/\    <= \37330\    ; -- A2 /3 - TIMER.
  \T07\       <= \37332\    ; -- A2 /3 - TIMER.
  \T08DC/\    <= \37334\    ; -- A2 /3 - TIMER.
  \T08\       <= \37336\    ; -- A2 /3 - TIMER.
  \T09DC/\    <= \37338\    ; -- A2 /3 - TIMER.
  \T09\       <= \37340\    ; -- A2 /3 - TIMER.
  \T10DC/\    <= \37342\    ; -- A2 /3 - TIMER.
  \T10\       <= \37344\    ; -- A2 /3 - TIMER.
  \T11\       <= \37349\    ; -- A2 /3 - TIMER.
  \RT/\       <= \37350\    ; -- A2 /3 - TIMER.
  \OVF\       <= \37353\    ; -- A2 /3 - TIMER.
  \UNF\       <= \37354\    ; -- A2 /3 - TIMER.
  \T12SET\    <= \37355\    ; -- A2 /3 - TIMER.
  \T01/\      <= \37401\    ; -- A2 /3 - TIMER.
  \T02/\      <= \37405\    ; -- A2 /3 - TIMER.
  \T03/\      <= \37408\    ; -- A2 /3 - TIMER.
  \T04/\      <= \37412\    ; -- A2 /3 - TIMER.
  \T05/\      <= \37416\    ; -- A2 /3 - TIMER.
  \T06/\      <= \37423\    ; -- A2 /3 - TIMER.
  \T07/\      <= \37428\    ; -- A2 /3 - TIMER.
  \T08/\      <= \37433\    ; -- A2 /3 - TIMER.
  \T09/\      <= \37438\    ; -- A2 /3 - TIMER.
  \T10/\      <= \37443\    ; -- A2 /3 - TIMER.
  \T11/\      <= \37448\    ; -- A2 /3 - TIMER.
  \T12/\      <= \37451\    ; -- A2 /3 - TIMER.
  \OVF/\      <= \37455\    ; -- A2 /3 - TIMER.
  \UNF/\      <= \37456\    ; -- A2 /3 - TIMER.
  \NISQL/\    <= \30004\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \CSQG\      <= \30007\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \RBSQ\      <= \30009\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \WSQG/\     <= \30011\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR16\     <= \30017\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR14\     <= \30019\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR13\     <= \30021\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ5\       <= \30039\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ0/\      <= \30045\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ1/\      <= \30048\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ2/\      <= \30049\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ3/\      <= \30053\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ4/\      <= \30054\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ6/\      <= \30055\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ7/\      <= \30056\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \CON1\      <= \30057\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \CON2\      <= \30058\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \INKBT1\    <= \30061\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \INHINT\    <= \30104\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \IIP/\      <= \30105\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \IIP\       <= \30106\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \STRTFC\    <= \30107\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \FUTEXT\    <= \30110\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \RPTSET\    <= \30117\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQEXT/\    <= \30124\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \RPTFRC\    <= \30127\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR12\     <= \30133\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR11\     <= \30135\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \QC0\       <= \30141\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \QC0/\      <= \30145\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \QC1/\      <= \30148\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \QC2/\      <= \30151\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \QC3/\      <= \30152\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR10\     <= \30154\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR10/\    <= \30156\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQR12/\    <= \30157\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQEXT\     <= \30160\    ; -- A3 /1 - SQ REGISTER AND DECODING.
  \SQ5QC0/\   <= \30303\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC1\       <= \30305\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC2\       <= \30306\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC2/\      <= \30309\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \SQ5/\      <= \30310\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC11\      <= \30313\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \EXST1/\    <= \30316\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC6\       <= \30317\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC7\       <= \30318\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TC0\       <= \30319\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TCF0\      <= \30320\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NEXST0\    <= \30321\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TC0/\      <= \30322\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC3/\      <= \30323\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NEXST0/\   <= \30324\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC3\       <= \30326\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DCS0\      <= \30327\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DCA0\      <= \30328\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC4/\      <= \30329\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC4\       <= \30330\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC13/\     <= \30331\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC13\      <= \30333\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC5\       <= \30338\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC5/\      <= \30339\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC9/\      <= \30340\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \LXCH0\     <= \30341\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \QXCH0\     <= \30342\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \QXCH0/\    <= \30343\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC9\       <= \30345\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC8/\      <= \30346\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TS0\       <= \30348\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \EXST0/\    <= \30349\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TS0/\      <= \30350\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DXCH0\     <= \30352\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DAS0\      <= \30354\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC10/\     <= \30356\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC10\      <= \30357\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DAS0/\     <= \30401\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \BZF0\      <= \30403\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \BZF0/\     <= \30404\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \BMF0\      <= \30405\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \BMF0/\     <= \30406\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC16/\     <= \30409\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC15/\     <= \30410\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC16\      <= \30411\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC17\      <= \30412\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC15\      <= \30413\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \CCS0\      <= \30415\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \CCS0/\     <= \30416\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DAS1/\     <= \30419\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DAS1\      <= \30421\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC12/\     <= \30422\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC12\      <= \30423\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \ADS0\      <= \30424\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \INCR0\     <= \30425\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MSU0\      <= \30426\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MSU0/\     <= \30427\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \AUG0\      <= \30428\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \AUG0/\     <= \30429\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DIM0\      <= \30430\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DIM0/\     <= \30431\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP3\       <= \30432\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP3/\      <= \30433\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP1\       <= \30435\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP1/\      <= \30436\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP0\       <= \30437\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MP0/\      <= \30439\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TCSAJ3\    <= \30441\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \TCSAJ3/\   <= \30442\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \RSM3\      <= \30443\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \RSM3/\     <= \30444\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \SU0\       <= \30445\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MASK0\     <= \30446\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \MASK0/\    <= \30447\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \AD0\       <= \30448\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NDX0\      <= \30449\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NDX0/\     <= \30450\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NDXX1\     <= \30451\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \NDXX1/\    <= \30452\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \GOJ1\      <= \30453\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \GOJ1/\     <= \30454\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \IC14\      <= \30456\    ; -- A3 /2 - SQ REGISTER AND DECODING.
  \DIVSTG\    <= \36101\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \T12USE/\   <= \36102\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST0/\      <= \36106\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \MP3A\      <= \36108\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST1/\      <= \36117\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \STG1\      <= \36120\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST1D\      <= \36121\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST1376/\   <= \36126\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV1376\    <= \36127\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV1376/\   <= \36128\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \STG2\      <= \36137\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \STD2\      <= \36138\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST3/\      <= \36141\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST4/\      <= \36145\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \STG3\      <= \36151\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST376\     <= \36153\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \ST376/\    <= \36154\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV3764\    <= \36157\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DIV/\      <= \36202\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV0\       <= \36204\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV0/\      <= \36205\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV376\     <= \36206\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV376/\    <= \36207\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV4\       <= \36208\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV1\       <= \36209\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV1/\      <= \36210\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \SGUM\      <= \36214\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \BR1\       <= \36220\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \BR1/\      <= \36226\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \BR2\       <= \36238\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \BR2/\      <= \36246\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \TRSM/\     <= \36263\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DVST/\     <= \36264\    ; -- A4 /1 - STAGE BRANCH DECODING.
  \DV4/\      <= \36301\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \READ0\     <= \36305\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \READ0/\    <= \36306\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WRITE0\    <= \36308\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WRITE0/\   <= \36309\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RAND0\     <= \36310\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WAND0\     <= \36312\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \INOUT/\    <= \36313\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \INOUT\     <= \36314\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \ROR0\      <= \36315\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WOR0\      <= \36316\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WOR0/\     <= \36317\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RXOR0\     <= \36318\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RXOR0/\    <= \36319\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RUPT0\     <= \36320\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RUPT0/\    <= \36321\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \8PP4\      <= \36322\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RUPT1\     <= \36323\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RUPT1/\    <= \36324\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \PRINC\     <= \36327\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RRPA\      <= \36331\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \3XP7\      <= \36332\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \9XP1\      <= \36336\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \5XP28\     <= \36341\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \5XP11\     <= \36344\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \WCH/\      <= \36350\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \2XP3\      <= \36352\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \R15\       <= \36402\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RB2\       <= \36403\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \1XP10\     <= \36404\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \2PP1\      <= \36405\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \2XP5\      <= \36408\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \RSC/\      <= \36410\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \3XP2\      <= \36416\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR1B2\     <= \36417\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR1B2/\    <= \36418\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR12B\     <= \36419\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR12B/\    <= \36420\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BRDIF/\    <= \36421\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR1B2B\    <= \36422\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \BR1B2B/\   <= \36423\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \4XP5\      <= \36429\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \8XP5\      <= \36432\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \4XP11\     <= \36433\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \8XP6\      <= \36434\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \B15X\      <= \36443\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \5XP4\      <= \36445\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \6XP5\      <= \36447\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \KRPT\      <= \36448\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \TL15\      <= \36449\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \MP0T10\    <= \36450\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \TSGN2\     <= \36455\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \7XP19\     <= \36457\    ; -- A4 /2 - STAGE BRANCH DECODING.
  \NISQ/\     <= \39113\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \DVST\      <= \39115\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \2XP7\      <= \39117\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \3XP6\      <= \39122\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \TPZG/\     <= \39126\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \PARTC\     <= \39132\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \5XP12\     <= \39136\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \TSGN/\     <= \39137\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \7XP9\      <= \39147\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \7XP4\      <= \39150\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \PTWOX\     <= \39151\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \TSUDO/\    <= \39205\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \RAD\       <= \39207\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \8XP15\     <= \39210\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \8XP3\      <= \39212\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \RSTRT\     <= \39219\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \8XP12\     <= \39220\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \9XP5\      <= \39224\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \10XP6\     <= \39229\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \10XP1\     <= \39231\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \10XP7\     <= \39236\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \10XP8\     <= \39238\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \11XP2\     <= \39240\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \GNHNC\     <= \39249\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \PINC/\     <= \39255\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \PINC\      <= \39256\    ; -- A5 /1 - CROSS POINT GENERATOR NQI.
  \RL10BB\    <= \39304\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \R6\        <= \39306\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \2XP8\      <= \39308\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \RSCT\      <= \39309\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \RQ\        <= \39314\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \RL/\       <= \39321\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \RA/\       <= \39322\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \TRSM\      <= \39323\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \WY12/\     <= \39331\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \5XP9\      <= \39332\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \WY/\       <= \39333\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \5XP13\     <= \39337\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \5XP15\     <= \39339\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \5XP21\     <= \39340\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \SCAD\      <= \39346\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \SCAD/\     <= \39347\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \NDR100/\   <= \39350\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \OCTAD2\    <= \39352\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \OCTAD3\    <= \39353\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \OCTAD4\    <= \39354\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \OCTAD5\    <= \39355\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \OCTAD6\    <= \39356\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \DV1B1B\    <= \39402\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \5XP19\     <= \39407\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \6XP8\      <= \39419\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \6XP7\      <= \39420\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \6XP2\      <= \39421\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \U2BBK\     <= \39426\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \RSTSTG\    <= \39431\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \TMZ/\      <= \39440\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \10XP10\    <= \39442\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \DV4B1B\    <= \39446\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \11XP6\     <= \39450\    ; -- A5 /2 - CROSS POINT GENERATOR NQI.
  \DVXP1\     <= \40106\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \A2X/\      <= \40107\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \L2GD/\     <= \40108\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RB/\       <= \40109\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WYD/\      <= \40110\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \ZIP\       <= \40117\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \ZIPCI\     <= \40130\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RC/\       <= \40131\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RCH/\      <= \40132\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \TSGU/\     <= \40139\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WL/\       <= \40140\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RG/\       <= \40146\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \ZAP/\      <= \40152\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \ZAP\       <= \40154\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WB/\       <= \40155\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RU/\       <= \40156\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WZ/\       <= \40158\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \MCRO/\     <= \40160\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \RB1F\      <= \40201\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \CLXC\      <= \40202\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WQ/\       <= \40206\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \TOV/\      <= \40207\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WSC/\      <= \40208\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \WG/\       <= \40209\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \MONEX\     <= \40210\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \TWOX\      <= \40214\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \BXVX\      <= \40216\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \PIFL/\     <= \40220\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \CGMC\      <= \40241\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \TIMR\      <= \40251\    ; -- A6 /1 - CROSS POINT GENERATOR II.
  \6XP10\     <= \40305\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \MONEX/\    <= \40311\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \POUT\      <= \40320\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \MOUT\      <= \40321\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \ZOUT\      <= \40322\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \7XP7\      <= \40327\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \7XP14\     <= \40331\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \WOVR\      <= \40341\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \8XP4\      <= \40349\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \8XP10\     <= \40350\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \RD_BANK\   <= \40357\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \EXT\       <= \40402\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \10XP9\     <= \40403\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \WA/\       <= \40414\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \RUS/\      <= \40419\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \RZ/\       <= \40420\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \ST1\       <= \40423\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \ST2/\      <= \40424\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \ST2\       <= \40425\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \NEAC\      <= \40427\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \WS/\       <= \40430\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \CI/\       <= \40431\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \PONEX\     <= \40434\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \R1C/\      <= \40435\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \RB1/\      <= \40436\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \PSEUDO\    <= \40440\    ; -- A6 /2 - CROSS POINT GENERATOR II.
  \WALSG/\    <= \33101\    ; -- A7 /1 - SERVICE GATES.
  \WALSG\     <= \33102\    ; -- A7 /1 - SERVICE GATES.
  \WYLOG/\    <= \33109\    ; -- A7 /1 - SERVICE GATES.
  \WYHIG/\    <= \33112\    ; -- A7 /1 - SERVICE GATES.
  \CUG\       <= \33116\    ; -- A7 /1 - SERVICE GATES.
  \WYDG/\     <= \33126\    ; -- A7 /1 - SERVICE GATES.
  \WYDLOG/\   <= \33129\    ; -- A7 /1 - SERVICE GATES.
  \WBG/\      <= \33131\    ; -- A7 /1 - SERVICE GATES.
  \CBG\       <= \33136\    ; -- A7 /1 - SERVICE GATES.
  \WGNORM\    <= \33140\    ; -- A7 /1 - SERVICE GATES.
  \WG1G/\     <= \33141\    ; -- A7 /1 - SERVICE GATES.
  \WG2G/\     <= \33145\    ; -- A7 /1 - SERVICE GATES.
  \WG4G/\     <= \33146\    ; -- A7 /1 - SERVICE GATES.
  \WG5G/\     <= \33150\    ; -- A7 /1 - SERVICE GATES.
  \WG3G/\     <= \33152\    ; -- A7 /1 - SERVICE GATES.
  \WEDOPG/\   <= \33156\    ; -- A7 /1 - SERVICE GATES.
  \PIPSAM\    <= \33160\    ; -- A7 /1 - SERVICE GATES.
  \WZG/\      <= \33202\    ; -- A7 /1 - SERVICE GATES.
  \CZG\       <= \33208\    ; -- A7 /1 - SERVICE GATES.
  \WLG/\      <= \33214\    ; -- A7 /1 - SERVICE GATES.
  \CLG2G\     <= \33221\    ; -- A7 /1 - SERVICE GATES.
  \CLG1G\     <= \33224\    ; -- A7 /1 - SERVICE GATES.
  \WAG/\      <= \33229\    ; -- A7 /1 - SERVICE GATES.
  \CAG\       <= \33234\    ; -- A7 /1 - SERVICE GATES.
  \WSG/\      <= \33238\    ; -- A7 /1 - SERVICE GATES.
  \CSG\       <= \33242\    ; -- A7 /1 - SERVICE GATES.
  \WQG/\      <= \33247\    ; -- A7 /1 - SERVICE GATES.
  \CQG\       <= \33252\    ; -- A7 /1 - SERVICE GATES.
  \P04A\      <= \33257\    ; -- A7 /1 - SERVICE GATES.
  \WEBG/\     <= \33302\    ; -- A7 /2 - SERVICE GATES.
  \CEBG\      <= \33306\    ; -- A7 /2 - SERVICE GATES.
  \WFBG/\     <= \33308\    ; -- A7 /2 - SERVICE GATES.
  \CFBG\      <= \33310\    ; -- A7 /2 - SERVICE GATES.
  \WBBEG/\    <= \33313\    ; -- A7 /2 - SERVICE GATES.
  \RGG1\      <= \33316\    ; -- A7 /2 - SERVICE GATES.
  \RGG/\      <= \33317\    ; -- A7 /2 - SERVICE GATES.
  \RAG/\      <= \33323\    ; -- A7 /2 - SERVICE GATES.
  \REBG/\     <= \33328\    ; -- A7 /2 - SERVICE GATES.
  \RLG2\      <= \33329\    ; -- A7 /2 - SERVICE GATES.
  \RLG/\      <= \33330\    ; -- A7 /2 - SERVICE GATES.
  \RLG1\      <= \33331\    ; -- A7 /2 - SERVICE GATES.
  \RLG3\      <= \33333\    ; -- A7 /2 - SERVICE GATES.
  \RZG/\      <= \33338\    ; -- A7 /2 - SERVICE GATES.
  \RULOG/\    <= \33342\    ; -- A7 /2 - SERVICE GATES.
  \RUG/\      <= \33348\    ; -- A7 /2 - SERVICE GATES.
  \RUSG/\     <= \33349\    ; -- A7 /2 - SERVICE GATES.
  \RBHG/\     <= \33351\    ; -- A7 /2 - SERVICE GATES.
  \RBLG/\     <= \33353\    ; -- A7 /2 - SERVICE GATES.
  \CI01/\     <= \33356\    ; -- A7 /2 - SERVICE GATES.
  \RCG/\      <= \33402\    ; -- A7 /2 - SERVICE GATES.
  \RQG/\      <= \33406\    ; -- A7 /2 - SERVICE GATES.
  \RFBG/\     <= \33412\    ; -- A7 /2 - SERVICE GATES.
  \RBBEG/\    <= \33414\    ; -- A7 /2 - SERVICE GATES.
  \G2LSG\     <= \33415\    ; -- A7 /2 - SERVICE GATES.
  \G2LSG/\    <= \33416\    ; -- A7 /2 - SERVICE GATES.
  \L2GDG/\    <= \33420\    ; -- A7 /2 - SERVICE GATES.
  \A2XG/\     <= \33424\    ; -- A7 /2 - SERVICE GATES.
  \CGG\       <= \33430\    ; -- A7 /2 - SERVICE GATES.
  \YT0\       <= \33433\    ; -- A7 /2 - SERVICE GATES.
  \YT0/\      <= \33434\    ; -- A7 /2 - SERVICE GATES.
  \YT1\       <= \33436\    ; -- A7 /2 - SERVICE GATES.
  \YT1/\      <= \33437\    ; -- A7 /2 - SERVICE GATES.
  \YT2\       <= \33439\    ; -- A7 /2 - SERVICE GATES.
  \YT2/\      <= \33440\    ; -- A7 /2 - SERVICE GATES.
  \YT3\       <= \33442\    ; -- A7 /2 - SERVICE GATES.
  \YT3/\      <= \33443\    ; -- A7 /2 - SERVICE GATES.
  \YT4\       <= \33445\    ; -- A7 /2 - SERVICE GATES.
  \YT4/\      <= \33446\    ; -- A7 /2 - SERVICE GATES.
  \YT5\       <= \33448\    ; -- A7 /2 - SERVICE GATES.
  \YT5/\      <= \33449\    ; -- A7 /2 - SERVICE GATES.
  \YT6\       <= \33451\    ; -- A7 /2 - SERVICE GATES.
  \YT6/\      <= \33452\    ; -- A7 /2 - SERVICE GATES.
  \YT7\       <= \33454\    ; -- A7 /2 - SERVICE GATES.
  \YT7/\      <= \33455\    ; -- A7 /2 - SERVICE GATES.
  \CINORM\    <= \33457\    ; -- A7 /2 - SERVICE GATES.
  \CIFF\      <= \33459\    ; -- A7 /2 - SERVICE GATES.
  \RBBK\      <= \33460\    ; -- A7 /2 - SERVICE GATES.
  \CO04\      <= \51101\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \XUY01/\    <= \51110\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \SUMA01/\   <= \51112\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \CI02/\     <= \51114\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \SUMB01/\   <= \51115\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \A01/\      <= \51120\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \L01/\      <= \51126\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \Z01/\      <= \51135\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \G01/\      <= \51148\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \G01\       <= \51149\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \WL01\      <= \51152\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \WL01/\     <= \51154\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \RL01/\     <= \51157\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \CLEARA\    <= \51161\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \XUY02/\    <= \51210\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \SUMA02/\   <= \51212\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \CI03/\     <= \51214\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \SUMB02/\   <= \51215\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \A02/\      <= \51220\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \L02/\      <= \51226\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \Z02/\      <= \51235\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \G02/\      <= \51248\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \G02\       <= \51249\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \WL02\      <= \51252\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \WL02/\     <= \51254\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \RL02/\     <= \51257\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \S08A/\     <= \51261\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \S08A\      <= \51262\    ; -- A8 /1 - 4 BIT MODULE (1 OF 4).
  \XUY04/\    <= \51310\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \SUMA04/\   <= \51312\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CI05/\     <= \51314\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \SUMB04/\   <= \51315\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \A04/\      <= \51320\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \L04/\      <= \51326\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \Z04/\      <= \51335\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \G04/\      <= \51348\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \G04\       <= \51349\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \WL04\      <= \51352\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \WL04/\     <= \51354\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \RL04/\     <= \51357\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CLEARC\    <= \51361\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CLEARD\    <= \51362\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CO06\      <= \51401\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \XUY03/\    <= \51410\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \SUMA03/\   <= \51412\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CI04/\     <= \51414\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \SUMB03/\   <= \51415\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \A03/\      <= \51420\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \L03/\      <= \51426\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \Z03/\      <= \51435\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \G03/\      <= \51448\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \G03\       <= \51449\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \WL03\      <= \51452\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \WL03/\     <= \51454\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \RL03/\     <= \51457\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CLEARB\    <= \51461\    ; -- A8 /2 - 4 BIT MODULE (1 OF 4).
  \CO08\      <= \52101\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \XUY05/\    <= \52110\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \SUMA05/\   <= \52112\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \CI06/\     <= \52114\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \SUMB05/\   <= \52115\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \A05/\      <= \52120\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \L05/\      <= \52126\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \Z05/\      <= \52135\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \G05/\      <= \52148\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \G05\       <= \52149\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \WL05\      <= \52152\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \WL05/\     <= \52154\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \RL05/\     <= \52157\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \XUY06/\    <= \52210\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \SUMA06/\   <= \52212\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \CI07/\     <= \52214\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \SUMB06/\   <= \52215\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \A06/\      <= \52220\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \L06/\      <= \52226\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \Z06/\      <= \52235\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \G06/\      <= \52248\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \G06\       <= \52249\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \WL06\      <= \52252\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \WL06/\     <= \52254\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \RL06/\     <= \52257\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \PIPSAM/\   <= \52261\    ; -- A9 /1 - 4 BIT MODULE (2 OF 4).
  \XUY08/\    <= \52310\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \SUMA08/\   <= \52312\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \CI09/\     <= \52314\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \SUMB08/\   <= \52315\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \A08/\      <= \52320\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \L08/\      <= \52326\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \Z08/\      <= \52335\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \G08/\      <= \52348\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \G08\       <= \52349\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \WL08\      <= \52352\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \WL08/\     <= \52354\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \RL08/\     <= \52357\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \PIPGX-\    <= \52361\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \PIPGY+\    <= \52362\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \CO10\      <= \52401\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \XUY07/\    <= \52410\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \SUMA07/\   <= \52412\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \CI08/\     <= \52414\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \SUMB07/\   <= \52415\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \A07/\      <= \52420\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \L07/\      <= \52426\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \Z07/\      <= \52435\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \G07/\      <= \52448\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \G07\       <= \52449\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \WL07\      <= \52452\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \WL07/\     <= \52454\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \RL07/\     <= \52457\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \PIPGX+\    <= \52461\    ; -- A9 /2 - 4 BIT MODULE (2 OF 4).
  \CO12\      <= \53101\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \XUY09/\    <= \53110\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \SUMA09/\   <= \53112\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \CI10/\     <= \53114\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \SUMB09/\   <= \53115\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \A09/\      <= \53120\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \L09/\      <= \53126\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \Z09/\      <= \53135\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \G09/\      <= \53148\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \G09\       <= \53149\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \WL09\      <= \53152\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \WL09/\     <= \53154\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \RL09/\     <= \53157\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \PIPGY-\    <= \53161\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \XUY10/\    <= \53210\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \SUMA10/\   <= \53212\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \CI11/\     <= \53214\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \SUMB10/\   <= \53215\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \A10/\      <= \53220\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \L10/\      <= \53226\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \Z10/\      <= \53235\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \G10/\      <= \53248\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \G10\       <= \53249\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \WL10\      <= \53252\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \WL10/\     <= \53254\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \RL10/\     <= \53257\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \PIPGZ+\    <= \53261\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \PIPGZ-\    <= \53262\    ; -- A10/1 - 4 BIT MODULE (3 OF 4).
  \XUY12/\    <= \53310\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \SUMA12/\   <= \53312\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \CI13/\     <= \53314\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \SUMB12/\   <= \53315\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \A12/\      <= \53320\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \L12/\      <= \53326\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \Z12/\      <= \53335\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \G12/\      <= \53348\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \G12\       <= \53349\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \WL12\      <= \53352\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \WL12/\     <= \53354\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \RL12/\     <= \53357\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \PIPAX-/\   <= \53361\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \PIPAY+/\   <= \53362\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \CO14\      <= \53401\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \XUY11/\    <= \53410\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \SUMA11/\   <= \53412\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \CI12/\     <= \53414\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \SUMB11/\   <= \53415\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \A11/\      <= \53420\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \L11/\      <= \53426\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \Z11/\      <= \53435\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \G11/\      <= \53448\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \G11\       <= \53449\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \WL11\      <= \53452\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \WL11/\     <= \53454\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \RL11/\     <= \53457\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \PIPAX+/\   <= \53461\    ; -- A10/2 - 4 BIT MODULE (3 OF 4).
  \CO16\      <= \54101\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \XUY13/\    <= \54110\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \SUMA13/\   <= \54112\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \CI14/\     <= \54114\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \SUMB13/\   <= \54115\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \A13/\      <= \54120\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \L13/\      <= \54126\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \Z13/\      <= \54135\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \G13/\      <= \54148\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \G13\       <= \54149\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WL13\      <= \54152\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WL13/\     <= \54154\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \RL13/\     <= \54157\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WHOMP/\    <= \54161\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \XUY14/\    <= \54210\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \SUMA14/\   <= \54212\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \CI15/\     <= \54214\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \SUMB14/\   <= \54215\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \A14/\      <= \54220\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \L14/\      <= \54226\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \Z14/\      <= \54235\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \G14/\      <= \54248\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \G14\       <= \54249\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WL14\      <= \54252\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WL14/\     <= \54254\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \RL14/\     <= \54257\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \GTRST/\    <= \54261\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \WHOMP\     <= \54262\    ; -- A11/1 - 4 BIT MODULE (4 OF 4).
  \XUY16/\    <= \54310\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \SUMA16/\   <= \54312\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \EAC/\      <= \54314\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \SUMB16/\   <= \54315\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \A16/\      <= \54320\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \L16/\      <= \54326\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \RL16\      <= \54328\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \Z16/\      <= \54335\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \G16/\      <= \54348\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \G16\       <= \54349\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \WL16\      <= \54352\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \WL16/\     <= \54354\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \RL16/\     <= \54357\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \PIPAZ+/\   <= \54361\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \PIPAZ-/\   <= \54362\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \CO02\      <= \54401\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \XUY15/\    <= \54410\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \SUMA15/\   <= \54412\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \CI16/\     <= \54414\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \SUMB15/\   <= \54415\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \A15/\      <= \54420\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \L15/\      <= \54426\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \Z15/\      <= \54435\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \G15/\      <= \54448\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \G15\       <= \54449\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \WL15\      <= \54452\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \WL15/\     <= \54454\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \RL15/\     <= \54457\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \PIPAY-/\   <= \54461\    ; -- A11/2 - 4 BIT MODULE (4 OF 4).
  \G01A/\     <= \34101\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA03\      <= \34108\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA03/\     <= \34110\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA06\      <= \34118\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA06/\     <= \34120\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA09\      <= \34129\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA09/\     <= \34131\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA12\      <= \34140\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA12/\     <= \34143\    ; -- A12/1 - PARITY AND S REGISTER.
  \G16A/\     <= \34146\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA15\      <= \34151\    ; -- A12/1 - PARITY AND S REGISTER.
  \PA15/\     <= \34153\    ; -- A12/1 - PARITY AND S REGISTER.
  \GNZRO\     <= \34155\    ; -- A12/1 - PARITY AND S REGISTER.
  \EXTPLS\    <= \34205\    ; -- A12/1 - PARITY AND S REGISTER.
  \RELPLS\    <= \34206\    ; -- A12/1 - PARITY AND S REGISTER.
  \RADRZ\     <= \34212\    ; -- A12/1 - PARITY AND S REGISTER.
  \RADRG\     <= \34213\    ; -- A12/1 - PARITY AND S REGISTER.
  \INHPLS\    <= \34215\    ; -- A12/1 - PARITY AND S REGISTER.
  \GEQZRO/\   <= \34218\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD09\     <= \34221\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD10\     <= \34222\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD11\     <= \34223\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD09/\    <= \34224\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD10/\    <= \34225\    ; -- A12/1 - PARITY AND S REGISTER.
  \EAD11/\    <= \34226\    ; -- A12/1 - PARITY AND S REGISTER.
  \PB09\      <= \34231\    ; -- A12/1 - PARITY AND S REGISTER.
  \PB09/\     <= \34233\    ; -- A12/1 - PARITY AND S REGISTER.
  \PB15\      <= \34236\    ; -- A12/1 - PARITY AND S REGISTER.
  \PB15/\     <= \34237\    ; -- A12/1 - PARITY AND S REGISTER.
  \PC15\      <= \34240\    ; -- A12/1 - PARITY AND S REGISTER.
  \PC15/\     <= \34242\    ; -- A12/1 - PARITY AND S REGISTER.
  \PALE\      <= \34251\    ; -- A12/1 - PARITY AND S REGISTER.
  \BRXP3\     <= \34253\    ; -- A12/1 - PARITY AND S REGISTER.
  \G01ED\     <= \34301\    ; -- A12/2 - PARITY AND S REGISTER.
  \S08\       <= \34306\    ; -- A12/2 - PARITY AND S REGISTER.
  \S08/\      <= \34307\    ; -- A12/2 - PARITY AND S REGISTER.
  \G02ED\     <= \34309\    ; -- A12/2 - PARITY AND S REGISTER.
  \S09\       <= \34314\    ; -- A12/2 - PARITY AND S REGISTER.
  \S09/\      <= \34315\    ; -- A12/2 - PARITY AND S REGISTER.
  \G03ED\     <= \34317\    ; -- A12/2 - PARITY AND S REGISTER.
  \S10\       <= \34322\    ; -- A12/2 - PARITY AND S REGISTER.
  \S10/\      <= \34323\    ; -- A12/2 - PARITY AND S REGISTER.
  \G04ED\     <= \34325\    ; -- A12/2 - PARITY AND S REGISTER.
  \T12A\      <= \34329\    ; -- A12/2 - PARITY AND S REGISTER.
  \S11\       <= \34330\    ; -- A12/2 - PARITY AND S REGISTER.
  \S11/\      <= \34331\    ; -- A12/2 - PARITY AND S REGISTER.
  \G05ED\     <= \34333\    ; -- A12/2 - PARITY AND S REGISTER.
  \S12\       <= \34338\    ; -- A12/2 - PARITY AND S REGISTER.
  \S12/\      <= \34339\    ; -- A12/2 - PARITY AND S REGISTER.
  \SHIFT/\    <= \34340\    ; -- A12/2 - PARITY AND S REGISTER.
  \G06ED\     <= \34341\    ; -- A12/2 - PARITY AND S REGISTER.
  \G07ED\     <= \34342\    ; -- A12/2 - PARITY AND S REGISTER.
  \CYR/\      <= \34348\    ; -- A12/2 - PARITY AND S REGISTER.
  \SR/\       <= \34350\    ; -- A12/2 - PARITY AND S REGISTER.
  \CYL/\      <= \34352\    ; -- A12/2 - PARITY AND S REGISTER.
  \EDOP/\     <= \34354\    ; -- A12/2 - PARITY AND S REGISTER.
  \GINH\      <= \34358\    ; -- A12/2 - PARITY AND S REGISTER.
  \SHIFT\     <= \34362\    ; -- A12/2 - PARITY AND S REGISTER.
  \S01\       <= \34404\    ; -- A12/2 - PARITY AND S REGISTER.
  \S01/\      <= \34406\    ; -- A12/2 - PARITY AND S REGISTER.
  \S02\       <= \34411\    ; -- A12/2 - PARITY AND S REGISTER.
  \S02/\      <= \34413\    ; -- A12/2 - PARITY AND S REGISTER.
  \S03\       <= \34418\    ; -- A12/2 - PARITY AND S REGISTER.
  \S03/\      <= \34420\    ; -- A12/2 - PARITY AND S REGISTER.
  \S04\       <= \34425\    ; -- A12/2 - PARITY AND S REGISTER.
  \S04/\      <= \34427\    ; -- A12/2 - PARITY AND S REGISTER.
  \S05\       <= \34432\    ; -- A12/2 - PARITY AND S REGISTER.
  \S05/\      <= \34434\    ; -- A12/2 - PARITY AND S REGISTER.
  \S06\       <= \34439\    ; -- A12/2 - PARITY AND S REGISTER.
  \S06/\      <= \34441\    ; -- A12/2 - PARITY AND S REGISTER.
  \WGA/\      <= \34446\    ; -- A12/2 - PARITY AND S REGISTER.
  \S07\       <= \34447\    ; -- A12/2 - PARITY AND S REGISTER.
  \S07/\      <= \34449\    ; -- A12/2 - PARITY AND S REGISTER.
  \L02A/\     <= \34463\    ; -- A12/2 - PARITY AND S REGISTER.
  \L15A/\     <= \34465\    ; -- A12/2 - PARITY AND S REGISTER.
  \G01A\      <= \34466\    ; -- A12/2 - PARITY AND S REGISTER.
  \MSTRTP\    <= \41105\    ; -- A13/1 - ALARMS.
  \CKTAL/\    <= \41117\    ; -- A13/1 - ALARMS.
  \ALGA\      <= \41118\    ; -- A13/1 - ALARMS.
  \G16SW/\    <= \41131\    ; -- A13/1 - ALARMS.
  \CTPLS/\    <= \41134\    ; -- A13/1 - ALARMS.
  \DOFILT\    <= \41147\    ; -- A13/1 - ALARMS.
  \DLKPLS\    <= \41154\    ; -- A13/1 - ALARMS.
  \SYNC4/\    <= \41219\    ; -- A13/1 - ALARMS.
  \SYNC14/\   <= \41221\    ; -- A13/1 - ALARMS.
  \AGCWAR\    <= \41226\    ; -- A13/1 - ALARMS.
  \WARN\      <= \41227\    ; -- A13/1 - ALARMS.
  \CGCWAR\    <= \41228\    ; -- A13/1 - ALARMS.
  \TMPCAU\    <= \41230\    ; -- A13/1 - ALARMS.
  \OSCALM\    <= \41233\    ; -- A13/1 - ALARMS.
  \SBYEXT\    <= \41236\    ; -- A13/1 - ALARMS.
  \RESTRT\    <= \41240\    ; -- A13/1 - ALARMS.
  \F08B/\     <= \41241\    ; -- A13/1 - ALARMS.
  \CON3\      <= \41242\    ; -- A13/1 - ALARMS.
  \SCADBL\    <= \41243\    ; -- A13/1 - ALARMS.
  \STRT1\     <= \41246\    ; -- A13/1 - ALARMS.
  \ROP/\      <= \42101\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \SETAB/\    <= \42116\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \SETCD/\    <= \42117\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \SBFSET\    <= \42122\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \STBF\      <= \42124\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \TPGF\      <= \42143\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \STRGAT\    <= \42146\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \WHOMPA\    <= \42157\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \RSTK/\     <= \42219\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \FNERAS/\   <= \42225\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \REDRST\    <= \42241\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \SBESET\    <= \42245\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \STBE\      <= \42247\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \TPGE\      <= \42248\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \TPARG/\    <= \42249\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \ERAS/\     <= \42252\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \ERAS\      <= \42254\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \NOTEST/\   <= \42257\    ; -- A14/1 - MEMORY TIMING & ADDRESSING.
  \XB0\       <= \42301\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB0/\      <= \42302\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB1\       <= \42307\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB1/\      <= \42308\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB2\       <= \42312\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB2/\      <= \42313\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB3\       <= \42317\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB3/\      <= \42318\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB4\       <= \42322\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB4/\      <= \42323\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB5\       <= \42327\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB5/\      <= \42328\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB6\       <= \42332\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB6/\      <= \42333\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB7\       <= \42337\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XB7/\      <= \42339\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB0\       <= \42342\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB0/\      <= \42343\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB1\       <= \42346\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB1/\      <= \42347\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB2\       <= \42349\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB2/\      <= \42350\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB3\       <= \42352\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \YB3/\      <= \42353\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \RILP1\     <= \42355\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \RILP1/\    <= \42356\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \CXB1/\     <= \42357\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT0\       <= \42401\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT0/\      <= \42402\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT1\       <= \42405\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT1/\      <= \42406\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT2\       <= \42409\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT2/\      <= \42410\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT3\       <= \42413\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT3/\      <= \42414\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT4\       <= \42417\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT4/\      <= \42418\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT5\       <= \42421\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT5/\      <= \42423\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT6\       <= \42425\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \RB1\       <= \42426\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT6/\      <= \42427\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT7\       <= \42429\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \XT7/\      <= \42431\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \RSCG/\     <= \42449\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \WSCG/\     <= \42452\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \R1C\       <= \42454\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \NOTEST\    <= \42459\    ; -- A14/2 - MEMORY TIMING & ADDRESSING.
  \FB16/\     <= \35102\    ; -- A15/1 - RUPT SERVICE.
  \FB16\      <= \35104\    ; -- A15/1 - RUPT SERVICE.
  \BK16\      <= \35105\    ; -- A15/1 - RUPT SERVICE.
  \FB14/\     <= \35108\    ; -- A15/1 - RUPT SERVICE.
  \FB14\      <= \35110\    ; -- A15/1 - RUPT SERVICE.
  \FB13/\     <= \35114\    ; -- A15/1 - RUPT SERVICE.
  \FB13\      <= \35115\    ; -- A15/1 - RUPT SERVICE.
  \FB12/\     <= \35119\    ; -- A15/1 - RUPT SERVICE.
  \FB12\      <= \35120\    ; -- A15/1 - RUPT SERVICE.
  \FB11/\     <= \35124\    ; -- A15/1 - RUPT SERVICE.
  \FB11\      <= \35125\    ; -- A15/1 - RUPT SERVICE.
  \EB11/\     <= \35130\    ; -- A15/1 - RUPT SERVICE.
  \EB11\      <= \35131\    ; -- A15/1 - RUPT SERVICE.
  \BBK3\      <= \35133\    ; -- A15/1 - RUPT SERVICE.
  \EB10/\     <= \35137\    ; -- A15/1 - RUPT SERVICE.
  \EB10\      <= \35138\    ; -- A15/1 - RUPT SERVICE.
  \BBK2\      <= \35140\    ; -- A15/1 - RUPT SERVICE.
  \EB9/\      <= \35145\    ; -- A15/1 - RUPT SERVICE.
  \EB9\       <= \35146\    ; -- A15/1 - RUPT SERVICE.
  \BBK1\      <= \35148\    ; -- A15/1 - RUPT SERVICE.
  \F11/\      <= \35205\    ; -- A15/1 - RUPT SERVICE.
  \F11\       <= \35206\    ; -- A15/1 - RUPT SERVICE.
  \F13\       <= \35207\    ; -- A15/1 - RUPT SERVICE.
  \F12/\      <= \35208\    ; -- A15/1 - RUPT SERVICE.
  \F12\       <= \35209\    ; -- A15/1 - RUPT SERVICE.
  \F13/\      <= \35210\    ; -- A15/1 - RUPT SERVICE.
  \F16\       <= \35213\    ; -- A15/1 - RUPT SERVICE.
  \F14\       <= \35215\    ; -- A15/1 - RUPT SERVICE.
  \F15\       <= \35216\    ; -- A15/1 - RUPT SERVICE.
  \F14/\      <= \35217\    ; -- A15/1 - RUPT SERVICE.
  \F15/\      <= \35218\    ; -- A15/1 - RUPT SERVICE.
  \F16/\      <= \35219\    ; -- A15/1 - RUPT SERVICE.
  \PRPOR3\    <= \35226\    ; -- A15/1 - RUPT SERVICE.
  \PRPOR4\    <= \35227\    ; -- A15/1 - RUPT SERVICE.
  \RPTAD6\    <= \35232\    ; -- A15/1 - RUPT SERVICE.
  \RPTA12\    <= \35233\    ; -- A15/1 - RUPT SERVICE.
  \RUPTOR/\   <= \35235\    ; -- A15/1 - RUPT SERVICE.
  \MINC/\     <= \35239\    ; -- A15/1 - RUPT SERVICE.
  \MINC\      <= \35240\    ; -- A15/1 - RUPT SERVICE.
  \PCDU/\     <= \35244\    ; -- A15/1 - RUPT SERVICE.
  \PCDU\      <= \35245\    ; -- A15/1 - RUPT SERVICE.
  \MCDU/\     <= \35249\    ; -- A15/1 - RUPT SERVICE.
  \MCDU\      <= \35250\    ; -- A15/1 - RUPT SERVICE.
  \WOVR/\     <= \35301\    ; -- A15/2 - RUPT SERVICE.
  \KRPTA/\    <= \35304\    ; -- A15/2 - RUPT SERVICE.
  \T6RPT\     <= \35307\    ; -- A15/2 - RUPT SERVICE.
  \KY1RST\    <= \35327\    ; -- A15/2 - RUPT SERVICE.
  \KY2RST\    <= \35333\    ; -- A15/2 - RUPT SERVICE.
  \PRPOR1\    <= \35344\    ; -- A15/2 - RUPT SERVICE.
  \DRPRST\    <= \35345\    ; -- A15/2 - RUPT SERVICE.
  \DNRPTA\    <= \35347\    ; -- A15/2 - RUPT SERVICE.
  \PRPOR2\    <= \35348\    ; -- A15/2 - RUPT SERVICE.
  \RRPA1/\    <= \35349\    ; -- A15/2 - RUPT SERVICE.
  \RPTAD3\    <= \35352\    ; -- A15/2 - RUPT SERVICE.
  \RPTAD4\    <= \35355\    ; -- A15/2 - RUPT SERVICE.
  \RPTAD5\    <= \35358\    ; -- A15/2 - RUPT SERVICE.
  \RC+X+P\    <= \43105\    ; -- A16/1 - INOUT I.
  \RC-X-P\    <= \43111\    ; -- A16/1 - INOUT I.
  \RC-X+P\    <= \43117\    ; -- A16/1 - INOUT I.
  \RC+X-P\    <= \43123\    ; -- A16/1 - INOUT I.
  \RC+X+Y\    <= \43129\    ; -- A16/1 - INOUT I.
  \RC-X-Y\    <= \43135\    ; -- A16/1 - INOUT I.
  \RC-X+Y\    <= \43141\    ; -- A16/1 - INOUT I.
  \RC+X-Y\    <= \43147\    ; -- A16/1 - INOUT I.
  \WCH05/\    <= \43149\    ; -- A16/1 - INOUT I.
  \CCH05\     <= \43154\    ; -- A16/1 - INOUT I.
  \CH1208\    <= \43159\    ; -- A16/1 - INOUT I.
  \TVCNAB\    <= \43160\    ; -- A16/1 - INOUT I.
  \RC+Y-R\    <= \43205\    ; -- A16/1 - INOUT I.
  \WCH06/\    <= \43207\    ; -- A16/1 - INOUT I.
  \CCH06\     <= \43211\    ; -- A16/1 - INOUT I.
  \RCH06/\    <= \43214\    ; -- A16/1 - INOUT I.
  \RCH05/\    <= \43217\    ; -- A16/1 - INOUT I.
  \RC-Y+R\    <= \43223\    ; -- A16/1 - INOUT I.
  \CH1207\    <= \43227\    ; -- A16/1 - INOUT I.
  \OT1207\    <= \43228\    ; -- A16/1 - INOUT I.
  \OT1207/\   <= \43229\    ; -- A16/1 - INOUT I.
  \RC-Y-R\    <= \43234\    ; -- A16/1 - INOUT I.
  \RC+Y+R\    <= \43239\    ; -- A16/1 - INOUT I.
  \RC+Z-R\    <= \43244\    ; -- A16/1 - INOUT I.
  \RC-Z+R\    <= \43249\    ; -- A16/1 - INOUT I.
  \RC-Z-R\    <= \43254\    ; -- A16/1 - INOUT I.
  \RC+Z+R\    <= \43259\    ; -- A16/1 - INOUT I.
  \ZOPCDU\    <= \43302\    ; -- A16/2 - INOUT I.
  \ENEROP\    <= \43310\    ; -- A16/2 - INOUT I.
  \STARON\    <= \43312\    ; -- A16/2 - INOUT I.
  \COARSE\    <= \43320\    ; -- A16/2 - INOUT I.
  \ZIMCDU\    <= \43322\    ; -- A16/2 - INOUT I.
  \ENERIM\    <= \43330\    ; -- A16/2 - INOUT I.
  \CH1209\    <= \43331\    ; -- A16/2 - INOUT I.
  \S4BTAK\    <= \43332\    ; -- A16/2 - INOUT I.
  \CH1210\    <= \43339\    ; -- A16/2 - INOUT I.
  \ZEROPT\    <= \43340\    ; -- A16/2 - INOUT I.
  \CH1211\    <= \43341\    ; -- A16/2 - INOUT I.
  \DISDAC\    <= \43342\    ; -- A16/2 - INOUT I.
  \WCH12/\    <= \43346\    ; -- A16/2 - INOUT I.
  \CCH12\     <= \43352\    ; -- A16/2 - INOUT I.
  \RCH12/\    <= \43356\    ; -- A16/2 - INOUT I.
  \ISSWAR\    <= \43401\    ; -- A16/2 - INOUT I.
  \COMACT\    <= \43412\    ; -- A16/2 - INOUT I.
  \UPLACT\    <= \43413\    ; -- A16/2 - INOUT I.
  \TMPOUT\    <= \43424\    ; -- A16/2 - INOUT I.
  \KYRLS\     <= \43427\    ; -- A16/2 - INOUT I.
  \VNFLSH\    <= \43435\    ; -- A16/2 - INOUT I.
  \OPEROR\    <= \43441\    ; -- A16/2 - INOUT I.
  \CH1212\    <= \43449\    ; -- A16/2 - INOUT I.
  \MROLGT\    <= \43450\    ; -- A16/2 - INOUT I.
  \S4BSEQ\    <= \43451\    ; -- A16/2 - INOUT I.
  \CH1213\    <= \43452\    ; -- A16/2 - INOUT I.
  \CH1214\    <= \43459\    ; -- A16/2 - INOUT I.
  \S4BOFF\    <= \43460\    ; -- A16/2 - INOUT I.
  \CHOR01/\   <= \44103\    ; -- A17/1 - INOUT II.
  \CHOR02/\   <= \44106\    ; -- A17/1 - INOUT II.
  \CHOR03/\   <= \44109\    ; -- A17/1 - INOUT II.
  \CHOR04/\   <= \44112\    ; -- A17/1 - INOUT II.
  \CHOR05/\   <= \44115\    ; -- A17/1 - INOUT II.
  \CHOR06/\   <= \44118\    ; -- A17/1 - INOUT II.
  \CHOR07/\   <= \44121\    ; -- A17/1 - INOUT II.
  \CHOR08/\   <= \44124\    ; -- A17/1 - INOUT II.
  \CHOR09/\   <= \44127\    ; -- A17/1 - INOUT II.
  \CHOR10/\   <= \44129\    ; -- A17/1 - INOUT II.
  \CHOR11/\   <= \44132\    ; -- A17/1 - INOUT II.
  \CHOR12/\   <= \44135\    ; -- A17/1 - INOUT II.
  \CHOR13/\   <= \44138\    ; -- A17/1 - INOUT II.
  \CHOR14/\   <= \44141\    ; -- A17/1 - INOUT II.
  \CHOR16/\   <= \44144\    ; -- A17/1 - INOUT II.
  \RCH30/\    <= \44146\    ; -- A17/1 - INOUT II.
  \RCH31/\    <= \44150\    ; -- A17/1 - INOUT II.
  \RCH32/\    <= \44154\    ; -- A17/1 - INOUT II.
  \RCH33/\    <= \44158\    ; -- A17/1 - INOUT II.
  \TRP31A\    <= \44211\    ; -- A17/1 - INOUT II.
  \TRP31B\    <= \44226\    ; -- A17/1 - INOUT II.
  \HNDRPT\    <= \44231\    ; -- A17/1 - INOUT II.
  \CH3201\    <= \44236\    ; -- A17/1 - INOUT II.
  \CH3206\    <= \44237\    ; -- A17/1 - INOUT II.
  \CH3202\    <= \44238\    ; -- A17/1 - INOUT II.
  \CH3207\    <= \44239\    ; -- A17/1 - INOUT II.
  \CH3203\    <= \44240\    ; -- A17/1 - INOUT II.
  \CH3208\    <= \44241\    ; -- A17/1 - INOUT II.
  \CH3204\    <= \44242\    ; -- A17/1 - INOUT II.
  \CH3209\    <= \44243\    ; -- A17/1 - INOUT II.
  \CH3205\    <= \44244\    ; -- A17/1 - INOUT II.
  \CH3210\    <= \44245\    ; -- A17/1 - INOUT II.
  \TRP32\     <= \44253\    ; -- A17/1 - INOUT II.
  \CH3316\    <= \44257\    ; -- A17/1 - INOUT II.
  \CH3314\    <= \44258\    ; -- A17/1 - INOUT II.
  \CH3313\    <= \44259\    ; -- A17/1 - INOUT II.
  \RLYB01\    <= \44305\    ; -- A17/2 - INOUT II.
  \RLYB02\    <= \44311\    ; -- A17/2 - INOUT II.
  \RLYB03\    <= \44317\    ; -- A17/2 - INOUT II.
  \RLYB04\    <= \44323\    ; -- A17/2 - INOUT II.
  \RLYB05\    <= \44329\    ; -- A17/2 - INOUT II.
  \RLYB06\    <= \44335\    ; -- A17/2 - INOUT II.
  \RLYB07\    <= \44341\    ; -- A17/2 - INOUT II.
  \RLYB08\    <= \44347\    ; -- A17/2 - INOUT II.
  \RLYB09\    <= \44353\    ; -- A17/2 - INOUT II.
  \RLYB10\    <= \44359\    ; -- A17/2 - INOUT II.
  \RLYB11\    <= \44405\    ; -- A17/2 - INOUT II.
  \RYWD12\    <= \44411\    ; -- A17/2 - INOUT II.
  \RYWD13\    <= \44417\    ; -- A17/2 - INOUT II.
  \RYWD14\    <= \44423\    ; -- A17/2 - INOUT II.
  \RYWD16\    <= \44429\    ; -- A17/2 - INOUT II.
  \WCH10/\    <= \44432\    ; -- A17/2 - INOUT II.
  \CCH10\     <= \44437\    ; -- A17/2 - INOUT II.
  \RCH10/\    <= \44441\    ; -- A17/2 - INOUT II.
  \WCH11/\    <= \44445\    ; -- A17/2 - INOUT II.
  \CCH11\     <= \44450\    ; -- A17/2 - INOUT II.
  \RCH11/\    <= \44454\    ; -- A17/2 - INOUT II.
  \XBC\       <= \44462\    ; -- A17/2 - INOUT II.
  \CH1501\    <= \45103\    ; -- A18/1 - INOUT III.
  \CH1502\    <= \45107\    ; -- A18/1 - INOUT III.
  \CH1503\    <= \45111\    ; -- A18/1 - INOUT III.
  \CH1504\    <= \45115\    ; -- A18/1 - INOUT III.
  \CH1505\    <= \45119\    ; -- A18/1 - INOUT III.
  \RCH15/\    <= \45124\    ; -- A18/1 - INOUT III.
  \TPOR/\     <= \45128\    ; -- A18/1 - INOUT III.
  \KYRPT1\    <= \45131\    ; -- A18/1 - INOUT III.
  \CH1311\    <= \45140\    ; -- A18/1 - INOUT III.
  \SBY\       <= \45148\    ; -- A18/1 - INOUT III.
  \STNDBY/\   <= \45153\    ; -- A18/1 - INOUT III.
  \STNDBY\    <= \45155\    ; -- A18/1 - INOUT III.
  \SBYLIT\    <= \45157\    ; -- A18/1 - INOUT III.
  \F17A/\     <= \45159\    ; -- A18/1 - INOUT III.
  \CH1601\    <= \45203\    ; -- A18/1 - INOUT III.
  \CH1602\    <= \45207\    ; -- A18/1 - INOUT III.
  \CH1603\    <= \45211\    ; -- A18/1 - INOUT III.
  \CH1604\    <= \45215\    ; -- A18/1 - INOUT III.
  \CH1605\    <= \45219\    ; -- A18/1 - INOUT III.
  \ERRST\     <= \45224\    ; -- A18/1 - INOUT III.
  \CH1606\    <= \45227\    ; -- A18/1 - INOUT III.
  \CH1607\    <= \45231\    ; -- A18/1 - INOUT III.
  \RCH16/\    <= \45236\    ; -- A18/1 - INOUT III.
  \KYRPT2\    <= \45244\    ; -- A18/1 - INOUT III.
  \MKRPT\     <= \45254\    ; -- A18/1 - INOUT III.
  \F17B/\     <= \45261\    ; -- A18/1 - INOUT III.
  \TEMPIN/\   <= \45262\    ; -- A18/1 - INOUT III.
  \CH1304\    <= \45304\    ; -- A18/2 - INOUT III.
  \CH1303\    <= \45309\    ; -- A18/2 - INOUT III.
  \CH1302\    <= \45315\    ; -- A18/2 - INOUT III.
  \CH1301\    <= \45319\    ; -- A18/2 - INOUT III.
  \RRRANG\    <= \45328\    ; -- A18/2 - INOUT III.
  \RRRARA\    <= \45329\    ; -- A18/2 - INOUT III.
  \LRXVEL\    <= \45330\    ; -- A18/2 - INOUT III.
  \LRYVEL\    <= \45331\    ; -- A18/2 - INOUT III.
  \LRZVEL\    <= \45332\    ; -- A18/2 - INOUT III.
  \LRRANG\    <= \45333\    ; -- A18/2 - INOUT III.
  \RADRPT\    <= \45342\    ; -- A18/2 - INOUT III.
  \RRSYNC\    <= \45345\    ; -- A18/2 - INOUT III.
  \LRSYNC\    <= \45346\    ; -- A18/2 - INOUT III.
  \RNRADP\    <= \45352\    ; -- A18/2 - INOUT III.
  \RNRADM\    <= \45358\    ; -- A18/2 - INOUT III.
  \TPORA/\    <= \45359\    ; -- A18/2 - INOUT III.
  \HERB\      <= \45360\    ; -- A18/2 - INOUT III.
  \F10AS0\    <= \45401\    ; -- A18/2 - INOUT III.
  \CNTOF9\    <= \45434\    ; -- A18/2 - INOUT III.
  \CH11\      <= \45437\    ; -- A18/2 - INOUT III.
  \CH12\      <= \45440\    ; -- A18/2 - INOUT III.
  \CH13\      <= \45442\    ; -- A18/2 - INOUT III.
  \CH14\      <= \45444\    ; -- A18/2 - INOUT III.
  \CH16\      <= \45446\    ; -- A18/2 - INOUT III.
  \END\       <= \45448\    ; -- A18/2 - INOUT III.
  \DLKRPT\    <= \45449\    ; -- A18/2 - INOUT III.
  \CH3312\    <= \45456\    ; -- A18/2 - INOUT III.
  \SH3MS/\    <= \46102\    ; -- A19/1 - INOUT IV.
  \ALT0\      <= \46109\    ; -- A19/1 - INOUT IV.
  \ALT1\      <= \46110\    ; -- A19/1 - INOUT IV.
  \ALRT0\     <= \46111\    ; -- A19/1 - INOUT IV.
  \ALRT1\     <= \46112\    ; -- A19/1 - INOUT IV.
  \CH1402\    <= \46116\    ; -- A19/1 - INOUT IV.
  \CH1403\    <= \46120\    ; -- A19/1 - INOUT IV.
  \ALTM\      <= \46129\    ; -- A19/1 - INOUT IV.
  \ALTSNC\    <= \46132\    ; -- A19/1 - INOUT IV.
  \OTLNKM\    <= \46143\    ; -- A19/1 - INOUT IV.
  \CH1401\    <= \46145\    ; -- A19/1 - INOUT IV.
  \OTLNK0\    <= \46147\    ; -- A19/1 - INOUT IV.
  \OTLNK1\    <= \46149\    ; -- A19/1 - INOUT IV.
  \F5ASB0\    <= \46152\    ; -- A19/1 - INOUT IV.
  \F5ASB0/\   <= \46153\    ; -- A19/1 - INOUT IV.
  \F5ASB2\    <= \46154\    ; -- A19/1 - INOUT IV.
  \F5ASB2/\   <= \46155\    ; -- A19/1 - INOUT IV.
  \F5BSB2\    <= \46156\    ; -- A19/1 - INOUT IV.
  \F5BSB2/\   <= \46157\    ; -- A19/1 - INOUT IV.
  \T2P\       <= \46160\    ; -- A19/1 - INOUT IV.
  \INLNKM\    <= \46203\    ; -- A19/1 - INOUT IV.
  \INLNKP\    <= \46206\    ; -- A19/1 - INOUT IV.
  \CCH33\     <= \46212\    ; -- A19/1 - INOUT IV.
  \CH3311\    <= \46215\    ; -- A19/1 - INOUT IV.
  \C45R/\     <= \46220\    ; -- A19/1 - INOUT IV.
  \CH3310\    <= \46221\    ; -- A19/1 - INOUT IV.
  \CH1305\    <= \46228\    ; -- A19/1 - INOUT IV.
  \CH1306\    <= \46229\    ; -- A19/1 - INOUT IV.
  \CH1404\    <= \46233\    ; -- A19/1 - INOUT IV.
  \THRSTD\    <= \46234\    ; -- A19/1 - INOUT IV.
  \CH1405\    <= \46238\    ; -- A19/1 - INOUT IV.
  \EMSD\      <= \46239\    ; -- A19/1 - INOUT IV.
  \THRST+\    <= \46247\    ; -- A19/1 - INOUT IV.
  \THRST-\    <= \46248\    ; -- A19/1 - INOUT IV.
  \EMS+\      <= \46254\    ; -- A19/1 - INOUT IV.
  \EMS-\      <= \46258\    ; -- A19/1 - INOUT IV.
  \UPRUPT\    <= \46303\    ; -- A19/2 - INOUT IV.
  \UPL0/\     <= \46304\    ; -- A19/2 - INOUT IV.
  \UPL1/\     <= \46305\    ; -- A19/2 - INOUT IV.
  \XLNK0/\    <= \46306\    ; -- A19/2 - INOUT IV.
  \XLNK1/\    <= \46307\    ; -- A19/2 - INOUT IV.
  \BLKUPL\    <= \46308\    ; -- A19/2 - INOUT IV.
  \F10B/\     <= \46309\    ; -- A19/2 - INOUT IV.
  \T1P\       <= \46310\    ; -- A19/2 - INOUT IV.
  \T3P\       <= \46311\    ; -- A19/2 - INOUT IV.
  \F09B/\     <= \46312\    ; -- A19/2 - INOUT IV.
  \T4P\       <= \46313\    ; -- A19/2 - INOUT IV.
  \F10A/\     <= \46314\    ; -- A19/2 - INOUT IV.
  \T5P\       <= \46315\    ; -- A19/2 - INOUT IV.
  \F06B/\     <= \46316\    ; -- A19/2 - INOUT IV.
  \T6P\       <= \46317\    ; -- A19/2 - INOUT IV.
  \CH1308\    <= \46321\    ; -- A19/2 - INOUT IV.
  \CH1309\    <= \46326\    ; -- A19/2 - INOUT IV.
  \RHCGO\     <= \46330\    ; -- A19/2 - INOUT IV.
  \BMAGXP\    <= \46339\    ; -- A19/2 - INOUT IV.
  \BMAGXM\    <= \46340\    ; -- A19/2 - INOUT IV.
  \BMAGYP\    <= \46348\    ; -- A19/2 - INOUT IV.
  \BMAGYM\    <= \46349\    ; -- A19/2 - INOUT IV.
  \BMAGZP\    <= \46358\    ; -- A19/2 - INOUT IV.
  \BMAGZM\    <= \46359\    ; -- A19/2 - INOUT IV.
  \CH1410\    <= \46404\    ; -- A19/2 - INOUT IV.
  \GYROD\     <= \46405\    ; -- A19/2 - INOUT IV.
  \CH1409\    <= \46409\    ; -- A19/2 - INOUT IV.
  \CH1408\    <= \46413\    ; -- A19/2 - INOUT IV.
  \CH1407\    <= \46417\    ; -- A19/2 - INOUT IV.
  \CH1406\    <= \46421\    ; -- A19/2 - INOUT IV.
  \GYXP\      <= \46424\    ; -- A19/2 - INOUT IV.
  \GYXM\      <= \46425\    ; -- A19/2 - INOUT IV.
  \GYYP\      <= \46426\    ; -- A19/2 - INOUT IV.
  \GYYM\      <= \46427\    ; -- A19/2 - INOUT IV.
  \GYZP\      <= \46432\    ; -- A19/2 - INOUT IV.
  \GYZM\      <= \46433\    ; -- A19/2 - INOUT IV.
  \GYENAB\    <= \46434\    ; -- A19/2 - INOUT IV.
  \GYRSET\    <= \46442\    ; -- A19/2 - INOUT IV.
  \GYRRST\    <= \46443\    ; -- A19/2 - INOUT IV.
  \FF1109/\   <= \46445\    ; -- A19/2 - INOUT IV.
  \FF1109\    <= \46446\    ; -- A19/2 - INOUT IV.
  \CH1109\    <= \46447\    ; -- A19/2 - INOUT IV.
  \W1110\     <= \46448\    ; -- A19/2 - INOUT IV.
  \FF1110/\   <= \46449\    ; -- A19/2 - INOUT IV.
  \FF1110\    <= \46450\    ; -- A19/2 - INOUT IV.
  \CH1110\    <= \46451\    ; -- A19/2 - INOUT IV.
  \FF1111/\   <= \46453\    ; -- A19/2 - INOUT IV.
  \FF1111\    <= \46454\    ; -- A19/2 - INOUT IV.
  \CH1111\    <= \46455\    ; -- A19/2 - INOUT IV.
  \FF1112/\   <= \46457\    ; -- A19/2 - INOUT IV.
  \FF1112\    <= \46458\    ; -- A19/2 - INOUT IV.
  \CH1112\    <= \46459\    ; -- A19/2 - INOUT IV.
  \C32A\      <= \31108\    ; -- A20/1 - COUNTER CELL I.
  \C32R\      <= \31112\    ; -- A20/1 - COUNTER CELL I.
  \C32P\      <= \31113\    ; -- A20/1 - COUNTER CELL I.
  \C32M\      <= \31114\    ; -- A20/1 - COUNTER CELL I.
  \C33A\      <= \31121\    ; -- A20/1 - COUNTER CELL I.
  \CG11\      <= \31123\    ; -- A20/1 - COUNTER CELL I.
  \C33R\      <= \31126\    ; -- A20/1 - COUNTER CELL I.
  \C33P\      <= \31127\    ; -- A20/1 - COUNTER CELL I.
  \C33M\      <= \31128\    ; -- A20/1 - COUNTER CELL I.
  \C24A\      <= \31134\    ; -- A20/1 - COUNTER CELL I.
  \C24R\      <= \31135\    ; -- A20/1 - COUNTER CELL I.
  \C25A\      <= \31141\    ; -- A20/1 - COUNTER CELL I.
  \C25R\      <= \31142\    ; -- A20/1 - COUNTER CELL I.
  \C26A\      <= \31149\    ; -- A20/1 - COUNTER CELL I.
  \CG21\      <= \31152\    ; -- A20/1 - COUNTER CELL I.
  \C26R\      <= \31153\    ; -- A20/1 - COUNTER CELL I.
  \CA3/\      <= \31154\    ; -- A20/1 - COUNTER CELL I.
  \CXB7/\     <= \31158\    ; -- A20/1 - COUNTER CELL I.
  \C34A\      <= \31208\    ; -- A20/1 - COUNTER CELL I.
  \C34R\      <= \31212\    ; -- A20/1 - COUNTER CELL I.
  \C34P\      <= \31213\    ; -- A20/1 - COUNTER CELL I.
  \C34M\      <= \31214\    ; -- A20/1 - COUNTER CELL I.
  \C35A\      <= \31221\    ; -- A20/1 - COUNTER CELL I.
  \CG12\      <= \31223\    ; -- A20/1 - COUNTER CELL I.
  \C35R\      <= \31226\    ; -- A20/1 - COUNTER CELL I.
  \C35P\      <= \31227\    ; -- A20/1 - COUNTER CELL I.
  \C35M\      <= \31228\    ; -- A20/1 - COUNTER CELL I.
  \C27A\      <= \31234\    ; -- A20/1 - COUNTER CELL I.
  \C27R\      <= \31235\    ; -- A20/1 - COUNTER CELL I.
  \C30A\      <= \31241\    ; -- A20/1 - COUNTER CELL I.
  \C30R\      <= \31242\    ; -- A20/1 - COUNTER CELL I.
  \C31A\      <= \31249\    ; -- A20/1 - COUNTER CELL I.
  \CG22\      <= \31252\    ; -- A20/1 - COUNTER CELL I.
  \C31R\      <= \31253\    ; -- A20/1 - COUNTER CELL I.
  \CXB2/\     <= \31256\    ; -- A20/1 - COUNTER CELL I.
  \C36A\      <= \31308\    ; -- A20/2 - COUNTER CELL I.
  \C36R\      <= \31312\    ; -- A20/2 - COUNTER CELL I.
  \C36P\      <= \31313\    ; -- A20/2 - COUNTER CELL I.
  \C36M\      <= \31314\    ; -- A20/2 - COUNTER CELL I.
  \C37A\      <= \31321\    ; -- A20/2 - COUNTER CELL I.
  \CG14\      <= \31323\    ; -- A20/2 - COUNTER CELL I.
  \C37R\      <= \31326\    ; -- A20/2 - COUNTER CELL I.
  \C37P\      <= \31327\    ; -- A20/2 - COUNTER CELL I.
  \C37M\      <= \31328\    ; -- A20/2 - COUNTER CELL I.
  \C50A\      <= \31334\    ; -- A20/2 - COUNTER CELL I.
  \C50R\      <= \31335\    ; -- A20/2 - COUNTER CELL I.
  \C51A\      <= \31341\    ; -- A20/2 - COUNTER CELL I.
  \C51R\      <= \31342\    ; -- A20/2 - COUNTER CELL I.
  \C52A\      <= \31349\    ; -- A20/2 - COUNTER CELL I.
  \CG24\      <= \31352\    ; -- A20/2 - COUNTER CELL I.
  \C52R\      <= \31353\    ; -- A20/2 - COUNTER CELL I.
  \CA4/\      <= \31354\    ; -- A20/2 - COUNTER CELL I.
  \CXB3/\     <= \31356\    ; -- A20/2 - COUNTER CELL I.
  \CA2/\      <= \31358\    ; -- A20/2 - COUNTER CELL I.
  \C40A\      <= \31408\    ; -- A20/2 - COUNTER CELL I.
  \C40R\      <= \31412\    ; -- A20/2 - COUNTER CELL I.
  \C40P\      <= \31413\    ; -- A20/2 - COUNTER CELL I.
  \C40M\      <= \31414\    ; -- A20/2 - COUNTER CELL I.
  \C41A\      <= \31421\    ; -- A20/2 - COUNTER CELL I.
  \CG13\      <= \31423\    ; -- A20/2 - COUNTER CELL I.
  \C41R\      <= \31426\    ; -- A20/2 - COUNTER CELL I.
  \C41P\      <= \31427\    ; -- A20/2 - COUNTER CELL I.
  \C41M\      <= \31428\    ; -- A20/2 - COUNTER CELL I.
  \C53A\      <= \31434\    ; -- A20/2 - COUNTER CELL I.
  \C53R\      <= \31435\    ; -- A20/2 - COUNTER CELL I.
  \C54A\      <= \31441\    ; -- A20/2 - COUNTER CELL I.
  \C54R\      <= \31442\    ; -- A20/2 - COUNTER CELL I.
  \C55A\      <= \31449\    ; -- A20/2 - COUNTER CELL I.
  \CG23\      <= \31452\    ; -- A20/2 - COUNTER CELL I.
  \C55R\      <= \31453\    ; -- A20/2 - COUNTER CELL I.
  \CXB4/\     <= \31456\    ; -- A20/2 - COUNTER CELL I.
  \CA6/\      <= \31458\    ; -- A20/2 - COUNTER CELL I.
  \CAD4\      <= \32008\    ; -- A21/1 - COUNTER CELL II.
  \32004K?\   <= \32014\    ; -- A21/1 - COUNTER CELL II.
  \CAD5\      <= \32035\    ; -- A21/1 - COUNTER CELL II.
  \DINC/\     <= \32045\    ; -- A21/1 - COUNTER CELL II.
  \CAD6\      <= \32046\    ; -- A21/1 - COUNTER CELL II.
  \DINC\      <= \32047\    ; -- A21/1 - COUNTER CELL II.
  \DINCNC/\   <= \32048\    ; -- A21/1 - COUNTER CELL II.
  \50SUM\     <= \32050\    ; -- A21/1 - COUNTER CELL II.
  \CAD1\      <= \32051\    ; -- A21/1 - COUNTER CELL II.
  \CAD2\      <= \32052\    ; -- A21/1 - COUNTER CELL II.
  \SHINC/\    <= \32059\    ; -- A21/1 - COUNTER CELL II.
  \SHINC\     <= \32060\    ; -- A21/1 - COUNTER CELL II.
  \CAD3\      <= \32063\    ; -- A21/1 - COUNTER CELL II.
  \30SUM\     <= \32064\    ; -- A21/1 - COUNTER CELL II.
  \SHANC/\    <= \32065\    ; -- A21/1 - COUNTER CELL II.
  \SHANC\     <= \32066\    ; -- A21/1 - COUNTER CELL II.
  \STORE1\    <= \32208\    ; -- A21/2 - COUNTER CELL II.
  \STORE1/\   <= \32209\    ; -- A21/2 - COUNTER CELL II.
  \STFET1/\   <= \32210\    ; -- A21/2 - COUNTER CELL II.
  \MON/\      <= \32215\    ; -- A21/2 - COUNTER CELL II.
  \FETCH1\    <= \32216\    ; -- A21/2 - COUNTER CELL II.
  \FETCH0\    <= \32217\    ; -- A21/2 - COUNTER CELL II.
  \FETCH0/\   <= \32219\    ; -- A21/2 - COUNTER CELL II.
  \INOTLD\    <= \32223\    ; -- A21/2 - COUNTER CELL II.
  \INOTRD\    <= \32227\    ; -- A21/2 - COUNTER CELL II.
  \MON+CH\    <= \32231\    ; -- A21/2 - COUNTER CELL II.
  \INCSET/\   <= \32247\    ; -- A21/2 - COUNTER CELL II.
  \INKL/\     <= \32249\    ; -- A21/2 - COUNTER CELL II.
  \INKL\      <= \32251\    ; -- A21/2 - COUNTER CELL II.
  \RSSB\      <= \32254\    ; -- A21/2 - COUNTER CELL II.
  \BKTF/\     <= \32255\    ; -- A21/2 - COUNTER CELL II.
  \CHINC/\    <= \32256\    ; -- A21/2 - COUNTER CELL II.
  \C42A\      <= \32508\    ; -- A21/3 - COUNTER CELL II.
  \C42R\      <= \32512\    ; -- A21/3 - COUNTER CELL II.
  \C42P\      <= \32513\    ; -- A21/3 - COUNTER CELL II.
  \C42M\      <= \32514\    ; -- A21/3 - COUNTER CELL II.
  \C43A\      <= \32521\    ; -- A21/3 - COUNTER CELL II.
  \CG15\      <= \32523\    ; -- A21/3 - COUNTER CELL II.
  \C43R\      <= \32526\    ; -- A21/3 - COUNTER CELL II.
  \C43P\      <= \32527\    ; -- A21/3 - COUNTER CELL II.
  \C43M\      <= \32528\    ; -- A21/3 - COUNTER CELL II.
  \C56A\      <= \32534\    ; -- A21/3 - COUNTER CELL II.
  \C56R\      <= \32535\    ; -- A21/3 - COUNTER CELL II.
  \C57A\      <= \32541\    ; -- A21/3 - COUNTER CELL II.
  \C57R\      <= \32542\    ; -- A21/3 - COUNTER CELL II.
  \C60A\      <= \32549\    ; -- A21/3 - COUNTER CELL II.
  \CTROR/\    <= \32550\    ; -- A21/3 - COUNTER CELL II.
  \CTROR\     <= \32552\    ; -- A21/3 - COUNTER CELL II.
  \C60R\      <= \32553\    ; -- A21/3 - COUNTER CELL II.
  \CA5/\      <= \32554\    ; -- A21/3 - COUNTER CELL II.
  \CXB5/\     <= \32556\    ; -- A21/3 - COUNTER CELL II.
  \CHINC\     <= \32558\    ; -- A21/3 - COUNTER CELL II.
  \C44A\      <= \32608\    ; -- A21/3 - COUNTER CELL II.
  \C44R\      <= \32612\    ; -- A21/3 - COUNTER CELL II.
  \C44P\      <= \32613\    ; -- A21/3 - COUNTER CELL II.
  \C44M\      <= \32614\    ; -- A21/3 - COUNTER CELL II.
  \C45A\      <= \32621\    ; -- A21/3 - COUNTER CELL II.
  \CG16\      <= \32623\    ; -- A21/3 - COUNTER CELL II.
  \C45R\      <= \32626\    ; -- A21/3 - COUNTER CELL II.
  \C45P\      <= \32627\    ; -- A21/3 - COUNTER CELL II.
  \C45M\      <= \32628\    ; -- A21/3 - COUNTER CELL II.
  \C46A\      <= \32634\    ; -- A21/3 - COUNTER CELL II.
  \C46R\      <= \32635\    ; -- A21/3 - COUNTER CELL II.
  \C46P\      <= \32639\    ; -- A21/3 - COUNTER CELL II.
  \C46M\      <= \32640\    ; -- A21/3 - COUNTER CELL II.
  \C47A\      <= \32649\    ; -- A21/3 - COUNTER CELL II.
  \CG26\      <= \32652\    ; -- A21/3 - COUNTER CELL II.
  \C47R\      <= \32653\    ; -- A21/3 - COUNTER CELL II.
  \CXB0/\     <= \32654\    ; -- A21/3 - COUNTER CELL II.
  \CXB6/\     <= \32656\    ; -- A21/3 - COUNTER CELL II.
  \RQ/\       <= \32658\    ; -- A21/3 - COUNTER CELL II.
  \DLKCLR\    <= \47102\    ; -- A22/1 - INOUT V.
  \RDOUT/\    <= \47105\    ; -- A22/1 - INOUT V.
  \ADVCTR\    <= \47106\    ; -- A22/1 - INOUT V.
  \1CNT\      <= \47109\    ; -- A22/1 - INOUT V.
  \DKCTR1/\   <= \47115\    ; -- A22/1 - INOUT V.
  \DKCTR1\    <= \47116\    ; -- A22/1 - INOUT V.
  \DKCTR2/\   <= \47123\    ; -- A22/1 - INOUT V.
  \DKCTR2\    <= \47124\    ; -- A22/1 - INOUT V.
  \DKCTR3/\   <= \47131\    ; -- A22/1 - INOUT V.
  \DKCTR3\    <= \47132\    ; -- A22/1 - INOUT V.
  \DKCTR4\    <= \47137\    ; -- A22/1 - INOUT V.
  \DKCTR4/\   <= \47138\    ; -- A22/1 - INOUT V.
  \16CNT\     <= \47139\    ; -- A22/1 - INOUT V.
  \32CNT\     <= \47142\    ; -- A22/1 - INOUT V.
  \DKCTR5\    <= \47143\    ; -- A22/1 - INOUT V.
  \DKCTR5/\   <= \47144\    ; -- A22/1 - INOUT V.
  \WDORDR\    <= \47154\    ; -- A22/1 - INOUT V.
  \CH1307\    <= \47158\    ; -- A22/1 - INOUT V.
  \ORDRBT\    <= \47159\    ; -- A22/1 - INOUT V.
  \F12B/\     <= \47161\    ; -- A22/1 - INOUT V.
  \F14H\      <= \47162\    ; -- A22/1 - INOUT V.
  \WCH13/\    <= \47202\    ; -- A22/1 - INOUT V.
  \CCH13\     <= \47207\    ; -- A22/1 - INOUT V.
  \RCH13/\    <= \47211\    ; -- A22/1 - INOUT V.
  \WCH14/\    <= \47215\    ; -- A22/1 - INOUT V.
  \CCH14\     <= \47220\    ; -- A22/1 - INOUT V.
  \RCH14/\    <= \47224\    ; -- A22/1 - INOUT V.
  \BSYNC/\    <= \47227\    ; -- A22/1 - INOUT V.
  \LOW0/\     <= \47229\    ; -- A22/1 - INOUT V.
  \LOW1/\     <= \47231\    ; -- A22/1 - INOUT V.
  \LOW2/\     <= \47233\    ; -- A22/1 - INOUT V.
  \LOW3/\     <= \47235\    ; -- A22/1 - INOUT V.
  \LOW4/\     <= \47237\    ; -- A22/1 - INOUT V.
  \LOW5/\     <= \47239\    ; -- A22/1 - INOUT V.
  \LOW6/\     <= \47241\    ; -- A22/1 - INOUT V.
  \LOW7/\     <= \47243\    ; -- A22/1 - INOUT V.
  \DATA/\     <= \47253\    ; -- A22/1 - INOUT V.
  \DKDAT/\    <= \47255\    ; -- A22/1 - INOUT V.
  \DKDATA\    <= \47256\    ; -- A22/1 - INOUT V.
  \DKDATB\    <= \47261\    ; -- A22/1 - INOUT V.
  \FS13/\     <= \47262\    ; -- A22/1 - INOUT V.
  \WRD1BP\    <= \47304\    ; -- A22/2 - INOUT V.
  \WRD1B1\    <= \47308\    ; -- A22/2 - INOUT V.
  \WRD2B2\    <= \47404\    ; -- A22/2 - INOUT V.
  \WRD2B3\    <= \47408\    ; -- A22/2 - INOUT V.
  \PIPAFL\    <= \48108\    ; -- A23/1 - INOUT VI.
  \WCH35/\    <= \48120\    ; -- A23/1 - INOUT VI.
  \CCH35\     <= \48124\    ; -- A23/1 - INOUT VI.
  \BOTHX\     <= \48127\    ; -- A23/1 - INOUT VI.
  \NOXM\      <= \48149\    ; -- A23/1 - INOUT VI.
  \NOXP\      <= \48151\    ; -- A23/1 - INOUT VI.
  \MISSX\     <= \48153\    ; -- A23/1 - INOUT VI.
  \PIPXP\     <= \48155\    ; -- A23/1 - INOUT VI.
  \PIPXM\     <= \48156\    ; -- A23/1 - INOUT VI.
  \F18B/\     <= \48157\    ; -- A23/1 - INOUT VI.
  \CH01\      <= \48202\    ; -- A23/1 - INOUT VI.
  \CH02\      <= \48204\    ; -- A23/1 - INOUT VI.
  \CH03\      <= \48206\    ; -- A23/1 - INOUT VI.
  \CH04\      <= \48208\    ; -- A23/1 - INOUT VI.
  \CH05\      <= \48211\    ; -- A23/1 - INOUT VI.
  \CH06\      <= \48213\    ; -- A23/1 - INOUT VI.
  \CH07\      <= \48215\    ; -- A23/1 - INOUT VI.
  \CH08\      <= \48218\    ; -- A23/1 - INOUT VI.
  \WCH34/\    <= \48221\    ; -- A23/1 - INOUT VI.
  \CCH34\     <= \48225\    ; -- A23/1 - INOUT VI.
  \BOTHY\     <= \48228\    ; -- A23/1 - INOUT VI.
  \PIPYP\     <= \48250\    ; -- A23/1 - INOUT VI.
  \PIPYM\     <= \48251\    ; -- A23/1 - INOUT VI.
  \NOYM\      <= \48252\    ; -- A23/1 - INOUT VI.
  \NOYP\      <= \48254\    ; -- A23/1 - INOUT VI.
  \MISSY\     <= \48256\    ; -- A23/1 - INOUT VI.
  \CH1416\    <= \48304\    ; -- A23/2 - INOUT VI.
  \CDUXD\     <= \48305\    ; -- A23/2 - INOUT VI.
  \CDUXDP\    <= \48308\    ; -- A23/2 - INOUT VI.
  \CDUXDM\    <= \48309\    ; -- A23/2 - INOUT VI.
  \CH1414\    <= \48314\    ; -- A23/2 - INOUT VI.
  \CDUYD\     <= \48315\    ; -- A23/2 - INOUT VI.
  \CDUYDP\    <= \48318\    ; -- A23/2 - INOUT VI.
  \CDUYDM\    <= \48319\    ; -- A23/2 - INOUT VI.
  \CH1413\    <= \48323\    ; -- A23/2 - INOUT VI.
  \CDUZD\     <= \48325\    ; -- A23/2 - INOUT VI.
  \CDUZDP\    <= \48326\    ; -- A23/2 - INOUT VI.
  \CDUZDM\    <= \48329\    ; -- A23/2 - INOUT VI.
  \CH1412\    <= \48334\    ; -- A23/2 - INOUT VI.
  \TRUND\     <= \48335\    ; -- A23/2 - INOUT VI.
  \TRNDP\     <= \48336\    ; -- A23/2 - INOUT VI.
  \TRNDM\     <= \48339\    ; -- A23/2 - INOUT VI.
  \CH1411\    <= \48344\    ; -- A23/2 - INOUT VI.
  \SHAFTD\    <= \48345\    ; -- A23/2 - INOUT VI.
  \SHFTDP\    <= \48348\    ; -- A23/2 - INOUT VI.
  \SHFTDM\    <= \48349\    ; -- A23/2 - INOUT VI.
  \POUT/\     <= \48351\    ; -- A23/2 - INOUT VI.
  \MOUT/\     <= \48353\    ; -- A23/2 - INOUT VI.
  \ZOUT/\     <= \48355\    ; -- A23/2 - INOUT VI.
  \T7PHS4/\   <= \48358\    ; -- A23/2 - INOUT VI.
  \T7PHS4\    <= \48359\    ; -- A23/2 - INOUT VI.
  \E5\        <= \48403\    ; -- A23/2 - INOUT VI.
  \CH0705\    <= \48404\    ; -- A23/2 - INOUT VI.
  \E6\        <= \48407\    ; -- A23/2 - INOUT VI.
  \CH0706\    <= \48408\    ; -- A23/2 - INOUT VI.
  \E7/\       <= \48410\    ; -- A23/2 - INOUT VI.
  \CH0707\    <= \48412\    ; -- A23/2 - INOUT VI.
  \CCH07\     <= \48413\    ; -- A23/2 - INOUT VI.
  \WCH07/\    <= \48415\    ; -- A23/2 - INOUT VI.
  \RCH07/\    <= \48417\    ; -- A23/2 - INOUT VI.
  \CH1108\    <= \48421\    ; -- A23/2 - INOUT VI.
  \OT1108\    <= \48422\    ; -- A23/2 - INOUT VI.
  \CH1113\    <= \48426\    ; -- A23/2 - INOUT VI.
  \OT1113\    <= \48427\    ; -- A23/2 - INOUT VI.
  \CH1114\    <= \48431\    ; -- A23/2 - INOUT VI.
  \OT1114\    <= \48432\    ; -- A23/2 - INOUT VI.
  \CH1116\    <= \48436\    ; -- A23/2 - INOUT VI.
  \OT1116\    <= \48437\    ; -- A23/2 - INOUT VI.
  \CH09\      <= \48440\    ; -- A23/2 - INOUT VI.
  \CH1216\    <= \48444\    ; -- A23/2 - INOUT VI.
  \ISSTDC\    <= \48445\    ; -- A23/2 - INOUT VI.
  \T6ON/\     <= \48447\    ; -- A23/2 - INOUT VI.
  \CH1316\    <= \48449\    ; -- A23/2 - INOUT VI.
  \CH1310\    <= \48453\    ; -- A23/2 - INOUT VI.
  \ALTEST\    <= \48454\    ; -- A23/2 - INOUT VI.
  \CH10\      <= \48458\    ; -- A23/2 - INOUT VI.
  \OVNHRP\    <= \49109\    ; -- A24/1 - INOUT VII.
  \WATCHP\    <= \49114\    ; -- A24/1 - INOUT VII.
  \WATCH/\    <= \49116\    ; -- A24/1 - INOUT VII.
  \WATCH\     <= \49117\    ; -- A24/1 - INOUT VII.
  \HIGH0/\    <= \49121\    ; -- A24/1 - INOUT VII.
  \HIGH1/\    <= \49124\    ; -- A24/1 - INOUT VII.
  \HIGH2/\    <= \49127\    ; -- A24/1 - INOUT VII.
  \HIGH3/\    <= \49130\    ; -- A24/1 - INOUT VII.
  \RCHG/\     <= \49133\    ; -- A24/1 - INOUT VII.
  \WCHG/\     <= \49137\    ; -- A24/1 - INOUT VII.
  \CCHG/\     <= \49141\    ; -- A24/1 - INOUT VII.
  \CHWL01/\   <= \49143\    ; -- A24/1 - INOUT VII.
  \CHWL02/\   <= \49145\    ; -- A24/1 - INOUT VII.
  \CHWL03/\   <= \49147\    ; -- A24/1 - INOUT VII.
  \CHWL04/\   <= \49149\    ; -- A24/1 - INOUT VII.
  \CHWL05/\   <= \49151\    ; -- A24/1 - INOUT VII.
  \CHWL06/\   <= \49153\    ; -- A24/1 - INOUT VII.
  \CHWL07/\   <= \49155\    ; -- A24/1 - INOUT VII.
  \CHWL08/\   <= \49157\    ; -- A24/1 - INOUT VII.
  \CHWL09/\   <= \49159\    ; -- A24/1 - INOUT VII.
  \PIPPLS/\   <= \49203\    ; -- A24/1 - INOUT VII.
  \PIPASW\    <= \49204\    ; -- A24/1 - INOUT VII.
  \FS05/\     <= \49205\    ; -- A24/1 - INOUT VII.
  \PIPDAT\    <= \49206\    ; -- A24/1 - INOUT VII.
  \PIPINT\    <= \49208\    ; -- A24/1 - INOUT VII.
  \800SET\    <= \49209\    ; -- A24/1 - INOUT VII.
  \800RST\    <= \49210\    ; -- A24/1 - INOUT VII.
  \3200A\     <= \49211\    ; -- A24/1 - INOUT VII.
  \3200B\     <= \49212\    ; -- A24/1 - INOUT VII.
  \3200C\     <= \49213\    ; -- A24/1 - INOUT VII.
  \3200D\     <= \49215\    ; -- A24/1 - INOUT VII.
  \12KPPS\    <= \49217\    ; -- A24/1 - INOUT VII.
  \RRRST\     <= \49218\    ; -- A24/1 - INOUT VII.
  \LRRST\     <= \49219\    ; -- A24/1 - INOUT VII.
  \25KPPS\    <= \49220\    ; -- A24/1 - INOUT VII.
  \CDUCLK\    <= \49223\    ; -- A24/1 - INOUT VII.
  \SB0/\      <= \49224\    ; -- A24/1 - INOUT VII.
  \SB1/\      <= \49226\    ; -- A24/1 - INOUT VII.
  \SB2/\      <= \49228\    ; -- A24/1 - INOUT VII.
  \F05A/\     <= \49230\    ; -- A24/1 - INOUT VII.
  \F05B/\     <= \49232\    ; -- A24/1 - INOUT VII.
  \F07B/\     <= \49234\    ; -- A24/1 - INOUT VII.
  \CHWL10/\   <= \49235\    ; -- A24/1 - INOUT VII.
  \NISQ\      <= \49237\    ; -- A24/1 - INOUT VII.
  \RCHAT/\    <= \49241\    ; -- A24/1 - INOUT VII.
  \RCHBT/\    <= \49245\    ; -- A24/1 - INOUT VII.
  \ELSNCN\    <= \49249\    ; -- A24/1 - INOUT VII.
  \ELSNCM\    <= \49250\    ; -- A24/1 - INOUT VII.
  \OT1110\    <= \49252\    ; -- A24/1 - INOUT VII.
  \OT1111\    <= \49253\    ; -- A24/1 - INOUT VII.
  \OT1112\    <= \49254\    ; -- A24/1 - INOUT VII.
  \NOZM\      <= \49303\    ; -- A24/2 - INOUT VII.
  \NOZP\      <= \49305\    ; -- A24/2 - INOUT VII.
  \MISSZ\     <= \49307\    ; -- A24/2 - INOUT VII.
  \BOTHZ\     <= \49309\    ; -- A24/2 - INOUT VII.
  \PIPZP\     <= \49329\    ; -- A24/2 - INOUT VII.
  \PIPZM\     <= \49330\    ; -- A24/2 - INOUT VII.
  \CNTRSB/\   <= \49331\    ; -- A24/2 - INOUT VII.
  \RSCT/\     <= \49332\    ; -- A24/2 - INOUT VII.
  \US2SG\     <= \49336\    ; -- A24/2 - INOUT VII.
  \U2BBKG/\   <= \49337\    ; -- A24/2 - INOUT VII.
  \GTSET\     <= \49343\    ; -- A24/2 - INOUT VII.
  \GTSET/\    <= \49344\    ; -- A24/2 - INOUT VII.
  \GTRST\     <= \49345\    ; -- A24/2 - INOUT VII.
  \GTONE\     <= \49346\    ; -- A24/2 - INOUT VII.
  \FS09/\     <= \49348\    ; -- A24/2 - INOUT VII.
  \F09D\      <= \49352\    ; -- A24/2 - INOUT VII.
  \F09A/\     <= \49353\    ; -- A24/2 - INOUT VII.
  \CI\        <= \49354\    ; -- A24/2 - INOUT VII.
  \F07D/\     <= \49357\    ; -- A24/2 - INOUT VII.
  \F07C/\     <= \49358\    ; -- A24/2 - INOUT VII.
  \F7CSB1/\   <= \49360\    ; -- A24/2 - INOUT VII.
  \FLASH\     <= \49409\    ; -- A24/2 - INOUT VII.
  \FLASH/\    <= \49410\    ; -- A24/2 - INOUT VII.
  \ONE\       <= \49411\    ; -- A24/2 - INOUT VII.
  \CDUSTB/\   <= \49413\    ; -- A24/2 - INOUT VII.
  \PHS3/\     <= \49414\    ; -- A24/2 - INOUT VII.
  \F04B/\     <= \49418\    ; -- A24/2 - INOUT VII.
  \IC11/\     <= \49419\    ; -- A24/2 - INOUT VII.
  \F05D\      <= \49420\    ; -- A24/2 - INOUT VII.
  \CHWL11/\   <= \49425\    ; -- A24/2 - INOUT VII.
  \CHWL12/\   <= \49427\    ; -- A24/2 - INOUT VII.
  \CHWL13/\   <= \49429\    ; -- A24/2 - INOUT VII.
  \CHWL14/\   <= \49431\    ; -- A24/2 - INOUT VII.
  \CHWL16/\   <= \49433\    ; -- A24/2 - INOUT VII.
  \MDT01\     <= \21A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT02\     <= \22A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT03\     <= \23A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT04\     <= \24A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT05\     <= \25A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT06\     <= \26A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT07\     <= \27A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT08\     <= \28A\      ; -- CH77/1 - RESTART MONITOR.
  \MDT09\     <= \29A\      ; -- CH77/1 - RESTART MONITOR.
  \DERHI\     <= \PULLD01\  ; -- CH77/1 - RESTART MONITOR.
  \DERLO\     <= \PULLD02\  ; -- CH77/1 - RESTART MONITOR.
  \MDT10\     <= \PULLD03\  ; -- CH77/1 - RESTART MONITOR.
  \MDT11\     <= \PULLD04\  ; -- CH77/1 - RESTART MONITOR.
  \MDT12\     <= \PULLD05\  ; -- CH77/1 - RESTART MONITOR.
  \MDT13\     <= \PULLD06\  ; -- CH77/1 - RESTART MONITOR.
  \MDT14\     <= \PULLD07\  ; -- CH77/1 - RESTART MONITOR.
  \MDT15\     <= \PULLD08\  ; -- CH77/1 - RESTART MONITOR.
  \MDT16\     <= \PULLD09\  ; -- CH77/1 - RESTART MONITOR.
  \MNHSBF\    <= \PULLD10\  ; -- CH77/1 - RESTART MONITOR.
  \MNHNC\     <= \PULLD11\  ; -- CH77/1 - RESTART MONITOR.
  \MNHRPT\    <= \PULLD12\  ; -- CH77/1 - RESTART MONITOR.
  \MTCSAI\    <= \PULLD13\  ; -- CH77/1 - RESTART MONITOR.
  \MSTRT\     <= \PULLD14\  ; -- CH77/1 - RESTART MONITOR.
  \MSTP\      <= \PULLD15\  ; -- CH77/1 - RESTART MONITOR.
  \MSBSTP\    <= \PULLD16\  ; -- CH77/1 - RESTART MONITOR.
  \MRDCH\     <= \PULLD17\  ; -- CH77/1 - RESTART MONITOR.
  \MLDCH\     <= \PULLD18\  ; -- CH77/1 - RESTART MONITOR.
  \MONPAR\    <= \PULLD19\  ; -- CH77/1 - RESTART MONITOR.
  \MONWBK\    <= \PULLD20\  ; -- CH77/1 - RESTART MONITOR.
  \MLOAD\     <= \PULLD21\  ; -- CH77/1 - RESTART MONITOR.
  \MREAD\     <= \PULLD22\  ; -- CH77/1 - RESTART MONITOR.
  \NHALGA\    <= \PULLD23\  ; -- CH77/1 - RESTART MONITOR.
  \DOSCAL\    <= \PULLD24\  ; -- CH77/1 - RESTART MONITOR.
  \DBLTST\    <= \PULLD25\  ; -- CH77/1 - RESTART MONITOR.
  \MAMU\      <= \PULLD26\  ; -- CH77/1 - RESTART MONITOR.
  \MWL01\     <= \PULLU01\  ; -- CH77/1 - RESTART MONITOR.
  \MWL02\     <= \PULLU02\  ; -- CH77/1 - RESTART MONITOR.
  \MWL03\     <= \PULLU03\  ; -- CH77/1 - RESTART MONITOR.
  \MWL04\     <= \PULLU04\  ; -- CH77/1 - RESTART MONITOR.
  \MWL05\     <= \PULLU05\  ; -- CH77/1 - RESTART MONITOR.
  \MWL06\     <= \PULLU06\  ; -- CH77/1 - RESTART MONITOR.
  \MT01\      <= \PULLU07\  ; -- CH77/1 - RESTART MONITOR.
  \MWSG\      <= \PULLU08\  ; -- CH77/1 - RESTART MONITOR.
  \MT12\      <= \PULLU09\  ; -- CH77/1 - RESTART MONITOR.
  \MWCH\      <= \PULLU10\  ; -- CH77/1 - RESTART MONITOR.
  \MRCH\      <= \PULLU11\  ; -- CH77/1 - RESTART MONITOR.
  \MPAL/\     <= \PULLU12\  ; -- CH77/1 - RESTART MONITOR.
  \MT05\      <= \PULLU13\  ; -- CH77/1 - RESTART MONITOR.
  \MTCAL/\    <= \PULLU14\  ; -- CH77/1 - RESTART MONITOR.
  \MRPTAL/\   <= \PULLU15\  ; -- CH77/1 - RESTART MONITOR.
  \MWATCH/\   <= \PULLU16\  ; -- CH77/1 - RESTART MONITOR.
  \MVFAIL/\   <= \PULLU17\  ; -- CH77/1 - RESTART MONITOR.
  \MCTRAL/\   <= \PULLU18\  ; -- CH77/1 - RESTART MONITOR.
  \MSCAFL/\   <= \PULLU19\  ; -- CH77/1 - RESTART MONITOR.
  \MSCDBL/\   <= \PULLU20\  ; -- CH77/1 - RESTART MONITOR.
  \GEM01\     <= \PULLU21\  ; -- CH77/1 - RESTART MONITOR.
  \GEM02\     <= \PULLU22\  ; -- CH77/1 - RESTART MONITOR.
  \GEM03\     <= \PULLU23\  ; -- CH77/1 - RESTART MONITOR.
  \GEM04\     <= \PULLU24\  ; -- CH77/1 - RESTART MONITOR.
  \GEM05\     <= \PULLU25\  ; -- CH77/1 - RESTART MONITOR.
  \GEM06\     <= \PULLU26\  ; -- CH77/1 - RESTART MONITOR.
  \GEM07\     <= \PULLU27\  ; -- CH77/1 - RESTART MONITOR.
  \GEM08\     <= \PULLU28\  ; -- CH77/1 - RESTART MONITOR.
  \GEM09\     <= \PULLU29\  ; -- CH77/1 - RESTART MONITOR.
  \GEM10\     <= \PULLU30\  ; -- CH77/1 - RESTART MONITOR.
  \GEM11\     <= \PULLU31\  ; -- CH77/1 - RESTART MONITOR.
  \GEM12\     <= \PULLU32\  ; -- CH77/1 - RESTART MONITOR.
  \GEM13\     <= \PULLU33\  ; -- CH77/1 - RESTART MONITOR.
  \GEM14\     <= \PULLU34\  ; -- CH77/1 - RESTART MONITOR.
  \GEM16\     <= \PULLU35\  ; -- CH77/1 - RESTART MONITOR.
  \GEMP\      <= \PULLU36\  ; -- CH77/1 - RESTART MONITOR.
  \SBE\       <= \PULLU37\  ; -- CH77/1 - RESTART MONITOR.
  \SBF\       <= \PULLU38\  ; -- CH77/1 - RESTART MONITOR.
  \ZID\       <= \PULLU39\  ; -- CH77/1 - RESTART MONITOR.
  \REX\       <= \PULLU40\  ; -- CH77/1 - RESTART MONITOR.
  \REY\       <= \PULLU41\  ; -- CH77/1 - RESTART MONITOR.
  \WEX\       <= \PULLU42\  ; -- CH77/1 - RESTART MONITOR.
  \WEY\       <= \PULLU43\  ; -- CH77/1 - RESTART MONITOR.
  \CLROPE\    <= \PULLU44\  ; -- CH77/1 - RESTART MONITOR.
  \FILTIN\    <= \PULLU45\  ; -- CH77/1 - RESTART MONITOR.
  \HIMOD\     <= \PULLU46\  ; -- CH77/1 - RESTART MONITOR.
  \IHENV\     <= \PULLU47\  ; -- CH77/1 - RESTART MONITOR.
  \IL01\      <= \PULLU48\  ; -- CH77/1 - RESTART MONITOR.
  \IL01/\     <= \PULLU49\  ; -- CH77/1 - RESTART MONITOR.
  \IL02\      <= \PULLU50\  ; -- CH77/1 - RESTART MONITOR.
  \IL02/\     <= \PULLU51\  ; -- CH77/1 - RESTART MONITOR.
  \IL03\      <= \PULLU52\  ; -- CH77/1 - RESTART MONITOR.
  \IL03/\     <= \PULLU53\  ; -- CH77/1 - RESTART MONITOR.
  \IL04\      <= \PULLU54\  ; -- CH77/1 - RESTART MONITOR.
  \IL04/\     <= \PULLU55\  ; -- CH77/1 - RESTART MONITOR.
  \IL05\      <= \PULLU56\  ; -- CH77/1 - RESTART MONITOR.
  \IL05/\     <= \PULLU57\  ; -- CH77/1 - RESTART MONITOR.
  \IL06\      <= \PULLU58\  ; -- CH77/1 - RESTART MONITOR.
  \IL06/\     <= \PULLU59\  ; -- CH77/1 - RESTART MONITOR.
  \IL07\      <= \PULLU60\  ; -- CH77/1 - RESTART MONITOR.
  \IL07/\     <= \PULLU61\  ; -- CH77/1 - RESTART MONITOR.
  \ILP\       <= \PULLU62\  ; -- CH77/1 - RESTART MONITOR.
  \ILP/\      <= \PULLU63\  ; -- CH77/1 - RESTART MONITOR.
  \LOMOD\     <= \PULLU64\  ; -- CH77/1 - RESTART MONITOR.
  \MBR1\      <= \PULLU65\  ; -- CH77/1 - RESTART MONITOR.
  \MBR2\      <= \PULLU66\  ; -- CH77/1 - RESTART MONITOR.
  \MGOJAM\    <= \PULLU67\  ; -- CH77/1 - RESTART MONITOR.
  \MGP/\      <= \PULLU68\  ; -- CH77/1 - RESTART MONITOR.
  \MIIP\      <= \PULLU69\  ; -- CH77/1 - RESTART MONITOR.
  \MINHL\     <= \PULLU70\  ; -- CH77/1 - RESTART MONITOR.
  \MINKL\     <= \PULLU71\  ; -- CH77/1 - RESTART MONITOR.
  \MNISQ\     <= \PULLU72\  ; -- CH77/1 - RESTART MONITOR.
  \MON800\    <= \PULLU73\  ; -- CH77/1 - RESTART MONITOR.
  \MONWT\     <= \PULLU74\  ; -- CH77/1 - RESTART MONITOR.
  \MOSCAL/\   <= \PULLU75\  ; -- CH77/1 - RESTART MONITOR.
  \MPIPAL/\   <= \PULLU76\  ; -- CH77/1 - RESTART MONITOR.
  \MRAG\      <= \PULLU77\  ; -- CH77/1 - RESTART MONITOR.
  \MREQIN\    <= \PULLU78\  ; -- CH77/1 - RESTART MONITOR.
  \MRGG\      <= \PULLU79\  ; -- CH77/1 - RESTART MONITOR.
  \MRLG\      <= \PULLU80\  ; -- CH77/1 - RESTART MONITOR.
  \MRSC\      <= \PULLU81\  ; -- CH77/1 - RESTART MONITOR.
  \MRULOG\    <= \PULLU82\  ; -- CH77/1 - RESTART MONITOR.
  \MSP\       <= \PULLU83\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ10\     <= \PULLU84\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ11\     <= \PULLU85\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ12\     <= \PULLU86\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ13\     <= \PULLU87\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ14\     <= \PULLU88\  ; -- CH77/1 - RESTART MONITOR.
  \MSQ16\     <= \PULLU89\  ; -- CH77/1 - RESTART MONITOR.
  \MSQEXT\    <= \PULLU90\  ; -- CH77/1 - RESTART MONITOR.
  \MST1\      <= \PULLU91\  ; -- CH77/1 - RESTART MONITOR.
  \MST2\      <= \PULLU92\  ; -- CH77/1 - RESTART MONITOR.
  \MST3\      <= \PULLU93\  ; -- CH77/1 - RESTART MONITOR.
  \MSTPIT/\   <= \PULLU94\  ; -- CH77/1 - RESTART MONITOR.
  \MT02\      <= \PULLU95\  ; -- CH77/1 - RESTART MONITOR.
  \MT03\      <= \PULLU96\  ; -- CH77/1 - RESTART MONITOR.
  \MT04\      <= \PULLU97\  ; -- CH77/1 - RESTART MONITOR.
  \MT06\      <= \PULLU98\  ; -- CH77/1 - RESTART MONITOR.
  \MT07\      <= \PULLU99\  ; -- CH77/1 - RESTART MONITOR.
  \MT08\      <= \PULLU100\ ; -- CH77/1 - RESTART MONITOR.
  \MT09\      <= \PULLU101\ ; -- CH77/1 - RESTART MONITOR.
  \MT10\      <= \PULLU102\ ; -- CH77/1 - RESTART MONITOR.
  \MT11\      <= \PULLU103\ ; -- CH77/1 - RESTART MONITOR.
  \MTCSA/\    <= \PULLU104\ ; -- CH77/1 - RESTART MONITOR.
  \MWAG\      <= \PULLU105\ ; -- CH77/1 - RESTART MONITOR.
  \MWARNF/\   <= \PULLU106\ ; -- CH77/1 - RESTART MONITOR.
  \MWBBEG\    <= \PULLU107\ ; -- CH77/1 - RESTART MONITOR.
  \MWBG\      <= \PULLU108\ ; -- CH77/1 - RESTART MONITOR.
  \MWEBG\     <= \PULLU109\ ; -- CH77/1 - RESTART MONITOR.
  \MWFBG\     <= \PULLU110\ ; -- CH77/1 - RESTART MONITOR.
  \MWG\       <= \PULLU111\ ; -- CH77/1 - RESTART MONITOR.
  \MWL07\     <= \PULLU112\ ; -- CH77/1 - RESTART MONITOR.
  \MWL08\     <= \PULLU113\ ; -- CH77/1 - RESTART MONITOR.
  \MWL09\     <= \PULLU114\ ; -- CH77/1 - RESTART MONITOR.
  \MWL10\     <= \PULLU115\ ; -- CH77/1 - RESTART MONITOR.
  \MWL11\     <= \PULLU116\ ; -- CH77/1 - RESTART MONITOR.
  \MWL12\     <= \PULLU117\ ; -- CH77/1 - RESTART MONITOR.
  \MWL13\     <= \PULLU118\ ; -- CH77/1 - RESTART MONITOR.
  \MWL14\     <= \PULLU119\ ; -- CH77/1 - RESTART MONITOR.
  \MWL15\     <= \PULLU120\ ; -- CH77/1 - RESTART MONITOR.
  \MWL16\     <= \PULLU121\ ; -- CH77/1 - RESTART MONITOR.
  \MWLG\      <= \PULLU122\ ; -- CH77/1 - RESTART MONITOR.
  \MWQG\      <= \PULLU123\ ; -- CH77/1 - RESTART MONITOR.
  \MWYG\      <= \PULLU124\ ; -- CH77/1 - RESTART MONITOR.
  \MWZG\      <= \PULLU125\ ; -- CH77/1 - RESTART MONITOR.
  \OUTCOM\    <= \PULLU126\ ; -- CH77/1 - RESTART MONITOR.
  \Q2A\       <= \PULLU127\ ; -- CH77/1 - RESTART MONITOR.
  \RESETA\    <= \PULLU128\ ; -- CH77/1 - RESTART MONITOR.
  \RESETB\    <= \PULLU129\ ; -- CH77/1 - RESTART MONITOR.
  \RESETC\    <= \PULLU130\ ; -- CH77/1 - RESTART MONITOR.
  \RESETD\    <= \PULLU131\ ; -- CH77/1 - RESTART MONITOR.
  \ROPER\     <= \PULLU132\ ; -- CH77/1 - RESTART MONITOR.
  \ROPES\     <= \PULLU133\ ; -- CH77/1 - RESTART MONITOR.
  \ROPET\     <= \PULLU134\ ; -- CH77/1 - RESTART MONITOR.
  \RSTKX/\    <= \PULLU135\ ; -- CH77/1 - RESTART MONITOR.
  \RSTKY/\    <= \PULLU136\ ; -- CH77/1 - RESTART MONITOR.
  \SBYREL/\   <= \PULLU137\ ; -- CH77/1 - RESTART MONITOR.
  \SCAS10\    <= \PULLU138\ ; -- CH77/1 - RESTART MONITOR.
  \SCAS17\    <= \PULLU139\ ; -- CH77/1 - RESTART MONITOR.
  \SETAB\     <= \PULLU140\ ; -- CH77/1 - RESTART MONITOR.
  \SETCD\     <= \PULLU141\ ; -- CH77/1 - RESTART MONITOR.
  \SETEK\     <= \PULLU142\ ; -- CH77/1 - RESTART MONITOR.
  \STR14\     <= \PULLU143\ ; -- CH77/1 - RESTART MONITOR.
  \STR19\     <= \PULLU144\ ; -- CH77/1 - RESTART MONITOR.
  \STR210\    <= \PULLU145\ ; -- CH77/1 - RESTART MONITOR.
  \STR311\    <= \PULLU146\ ; -- CH77/1 - RESTART MONITOR.
  \STR412\    <= \PULLU147\ ; -- CH77/1 - RESTART MONITOR.
  \STR58\     <= \PULLU148\ ; -- CH77/1 - RESTART MONITOR.
  \STR912\    <= \PULLU149\ ; -- CH77/1 - RESTART MONITOR.
  \XB0E\      <= \PULLU151\ ; -- CH77/1 - RESTART MONITOR.
  \XB1E\      <= \PULLU152\ ; -- CH77/1 - RESTART MONITOR.
  \XB2E\      <= \PULLU153\ ; -- CH77/1 - RESTART MONITOR.
  \XB3E\      <= \PULLU154\ ; -- CH77/1 - RESTART MONITOR.
  \XB4E\      <= \PULLU155\ ; -- CH77/1 - RESTART MONITOR.
  \XB5E\      <= \PULLU156\ ; -- CH77/1 - RESTART MONITOR.
  \XB6E\      <= \PULLU157\ ; -- CH77/1 - RESTART MONITOR.
  \XB7E\      <= \PULLU158\ ; -- CH77/1 - RESTART MONITOR.
  \XT0E\      <= \PULLU159\ ; -- CH77/1 - RESTART MONITOR.
  \XT1E\      <= \PULLU160\ ; -- CH77/1 - RESTART MONITOR.
  \XT2E\      <= \PULLU161\ ; -- CH77/1 - RESTART MONITOR.
  \XT3E\      <= \PULLU162\ ; -- CH77/1 - RESTART MONITOR.
  \XT4E\      <= \PULLU163\ ; -- CH77/1 - RESTART MONITOR.
  \XT5E\      <= \PULLU164\ ; -- CH77/1 - RESTART MONITOR.
  \XT6E\      <= \PULLU165\ ; -- CH77/1 - RESTART MONITOR.
  \XT7E\      <= \PULLU166\ ; -- CH77/1 - RESTART MONITOR.
  \YB0E\      <= \PULLU167\ ; -- CH77/1 - RESTART MONITOR.
  \YB1E\      <= \PULLU168\ ; -- CH77/1 - RESTART MONITOR.
  \YB2E\      <= \PULLU169\ ; -- CH77/1 - RESTART MONITOR.
  \YB3E\      <= \PULLU170\ ; -- CH77/1 - RESTART MONITOR.
  \YT0E\      <= \PULLU171\ ; -- CH77/1 - RESTART MONITOR.
  \YT1E\      <= \PULLU172\ ; -- CH77/1 - RESTART MONITOR.
  \YT2E\      <= \PULLU173\ ; -- CH77/1 - RESTART MONITOR.
  \YT3E\      <= \PULLU174\ ; -- CH77/1 - RESTART MONITOR.
  \YT4E\      <= \PULLU175\ ; -- CH77/1 - RESTART MONITOR.
  \YT5E\      <= \PULLU176\ ; -- CH77/1 - RESTART MONITOR.
  \YT6E\      <= \PULLU177\ ; -- CH77/1 - RESTART MONITOR.
  \YT7E\      <= \PULLU178\ ; -- CH77/1 - RESTART MONITOR.

  -- ****************************
  -- ***                      ***
  -- ***  OUTPUT assignment.  ***
  -- ***                      ***
  -- ****************************

  ECADR(11)  <= \EAD11\; -- MSB of Erasable Address.
  ECADR(10)  <= \EAD10\;
  ECADR( 9)  <= \EAD09\;
  ECADR( 8)  <= \S08\;
  ECADR( 7)  <= \S07\;
  ECADR( 6)  <= \S06\;
  ECADR( 5)  <= \S05\;
  ECADR( 4)  <= \S04\;
  ECADR( 3)  <= \S03\;
  ECADR( 2)  <= \S02\;
  ECADR( 1)  <= \S01\;   -- LSB of Erasable Address.

  FCADR(16)  <= \F16\;   -- MSB of Fixed Address.
  FCADR(15)  <= \F15\;
  FCADR(14)  <= \F14\;
  FCADR(13)  <= \F13\;
  FCADR(12)  <= \F12\;
  FCADR(11)  <= \F11\;
  FCADR(10)  <= \S10\;
  FCADR( 9)  <= \S09\;
  FCADR( 8)  <= \S08\;
  FCADR( 7)  <= \S07\;
  FCADR( 6)  <= \S06\;
  FCADR( 5)  <= \S05\;
  FCADR( 4)  <= \S04\;
  FCADR( 3)  <= \S03\;
  FCADR( 2)  <= \S02\;
  FCADR( 1)  <= \S01\;   -- LSB of Fixed Address.

  GEMXX(15)  <= \GEM16\; -- MSB of data from G regsiter to Erasable memory.
  GEMXX(14)  <= \GEM14\;
  GEMXX(13)  <= \GEM13\;
  GEMXX(12)  <= \GEM12\;
  GEMXX(11)  <= \GEM11\;
  GEMXX(10)  <= \GEM10\;
  GEMXX( 9)  <= \GEM09\;
  GEMXX( 8)  <= \GEM08\;
  GEMXX( 7)  <= \GEM07\;
  GEMXX( 6)  <= \GEM06\;
  GEMXX( 5)  <= \GEM05\;
  GEMXX( 4)  <= \GEM04\;
  GEMXX( 3)  <= \GEM03\;
  GEMXX( 2)  <= \GEM02\;
  GEMXX( 1)  <= \GEM01\; -- LSB of data from G register to Erasable memory.
  GEMXX( 0)  <= \GEMP\;  -- Parity of data to Erasable memory.

  EWRITE     <= \ZID\;   -- Erasable write signal.
  EREAD      <= \SBE\;   -- Erasable read  signal.
  ESTART     <= \SETEK\; -- Start of erasable cycle.
  FREAD      <= \SBF\;   -- Fixed read signal.

  OUTPUTS.\3200A\      <= \3200A\;
  OUTPUTS.\CDUXDP\     <= \CDUXDP\;
  OUTPUTS.\3200B\      <= \3200B\;
  OUTPUTS.\CDUXDM\     <= \CDUXDM\;
  OUTPUTS.\3200C\      <= \3200C\;
  OUTPUTS.\CDUYDP\     <= \CDUYDP\;
  OUTPUTS.\3200D\      <= \3200D\;
  OUTPUTS.\CDUYDM\     <= \CDUYDM\;
  OUTPUTS.\25KPPS\     <= \25KPPS\;
  OUTPUTS.\CDUCLK\     <= \CDUCLK\;
  OUTPUTS.\12KPPS\     <= \12KPPS\;
  OUTPUTS.\PIPINT\     <= \PIPINT\;
  OUTPUTS.\800SET\     <= \800SET\;
  OUTPUTS.\PIPASW\     <= \PIPASW\;
  OUTPUTS.\800RST\     <= \800RST\;
  OUTPUTS.\PIPDAT\     <= \PIPDAT\;
  OUTPUTS.\GYENAB\     <= \GYENAB\;
  OUTPUTS.\CLK\        <= \CLK\;
  OUTPUTS.\CDUZDP\     <= \CDUZDP\;
  OUTPUTS.\RRRST\      <= \RRRST\;
  OUTPUTS.\CDUZDM\     <= \CDUZDM\;
  OUTPUTS.\LRRST\      <= \LRRST\;
  OUTPUTS.\OT1114\     <= \OT1114\;
  OUTPUTS.\RC-X+P\     <= \RC-X+P\;
  OUTPUTS.\OT1113\     <= \OT1113\;
  OUTPUTS.\RC+X-Y\     <= \RC+X-Y\;
  OUTPUTS.\OT1112\     <= \OT1112\;
  OUTPUTS.\RC+X+Y\     <= \RC+X+Y\;
  OUTPUTS.\OT1111\     <= \OT1111\;
  OUTPUTS.\RC+X-P\     <= \RC+X-P\;
  OUTPUTS.\OT1110\     <= \OT1110\;
  OUTPUTS.\RC+X+P\     <= \RC+X+P\;
  OUTPUTS.\OT1108\     <= \OT1108\;
  OUTPUTS.\TMPCAU\     <= \TMPCAU\;
  OUTPUTS.\OPEROR\     <= \OPEROR\;
  OUTPUTS.\ISSTDC\     <= \ISSTDC\;
  OUTPUTS.\ELSNCM\     <= \ELSNCM\;
  OUTPUTS.\OT1116\     <= \OT1116\;
  OUTPUTS.\VNFLSH\     <= \VNFLSH\;
  OUTPUTS.\ENERIM\     <= \ENERIM\;
  OUTPUTS.\CGCWAR\     <= \CGCWAR\;
  OUTPUTS.\ZIMCDU\     <= \ZIMCDU\;
  OUTPUTS.\KYRLS\      <= \KYRLS\;
  OUTPUTS.\COARSE\     <= \COARSE\;
  OUTPUTS.\UPLACT\     <= \UPLACT\;
  OUTPUTS.\ENEROP\     <= \ENEROP\;
  OUTPUTS.\S4BOFF\     <= \S4BOFF\;
  OUTPUTS.\ZEROPT\     <= \ZEROPT\;
  OUTPUTS.\S4BSEQ\     <= \S4BSEQ\;
  OUTPUTS.\MROLGT\     <= \MROLGT\;
  OUTPUTS.\RESTRT\     <= \RESTRT\;
  OUTPUTS.\ZOPCDU\     <= \ZOPCDU\;
  OUTPUTS.\SBYLIT\     <= \SBYLIT\;
  OUTPUTS.\ALTSNC\     <= \ALTSNC\;
  OUTPUTS.\COMACT\     <= \COMACT\;
  OUTPUTS.\OT1207/\    <= \OT1207/\;
  OUTPUTS.\ISSWAR\     <= \ISSWAR\;
  OUTPUTS.\OT1207\     <= \OT1207\;
  OUTPUTS.\RYWD16\     <= \RYWD16\;
  OUTPUTS.\S4BTAK\     <= \S4BTAK\;
  OUTPUTS.\RYWD14\     <= \RYWD14\;
  OUTPUTS.\DISDAC\     <= \DISDAC\;
  OUTPUTS.\RYWD13\     <= \RYWD13\;
  OUTPUTS.\STARON\     <= \STARON\;
  OUTPUTS.\RYWD12\     <= \RYWD12\;
  OUTPUTS.\TVCNAB\     <= \TVCNAB\;
  OUTPUTS.\RLYB11\     <= \RLYB11\;
  OUTPUTS.\RC-Z-R\     <= \RC-Z-R\;
  OUTPUTS.\RLYB10\     <= \RLYB10\;
  OUTPUTS.\RC-Z+R\     <= \RC-Z+R\;
  OUTPUTS.\RLYB09\     <= \RLYB09\;
  OUTPUTS.\RC+Z-R\     <= \RC+Z-R\;
  OUTPUTS.\RLYB08\     <= \RLYB08\;
  OUTPUTS.\RC+Z+R\     <= \RC+Z+R\;
  OUTPUTS.\RLYB07\     <= \RLYB07\;
  OUTPUTS.\RC-Y-R\     <= \RC-Y-R\;
  OUTPUTS.\RLYB06\     <= \RLYB06\;
  OUTPUTS.\RC-Y+R\     <= \RC-Y+R\;
  OUTPUTS.\RLYB05\     <= \RLYB05\;
  OUTPUTS.\RC+Y-R\     <= \RC+Y-R\;
  OUTPUTS.\RLYB04\     <= \RLYB04\;
  OUTPUTS.\RC+Y+R\     <= \RC+Y+R\;
  OUTPUTS.\RLYB03\     <= \RLYB03\;
  OUTPUTS.\RC-X-Y\     <= \RC-X-Y\;
  OUTPUTS.\RLYB02\     <= \RLYB02\;
  OUTPUTS.\RC-X+Y\     <= \RC-X+Y\;
  OUTPUTS.\RLYB01\     <= \RLYB01\;
  OUTPUTS.\RC-X-P\     <= \RC-X-P\;
  OUTPUTS.\ELSNCN\     <= \ELSNCN\;
  OUTPUTS.\THRST+\     <= \THRST+\;
  OUTPUTS.\LRRANG\     <= \LRRANG\;
  OUTPUTS.\SHFTDP\     <= \SHFTDP\;
  OUTPUTS.\THRST-\     <= \THRST-\;
  OUTPUTS.\LRZVEL\     <= \LRZVEL\;
  OUTPUTS.\SHFTDM\     <= \SHFTDM\;
  OUTPUTS.\EMS+\       <= \EMS+\;
  OUTPUTS.\LRYVEL\     <= \LRYVEL\;
  OUTPUTS.\TRNDP\      <= \TRNDP\;
  OUTPUTS.\EMS-\       <= \EMS-\;
  OUTPUTS.\LRXVEL\     <= \LRXVEL\;
  OUTPUTS.\TRNDM\      <= \TRNDM\;
  OUTPUTS.\ALT1\       <= \ALT1\;
  OUTPUTS.\RRRANG\     <= \RRRANG\;
  OUTPUTS.\GYRSET\     <= \GYRSET\;
  OUTPUTS.\ALT0\       <= \ALT0\;
  OUTPUTS.\RRRARA\     <= \RRRARA\;
  OUTPUTS.\GYRRST\     <= \GYRRST\;
  OUTPUTS.\ALRT1\      <= \ALRT1\;
  OUTPUTS.\RRSYNC\     <= \RRSYNC\;
  OUTPUTS.\OTLNK0\     <= \OTLNK0\;
  OUTPUTS.\ALRT0\      <= \ALRT0\;
  OUTPUTS.\LRSYNC\     <= \LRSYNC\;
  OUTPUTS.\OTLNK1\     <= \OTLNK1\;
  OUTPUTS.\DKDATB\     <= \DKDATB\;
  OUTPUTS.\DKDATA\     <= \DKDATA\;
  OUTPUTS.\GYZM\       <= \GYZM\;
  OUTPUTS.\GYYM\       <= \GYYM\;
  OUTPUTS.\GYXM\       <= \GYXM\;
  OUTPUTS.\GYZP\       <= \GYZP\;
  OUTPUTS.\GYYP\       <= \GYYP\;
  OUTPUTS.\GYXP\       <= \GYXP\;

  SYSERROR <=    not( \11B\ ) -- MDT01 (latched and inverted MPAL/   ) PARITY FAIL (E OR F MEMORY).
              or not( \13B\ ) -- MDT02 (latched              MT05    ) PARITY FAIL (E MEMORY).
              or not( \14B\ ) -- MDT03 (latched and inverted MTCAL/  ) TC TRAP.
              or not( \15B\ ) -- MDT04 (latched and inverted MRPTAL/ ) RUPT LOCK.
              or not( \16B\ ) -- MDT05 (latched and inverted MWATCH/ ) NIGHT WATCHMAN.
              or not( \17B\ ) -- MDT06 (latched and inverted MVFAIL/ ) VOLTAGE FAIL.
              or not( \18B\ ) -- MDT07 (latched and inverted MCTRAL/ ) COUNTER FAIL.
              or not( \19B\ ) -- MDT08 (latched and inverted MSCAFL/ ) SCALER FAIL.
              or not( \20B\ ) -- MDT09 (latched and inverted MSCDBL/ ) SCALER DOUBLE FREQUENCY ALARM.
              or \STOP\;

  VGADEBUG(  0,  0 ) <= not \11B\; -- MDT01 (latched and inverted MPAL/   ) PARITY FAIL (E OR F MEMORY).
  VGADEBUG(  1,  0 ) <= not \13B\; -- MDT02 (latched              MT05    ) PARITY FAIL (E MEMORY).
  VGADEBUG(  2,  0 ) <= not \14B\; -- MDT03 (latched and inverted MTCAL/  ) TC TRAP.
  VGADEBUG(  3,  0 ) <= not \15B\; -- MDT04 (latched and inverted MRPTAL/ ) RUPT LOCK.
  VGADEBUG(  4,  0 ) <= not \16B\; -- MDT05 (latched and inverted MWATCH/ ) NIGHT WATCHMAN.
  VGADEBUG(  5,  0 ) <= not \17B\; -- MDT06 (latched and inverted MVFAIL/ ) VOLTAGE FAIL.
  VGADEBUG(  6,  0 ) <= not \18B\; -- MDT07 (latched and inverted MCTRAL/ ) COUNTER FAIL.
  VGADEBUG(  7,  0 ) <= not \19B\; -- MDT08 (latched and inverted MSCAFL/ ) SCALER FAIL.
  VGADEBUG(  8,  0 ) <= not \20B\; -- MDT09 (latched and inverted MSCDBL/ ) SCALER DOUBLE FREQUENCY ALARM.
  VGADEBUG(  9,  0 ) <= \STOP\;
  VGADEBUG( 10,  0 ) <= \STOPA\;
  VGADEBUG( 11,  0 ) <= \SBY\;
  VGADEBUG( 12,  0 ) <= \ALGA\;
  VGADEBUG( 13,  0 ) <= \STRT1\;
  VGADEBUG( 14,  0 ) <= \STRT2\;
  VGADEBUG( 15,  0 ) <= \GOJAM\;

  VGADEBUG(  0,  1 ) <= \CLOCK\;
  VGADEBUG(  1,  1 ) <= \CLK\;
  VGADEBUG(  2,  1 ) <= not \RINGA/\;
  VGADEBUG(  3,  1 ) <= not \RINGB/\;
  VGADEBUG(  4,  1 ) <= not \ODDSET/\;
  VGADEBUG(  5,  1 ) <= not \EVNSET/\;

  VGADEBUG(  0,  2 ) <= \T01\;
  VGADEBUG(  1,  2 ) <= \T02\;
  VGADEBUG(  2,  2 ) <= \T03\;
  VGADEBUG(  3,  2 ) <= \T04\;
  VGADEBUG(  4,  2 ) <= \T05\;
  VGADEBUG(  5,  2 ) <= \T06\;
  VGADEBUG(  6,  2 ) <= \T07\;
  VGADEBUG(  7,  2 ) <= \T08\;
  VGADEBUG(  8,  2 ) <= \T09\;
  VGADEBUG(  9,  2 ) <= \T10\;
  VGADEBUG( 10,  2 ) <= \T11\;
  VGADEBUG( 11,  2 ) <= \T12\;
  VGADEBUG( 12,  2 ) <= \T12SET\;
  --        13
  VGADEBUG( 14,  2 ) <= \P01\;
  VGADEBUG( 15,  2 ) <= \P02\;
  VGADEBUG( 16,  2 ) <= \P03\;
  VGADEBUG( 17,  2 ) <= \P04\;
  VGADEBUG( 18,  2 ) <= \P05\;
  VGADEBUG( 19,  2 ) <= not \P01/\;
  VGADEBUG( 20,  2 ) <= not \P02/\;
  VGADEBUG( 21,  2 ) <= not \P03/\;
  VGADEBUG( 22,  2 ) <= not \P04/\;
  VGADEBUG( 23,  2 ) <= not \P05/\;
  VGADEBUG( 24,  2 ) <= \SB0\;
  VGADEBUG( 25,  2 ) <= \SB1\;
  VGADEBUG( 26,  2 ) <= \SB2\;
  VGADEBUG( 27,  2 ) <= \SB4\;
  VGADEBUG( 28,  2 ) <= \EDSET\;

  VGADEBUG(  0,  3 ) <= \FS01\;
  VGADEBUG(  1,  3 ) <= \FS02\;
  VGADEBUG(  2,  3 ) <= \FS03\;
  VGADEBUG(  3,  3 ) <= \FS04\;
  VGADEBUG(  4,  3 ) <= \FS05\;
  VGADEBUG(  5,  3 ) <= \FS06\;
  VGADEBUG(  6,  3 ) <= \FS07\;
  VGADEBUG(  7,  3 ) <= \FS08\;
  VGADEBUG(  8,  3 ) <= \FS09\;
  VGADEBUG(  9,  3 ) <= \FS10\;
  VGADEBUG( 10,  3 ) <= \FS11\;
  VGADEBUG( 11,  3 ) <= \FS12\;
  VGADEBUG( 12,  3 ) <= \FS13\;
  VGADEBUG( 13,  3 ) <= \FS14\;
  VGADEBUG( 14,  3 ) <= \FS15\;
  VGADEBUG( 15,  3 ) <= \FS16\;
  VGADEBUG( 16,  3 ) <= \FS17\;
  VGADEBUG( 17,  3 ) <= \FS18\;
  VGADEBUG( 18,  3 ) <= \FS19\;
  VGADEBUG( 19,  3 ) <= \FS20\;
  VGADEBUG( 20,  3 ) <= \FS21\;
  VGADEBUG( 21,  3 ) <= \FS22\;
  VGADEBUG( 22,  3 ) <= \FS23\;
  VGADEBUG( 23,  3 ) <= \FS24\;
  VGADEBUG( 24,  3 ) <= \FS25\;
  VGADEBUG( 25,  3 ) <= \FS26\;
  VGADEBUG( 26,  3 ) <= \FS27\;
  VGADEBUG( 27,  3 ) <= \FS28\;
  VGADEBUG( 28,  3 ) <= \FS29\;
  VGADEBUG( 29,  3 ) <= \FS30\;
  VGADEBUG( 30,  3 ) <= \FS31\;
  VGADEBUG( 31,  3 ) <= \FS32\;
  VGADEBUG( 32,  3 ) <= \FS33\;

  VGADEBUG(  0,  4 ) <= \SAP\;
  VGADEBUG(  1,  4 ) <= \SA01\;
  VGADEBUG(  2,  4 ) <= \SA02\;
  VGADEBUG(  3,  4 ) <= \SA03\;
  VGADEBUG(  4,  4 ) <= \SA04\;
  VGADEBUG(  5,  4 ) <= \SA05\;
  VGADEBUG(  6,  4 ) <= \SA06\;
  VGADEBUG(  7,  4 ) <= \SA07\;
  VGADEBUG(  8,  4 ) <= \SA08\;
  VGADEBUG(  9,  4 ) <= \SA09\;
  VGADEBUG( 10,  4 ) <= \SA10\;
  VGADEBUG( 11,  4 ) <= \SA11\;
  VGADEBUG( 12,  4 ) <= \SA12\;
  VGADEBUG( 13,  4 ) <= \SA13\;
  VGADEBUG( 14,  4 ) <= \SA14\;
  VGADEBUG( 15,  4 ) <= \SA16\;
  --        16
  --        17
  --        18
  VGADEBUG( 19,  4 ) <= \SBE\;   -- EREAD
  VGADEBUG( 20,  4 ) <= \ZID\;   -- EWRITE
  VGADEBUG( 21,  4 ) <= \SETEK\; -- ESTART
  VGADEBUG( 22,  4 ) <= \SBF\;   -- FREAD

  VGADEBUG(  0,  5 ) <= \GEMP\;
  VGADEBUG(  1,  5 ) <= \GEM01\;
  VGADEBUG(  2,  5 ) <= \GEM02\;
  VGADEBUG(  3,  5 ) <= \GEM03\;
  VGADEBUG(  4,  5 ) <= \GEM04\;
  VGADEBUG(  5,  5 ) <= \GEM05\;
  VGADEBUG(  6,  5 ) <= \GEM06\;
  VGADEBUG(  7,  5 ) <= \GEM07\;
  VGADEBUG(  8,  5 ) <= \GEM08\;
  VGADEBUG(  9,  5 ) <= \GEM09\;
  VGADEBUG( 10,  5 ) <= \GEM10\;
  VGADEBUG( 11,  5 ) <= \GEM11\;
  VGADEBUG( 12,  5 ) <= \GEM12\;
  VGADEBUG( 13,  5 ) <= \GEM13\;
  VGADEBUG( 14,  5 ) <= \GEM14\;
  VGADEBUG( 15,  5 ) <= \GEM16\;
  --        16
  --        17
  --        18
  VGADEBUG( 19,  5 ) <= \SBE\;   -- EREAD
  VGADEBUG( 20,  5 ) <= \ZID\;   -- EWRITE
  VGADEBUG( 21,  5 ) <= \SETEK\; -- ESTART
  --        22

  VGADEBUG(  0,  6 ) <= \S01\;
  VGADEBUG(  1,  6 ) <= \S02\;
  VGADEBUG(  2,  6 ) <= \S03\;
  VGADEBUG(  3,  6 ) <= \S04\;
  VGADEBUG(  4,  6 ) <= \S05\;
  VGADEBUG(  5,  6 ) <= \S06\;
  VGADEBUG(  6,  6 ) <= \S07\;
  VGADEBUG(  7,  6 ) <= \S08\;
  VGADEBUG(  8,  6 ) <= \EAD09\;
  VGADEBUG(  9,  6 ) <= \EAD10\;
  VGADEBUG( 10,  6 ) <= \EAD11\;
  --        11
  --        12
  --        13
  --        14
  --        15
  --        16
  --        17
  --        18
  VGADEBUG( 19,  6 ) <= \SBE\;   -- EREAD
  VGADEBUG( 20,  6 ) <= \ZID\;   -- EWRITE
  VGADEBUG( 21,  6 ) <= \SETEK\; -- ESTART
  --        22

  VGADEBUG(  0,  7 ) <= \S01\;
  VGADEBUG(  1,  7 ) <= \S02\;
  VGADEBUG(  2,  7 ) <= \S03\;
  VGADEBUG(  3,  7 ) <= \S04\;
  VGADEBUG(  4,  7 ) <= \S05\;
  VGADEBUG(  5,  7 ) <= \S06\;
  VGADEBUG(  6,  7 ) <= \S07\;
  VGADEBUG(  7,  7 ) <= \S08\;
  VGADEBUG(  8,  7 ) <= \S09\;
  VGADEBUG(  9,  7 ) <= \S10\;
  VGADEBUG( 10,  7 ) <= \F11\;
  VGADEBUG( 11,  7 ) <= \F12\;
  VGADEBUG( 12,  7 ) <= \F13\;
  VGADEBUG( 13,  7 ) <= \F14\;
  VGADEBUG( 14,  7 ) <= \F15\;
  VGADEBUG( 15,  7 ) <= \F16\;
  --        16
  --        17
  --        18
  --        19
  --        20
  --        21
  VGADEBUG( 22,  7 ) <= \SBF\;   -- FREAD

  VGADEBUG(  0,  8 ) <= \S01\;
  VGADEBUG(  1,  8 ) <= \S02\;
  VGADEBUG(  2,  8 ) <= \S03\;
  VGADEBUG(  3,  8 ) <= \S04\;
  VGADEBUG(  4,  8 ) <= \S05\;
  VGADEBUG(  5,  8 ) <= \S06\;
  VGADEBUG(  6,  8 ) <= \S07\;
  VGADEBUG(  7,  8 ) <= \S08\;
  VGADEBUG(  8,  8 ) <= \S09\;
  VGADEBUG(  9,  8 ) <= \S10\;
  VGADEBUG( 10,  8 ) <= \S11\;
  VGADEBUG( 11,  8 ) <= \S12\;

  VGADEBUG(  9,  9 ) <= \MSQ10\;
  VGADEBUG( 10,  9 ) <= \MSQ11\;
  VGADEBUG( 11,  9 ) <= \MSQ12\;
  VGADEBUG( 12,  9 ) <= \MSQ13\;
  VGADEBUG( 13,  9 ) <= \MSQ14\;
  --        14
  VGADEBUG( 15,  9 ) <= \MSQ16\;
  VGADEBUG( 16,  9 ) <= \MSQEXT\;
  --        17
  --        18
  VGADEBUG( 19,  9 ) <= \CSQG\;
  VGADEBUG( 20,  9 ) <= not \WSQG/\;

  VGADEBUG(  0, 10 ) <= \WL01\;
  VGADEBUG(  1, 10 ) <= \WL02\;
  VGADEBUG(  2, 10 ) <= \WL03\;
  VGADEBUG(  3, 10 ) <= \WL04\;
  VGADEBUG(  4, 10 ) <= \WL05\;
  VGADEBUG(  5, 10 ) <= \WL06\;
  VGADEBUG(  6, 10 ) <= \WL07\;
  VGADEBUG(  7, 10 ) <= \WL08\;
  VGADEBUG(  8, 10 ) <= \WL09\;
  VGADEBUG(  9, 10 ) <= \WL10\;
  VGADEBUG( 10, 10 ) <= \WL11\;
  VGADEBUG( 11, 10 ) <= \WL12\;
  VGADEBUG( 12, 10 ) <= \WL13\;
  VGADEBUG( 13, 10 ) <= \WL14\;
  VGADEBUG( 14, 10 ) <= \WL15\;
  VGADEBUG( 15, 10 ) <= \WL16\;

  VGADEBUG(  0, 11 ) <= not \51103\; -- X01
  VGADEBUG(  1, 11 ) <= not \51203\; -- X02
  VGADEBUG(  2, 11 ) <= not \51403\; -- X03
  VGADEBUG(  3, 11 ) <= not \51303\; -- X04
  VGADEBUG(  4, 11 ) <= not \52103\; -- X05
  VGADEBUG(  5, 11 ) <= not \52203\; -- X06
  VGADEBUG(  6, 11 ) <= not \52403\; -- X07
  VGADEBUG(  7, 11 ) <= not \52303\; -- X08
  VGADEBUG(  8, 11 ) <= not \53103\; -- X09
  VGADEBUG(  9, 11 ) <= not \53203\; -- X10
  VGADEBUG( 10, 11 ) <= not \53403\; -- X11
  VGADEBUG( 11, 11 ) <= not \53303\; -- X12
  VGADEBUG( 12, 11 ) <= not \54103\; -- X13
  VGADEBUG( 13, 11 ) <= not \54203\; -- X14
  VGADEBUG( 14, 11 ) <= not \54403\; -- X15
  VGADEBUG( 15, 11 ) <= not \54303\; -- X16

  VGADEBUG(  0, 12 ) <= not \51107\; -- Y01
  VGADEBUG(  1, 12 ) <= not \51207\; -- Y02
  VGADEBUG(  2, 12 ) <= not \51407\; -- Y03
  VGADEBUG(  3, 12 ) <= not \51307\; -- Y04
  VGADEBUG(  4, 12 ) <= not \52107\; -- Y05
  VGADEBUG(  5, 12 ) <= not \52207\; -- Y06
  VGADEBUG(  6, 12 ) <= not \53407\; -- Y07
  VGADEBUG(  7, 12 ) <= not \52307\; -- Y08
  VGADEBUG(  8, 12 ) <= not \53107\; -- Y09
  VGADEBUG(  9, 12 ) <= not \53207\; -- Y10
  VGADEBUG( 10, 12 ) <= not \53407\; -- Y11
  VGADEBUG( 11, 12 ) <= not \53307\; -- Y12
  VGADEBUG( 12, 12 ) <= not \54107\; -- Y13
  VGADEBUG( 13, 12 ) <= not \54207\; -- Y14
  VGADEBUG( 14, 12 ) <= not \54407\; -- Y15
  VGADEBUG( 15, 12 ) <= not \54307\; -- Y16

  VGADEBUG(  0, 13 ) <= not \A01/\; -- A01
  VGADEBUG(  1, 13 ) <= not \A02/\; -- A02
  VGADEBUG(  2, 13 ) <= not \A03/\; -- A03
  VGADEBUG(  3, 13 ) <= not \A04/\; -- A04
  VGADEBUG(  4, 13 ) <= not \A05/\; -- A05
  VGADEBUG(  5, 13 ) <= not \A06/\; -- A06
  VGADEBUG(  6, 13 ) <= not \A07/\; -- A07
  VGADEBUG(  7, 13 ) <= not \A08/\; -- A08
  VGADEBUG(  8, 13 ) <= not \A09/\; -- A09
  VGADEBUG(  9, 13 ) <= not \A10/\; -- A10
  VGADEBUG( 10, 13 ) <= not \A11/\; -- A11
  VGADEBUG( 11, 13 ) <= not \A12/\; -- A12
  VGADEBUG( 12, 13 ) <= not \A13/\; -- A13
  VGADEBUG( 13, 13 ) <= not \A14/\; -- A14
  VGADEBUG( 14, 13 ) <= not \A15/\; -- A15
  VGADEBUG( 15, 13 ) <= not \A16/\; -- A16

  VGADEBUG(  0, 14 ) <= not \L01/\; -- L01
  VGADEBUG(  1, 14 ) <= not \L02/\; -- L02
  VGADEBUG(  2, 14 ) <= not \L03/\; -- L03
  VGADEBUG(  3, 14 ) <= not \L04/\; -- L04
  VGADEBUG(  4, 14 ) <= not \L05/\; -- L05
  VGADEBUG(  5, 14 ) <= not \L06/\; -- L06
  VGADEBUG(  6, 14 ) <= not \L07/\; -- L07
  VGADEBUG(  7, 14 ) <= not \L08/\; -- L08
  VGADEBUG(  8, 14 ) <= not \L09/\; -- L09
  VGADEBUG(  9, 14 ) <= not \L10/\; -- L10
  VGADEBUG( 10, 14 ) <= not \L11/\; -- L11
  VGADEBUG( 11, 14 ) <= not \L12/\; -- L12
  VGADEBUG( 12, 14 ) <= not \L13/\; -- L13
  VGADEBUG( 13, 14 ) <= not \L14/\; -- L14
  VGADEBUG( 14, 14 ) <= not \L15/\; -- L15
  VGADEBUG( 15, 14 ) <= not \L16/\; -- L16

  VGADEBUG(  0, 15 ) <= not \51130\; -- Q01
  VGADEBUG(  1, 15 ) <= not \51230\; -- Q02
  VGADEBUG(  2, 15 ) <= not \51430\; -- Q03
  VGADEBUG(  3, 15 ) <= not \51330\; -- Q04
  VGADEBUG(  4, 15 ) <= not \52130\; -- Q05
  VGADEBUG(  5, 15 ) <= not \52230\; -- Q06
  VGADEBUG(  6, 15 ) <= not \52430\; -- Q07
  VGADEBUG(  7, 15 ) <= not \52330\; -- Q08
  VGADEBUG(  8, 15 ) <= not \53130\; -- Q09
  VGADEBUG(  9, 15 ) <= not \53230\; -- Q10
  VGADEBUG( 10, 15 ) <= not \53430\; -- Q11
  VGADEBUG( 11, 15 ) <= not \53330\; -- Q12
  VGADEBUG( 12, 15 ) <= not \54130\; -- Q13
  VGADEBUG( 13, 15 ) <= not \54230\; -- Q14
  VGADEBUG( 14, 15 ) <= not \54430\; -- Q15
  VGADEBUG( 15, 15 ) <= not \54330\; -- Q16

  VGADEBUG(  0, 16 ) <= not \Z01/\; -- Z01
  VGADEBUG(  1, 16 ) <= not \Z02/\; -- Z02
  VGADEBUG(  2, 16 ) <= not \Z03/\; -- Z03
  VGADEBUG(  3, 16 ) <= not \Z04/\; -- Z04
  VGADEBUG(  4, 16 ) <= not \Z05/\; -- Z05
  VGADEBUG(  5, 16 ) <= not \Z06/\; -- Z06
  VGADEBUG(  6, 16 ) <= not \Z07/\; -- Z07
  VGADEBUG(  7, 16 ) <= not \Z08/\; -- Z08
  VGADEBUG(  8, 16 ) <= not \Z09/\; -- Z09
  VGADEBUG(  9, 16 ) <= not \Z10/\; -- Z10
  VGADEBUG( 10, 16 ) <= not \Z11/\; -- Z11
  VGADEBUG( 11, 16 ) <= not \Z12/\; -- Z12
  VGADEBUG( 12, 16 ) <= not \Z13/\; -- Z13
  VGADEBUG( 13, 16 ) <= not \Z14/\; -- Z14
  VGADEBUG( 14, 16 ) <= not \Z15/\; -- Z15
  VGADEBUG( 15, 16 ) <= not \Z16/\; -- Z16

  VGADEBUG(  0, 17 ) <= not \51139\; -- B01
  VGADEBUG(  1, 17 ) <= not \51239\; -- B02
  VGADEBUG(  2, 17 ) <= not \51439\; -- B03
  VGADEBUG(  3, 17 ) <= not \51339\; -- B04
  VGADEBUG(  4, 17 ) <= not \52139\; -- B05
  VGADEBUG(  5, 17 ) <= not \52239\; -- B06
  VGADEBUG(  6, 17 ) <= not \52439\; -- B07
  VGADEBUG(  7, 17 ) <= not \52339\; -- B08
  VGADEBUG(  8, 17 ) <= not \53139\; -- B09
  VGADEBUG(  9, 17 ) <= not \53239\; -- B10
  VGADEBUG( 10, 17 ) <= not \53439\; -- B11
  VGADEBUG( 11, 17 ) <= not \53339\; -- B12
  VGADEBUG( 12, 17 ) <= not \54139\; -- B13
  VGADEBUG( 13, 17 ) <= not \54239\; -- B14
  VGADEBUG( 14, 17 ) <= not \54439\; -- B15
  VGADEBUG( 15, 17 ) <= not \54339\; -- B16

  VGADEBUG(  0, 18 ) <= \51139\; -- C01
  VGADEBUG(  1, 18 ) <= \51239\; -- C02
  VGADEBUG(  2, 18 ) <= \51439\; -- C03
  VGADEBUG(  3, 18 ) <= \51339\; -- C04
  VGADEBUG(  4, 18 ) <= \52139\; -- C05
  VGADEBUG(  5, 18 ) <= \52239\; -- C06
  VGADEBUG(  6, 18 ) <= \52439\; -- C07
  VGADEBUG(  7, 18 ) <= \52339\; -- C08
  VGADEBUG(  8, 18 ) <= \53139\; -- C09
  VGADEBUG(  9, 18 ) <= \53239\; -- C10
  VGADEBUG( 10, 18 ) <= \53439\; -- C11
  VGADEBUG( 11, 18 ) <= \53339\; -- C12
  VGADEBUG( 12, 18 ) <= \54139\; -- C13
  VGADEBUG( 13, 18 ) <= \54239\; -- C14
  VGADEBUG( 14, 18 ) <= \54439\; -- C15
  VGADEBUG( 15, 18 ) <= \54339\; -- C16

  VGADEBUG(  0, 19 ) <= not \G01/\; -- G01
  VGADEBUG(  1, 19 ) <= not \G02/\; -- G02
  VGADEBUG(  2, 19 ) <= not \G03/\; -- G03
  VGADEBUG(  3, 19 ) <= not \G04/\; -- G04
  VGADEBUG(  4, 19 ) <= not \G05/\; -- G05
  VGADEBUG(  5, 19 ) <= not \G06/\; -- G06
  VGADEBUG(  6, 19 ) <= not \G07/\; -- G07
  VGADEBUG(  7, 19 ) <= not \G08/\; -- G08
  VGADEBUG(  8, 19 ) <= not \G09/\; -- G09
  VGADEBUG(  9, 19 ) <= not \G10/\; -- G10
  VGADEBUG( 10, 19 ) <= not \G11/\; -- G11
  VGADEBUG( 11, 19 ) <= not \G12/\; -- G12
  VGADEBUG( 12, 19 ) <= not \G13/\; -- G13
  VGADEBUG( 13, 19 ) <= not \G14/\; -- G14
  VGADEBUG( 14, 19 ) <= not \G15/\; -- G15
  VGADEBUG( 15, 19 ) <= not \G16/\; -- G16

  VGADEBUG(  0, 21 ) <= \XT0\;
  VGADEBUG(  1, 21 ) <= \XT1\;
  VGADEBUG(  2, 21 ) <= \XT2\;
  VGADEBUG(  3, 21 ) <= \XT3\;
  VGADEBUG(  4, 21 ) <= \XT4\;
  VGADEBUG(  5, 21 ) <= \XT5\;
  VGADEBUG(  6, 21 ) <= \XT6\;
  VGADEBUG(  7, 21 ) <= \XT7\;
  VGADEBUG(  8, 21 ) <= \XB0\;
  VGADEBUG(  9, 21 ) <= \XB1\;
  VGADEBUG( 10, 21 ) <= \XB2\;
  VGADEBUG( 11, 21 ) <= \XB3\;
  VGADEBUG( 12, 21 ) <= \XB4\;
  VGADEBUG( 13, 21 ) <= \XB5\;
  VGADEBUG( 14, 21 ) <= \XB6\;
  VGADEBUG( 15, 21 ) <= \XB7\;
  VGADEBUG( 16, 21 ) <= \YB0\;
  VGADEBUG( 17, 21 ) <= \YB1\;
  VGADEBUG( 18, 21 ) <= \YB2\;
  VGADEBUG( 19, 21 ) <= \YB3\;

  VGADEBUG(  3, 22 ) <= not \RCHBT/\;
  VGADEBUG(  4, 22 ) <= not \RCHAT/\;
  VGADEBUG( 10, 22 ) <= not \WCH10/\;
  VGADEBUG( 11, 22 ) <= not \WCH11/\;
  VGADEBUG( 32, 22 ) <= not \RCH32/\;

  VGADEBUG(  0, 23 ) <= \RLYB01\;
  VGADEBUG(  1, 23 ) <= \RLYB02\;
  VGADEBUG(  2, 23 ) <= \RLYB03\;
  VGADEBUG(  3, 23 ) <= \RLYB04\;
  VGADEBUG(  4, 23 ) <= \RLYB05\;
  VGADEBUG(  5, 23 ) <= \RLYB06\;
  VGADEBUG(  6, 23 ) <= \RLYB07\;
  VGADEBUG(  7, 23 ) <= \RLYB08\;
  VGADEBUG(  8, 23 ) <= \RLYB09\;
  VGADEBUG(  9, 23 ) <= \RLYB10\;
  VGADEBUG( 10, 23 ) <= \RLYB11\;
  VGADEBUG( 11, 23 ) <= \RYWD12\;
  VGADEBUG( 12, 23 ) <= \RYWD13\;
  VGADEBUG( 13, 23 ) <= \RYWD14\;
  VGADEBUG( 14, 23 ) <= \RYWD16\;
  --        15
  --        16
  --        17
  --        18
  --        19
  VGADEBUG( 20, 23 ) <= not \WCH10/\;

  VGADEBUG(  0, 24 ) <= \ISSWAR\;
  VGADEBUG(  1, 24 ) <= \COMACT\;
  VGADEBUG(  2, 24 ) <= \UPLACT\;
  VGADEBUG(  3, 24 ) <= \TMPOUT\;
  VGADEBUG(  4, 24 ) <= not \43430\; -- KYRLS
  VGADEBUG(  5, 24 ) <= not \43434\; -- VNFLSH
  VGADEBUG(  6, 24 ) <= not \43444\; -- OPEROR
  VGADEBUG(  7, 24 ) <= \OT1108\;
  VGADEBUG(  8, 24 ) <= not \FF1109/\;
  VGADEBUG(  9, 24 ) <= not \FF1110/\;
  VGADEBUG( 10, 24 ) <= not \FF1111/\;
  VGADEBUG( 11, 24 ) <= not \FF1112/\;
  VGADEBUG( 12, 24 ) <= \OT1113\;
  VGADEBUG( 13, 24 ) <= \OT1114\;
  VGADEBUG( 14, 24 ) <= \OT1116\;
  --        15
  --        16
  --        17
  --        18
  --        19
  VGADEBUG( 20, 24 ) <= not \WCH11/\;

  VGADEBUG(  0, 25 ) <= INPUTS.\MAINRS\;
  VGADEBUG(  1, 25 ) <= INPUTS.\IN3214\;
  VGADEBUG(  2, 25 ) <= INPUTS.\MKEY5\;
  VGADEBUG(  3, 25 ) <= INPUTS.\MKEY4\;
  VGADEBUG(  4, 25 ) <= INPUTS.\MKEY3\;
  VGADEBUG(  5, 25 ) <= INPUTS.\MKEY2\;
  VGADEBUG(  6, 25 ) <= INPUTS.\MKEY1\;
  --         7
  VGADEBUG(  8, 25 ) <= \35322\;
  VGADEBUG(  9, 25 ) <= not \35323\;

  VGADEBUG(  0, 28 ) <= not \MRPTAL/\; -- DEBUG
  VGADEBUG(  1, 28 ) <= \F14H\; -- DEBUG
  VGADEBUG(  2, 28 ) <= \F14B\; -- DEBUG
  VGADEBUG(  3, 28 ) <= \MIIP\; -- DEBUG
  VGADEBUG(  4, 28 ) <= \MINHL\; -- DEBUG
  VGADEBUG(  5, 28 ) <= \KRPT\; -- DEBUG
  VGADEBUG(  6, 28 ) <= \RUPT0\; -- DEBUG
  VGADEBUG(  7, 28 ) <= \RUPT1\; -- DEBUG
  VGADEBUG(  8, 28 ) <= \INHPLS\; -- DEBUG
  VGADEBUG(  9, 28 ) <= \RELPLS\; -- DEBUG
  VGADEBUG( 10, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 11, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 12, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 13, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 14, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 15, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 16, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 17, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 18, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 19, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 20, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 21, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 22, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 23, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 24, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 25, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 26, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 27, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 28, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 29, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 30, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 31, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 32, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 33, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 34, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 35, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 36, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 37, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 38, 28 ) <= '0'; -- DEBUG
  VGADEBUG( 39, 28 ) <= '0'; -- DEBUG

  VGADEBUG(  0, 29 ) <= \PA03\; -- DEBUG
  VGADEBUG(  1, 29 ) <= \PA06\; -- DEBUG
  VGADEBUG(  2, 29 ) <= \PA09\; -- DEBUG
  VGADEBUG(  3, 29 ) <= \PA12\; -- DEBUG
  VGADEBUG(  4, 29 ) <= \PA15\; -- DEBUG
  VGADEBUG(  5, 29 ) <= \PB09\; -- DEBUG
  VGADEBUG(  6, 29 ) <= \PB15\; -- DEBUG
  VGADEBUG(  7, 29 ) <= \PC15\; -- DEBUG
  VGADEBUG(  8, 29 ) <= '0'; -- DEBUG
  VGADEBUG(  9, 29 ) <= \CGG\; -- DEBUG
  VGADEBUG( 10, 29 ) <= \MONPAR\; -- DEBUG
  VGADEBUG( 11, 29 ) <= \SAP\; -- DEBUG
  VGADEBUG( 12, 29 ) <= \GEMP\; -- DEBUG
  VGADEBUG( 13, 29 ) <= \MSP\; -- DEBUG
  VGADEBUG( 14, 29 ) <= \SCAD\; -- DEBUG
  VGADEBUG( 15, 29 ) <= not \TPARG/\; -- DEBUG
  VGADEBUG( 16, 29 ) <= \8XP5\; -- DEBUG
  VGADEBUG( 17, 29 ) <= \PALE\; -- DEBUG
  VGADEBUG( 18, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 19, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 20, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 21, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 22, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 23, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 24, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 25, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 26, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 27, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 28, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 29, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 30, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 31, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 32, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 33, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 34, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 35, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 36, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 37, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 38, 29 ) <= '0'; -- DEBUG
  VGADEBUG( 39, 29 ) <= '0'; -- DEBUG

end Rtl;

-- **********************
-- ***                ***
-- ***  END OF FILE.  ***
-- ***                ***
-- **********************

