`ifdef ATCBUSDEC301_CONST_VH
`else
`define ATCBUSDEC301_CONST_VH

`define ATCBUSDEC301_PRODUCT_ID			32'h00033003

`ifdef ATCBUSDEC301_ADDR_WIDTH_24
`define ATCBUSDEC301_ADDR_WIDTH			24
`else
`ifndef ATCBUSDEC301_ADDR_WIDTH
`define ATCBUSDEC301_ADDR_WIDTH			32
`endif
`endif

`define ATCBUSDEC301_ADDR_MSB			(`ATCBUSDEC301_ADDR_WIDTH-1)

`ifdef ATCBUSDEC301_DATA_WIDTH_256
`define ATCBUSDEC301_DATA_WIDTH 256
`else
`ifdef ATCBUSDEC301_DATA_WIDTH_128
`define ATCBUSDEC301_DATA_WIDTH 128
`else
`ifdef ATCBUSDEC301_DATA_WIDTH_64
`define ATCBUSDEC301_DATA_WIDTH 64
`else
`define ATCBUSDEC301_DATA_WIDTH_32
`define ATCBUSDEC301_DATA_WIDTH 32
`endif
`endif
`endif

`define ATCBUSDEC301_SLV_0
`define	ATCBUSDEC301_SLV0_SIZE			1
`ifdef ATCBUSDEC301_SLV0_OFFSET
`else
`define	ATCBUSDEC301_SLV0_OFFSET		`ATCBUSDEC301_ADDR_DECODE_WIDTH'h0
`endif

`endif
