
// Copyright (c) 2006-2013 Arteris, Inc. All rights reserved.
// Copyright (c) 2013-2020 Qualcomm Technologies, Inc. All rights reserved.
// These files contain material which is the Confidential Information of Arteris and which is protected by various intellectual property rights.
// You may make, have made, use, reproduce, display or perform (publicly or otherwise), prepare
// derivative works based on, offer for sale, sell, distribute, import,
// disclose, license, sublicense, dispose of and otherwise exploit this RTL solely in
// accordance with your license agreement with Arteris, Inc or Arteris IP, SAS.
// If you have not agreed to all of the terms and conditions in such License
// Agreement, you should immediately return these files (including any copies)
// to your licensor Arteris, Inc or Arteris IP, SAS.
// The material in these files or portions thereof are protected under U.S. and foreign patent and patent applications.
// This software and hardware IP product is protected by patents as described at http://www.arteris.com/patents.


// Generated by FlexNoC
// Tool Version 4.7.0
// Platform     centos:7
// Date         Tue Sep 13 13:44:24 2022


// FlexNoC version    : 4.7.0
// PDD File           : /home/aptashko/GEMINI/design/ip/FlexNoC/rsnoc_arch_edit.pdd
// Exported Structure : /Specification.Architecture.Structure
// ExportOption       : /verilog

`timescale 1ps/1ps
module rsnoc_z_T_C_S_C_L_S_Ce_R ( En , I , O );
	input   En ;
	input   I  ;
	output  O  ;
//	reg  LatchedEn ;
//	always @( I or En )		if ( I == 0)
//			LatchedEn <= #1.0 ( En );
//assign O = LatchedEn && I;
assign O = I;
endmodule

`ifndef SIM_GATERCELL_RSTASYNC
`define SIM_GATERCELL_RSTASYNC
`timescale 1ps/1ps
module GaterCell_RstAsync ( CLKIN , CLKOUT , EN , RSTN , TE );
	input   CLKIN  ;
	output  CLKOUT ;
	input   EN     ;
	input   RSTN   ;
	input   TE     ;
	rsnoc_z_T_C_S_C_L_S_Ce_R uce( .En( EN | TE ) , .I( CLKIN ) , .O( CLKOUT ) );
endmodule
`endif


