`ifdef ATCBMC300_CONFIG_VH
`else
`define ATCBMC300_CONFIG_VH
`include "config.inc"
`include "ae350_config.vh"
`include "ae350_const.vh"

`ifdef  PLATFORM_FORCE_4GB_SPACE 
        `define ATCBMC300_ADDR_WIDTH 32
`else  //~PLATFORM_FORCE_4GB_SPACE 
        `ifdef NDS_BIU_ADDR_WIDTH
                `define ATCBMC300_ADDR_WIDTH `NDS_BIU_ADDR_WIDTH
        `else
                `define ATCBMC300_ADDR_WIDTH 32
        `endif
`endif  //PLATFORM_FORCE_4GB_SPACE 

`define ATCBMC300_ID_WIDTH   `AE350_AXI_ID_WIDTH
`ifdef NDS_L2C_BIU_DATA_WIDTH
	`define ATCBMC300_DATA_WIDTH `NDS_L2C_BIU_DATA_WIDTH
`else
	`define ATCBMC300_DATA_WIDTH `NDS_BIU_DATA_WIDTH
`endif

//-------------------------------------------------
// AXI Master Ports
//-------------------------------------------------

`ifdef NDS_IO_CLUSTER
	`define ATCBMC300_MST0_SUPPORT	// Cluster_AXI_MEM0
//	`define ATCBMC300_MST3_SUPPORT  // Cluster_AXI_MEM1
	`define ATCBMC300_MST4_SUPPORT	// Cluster_AXI_MMIO
`else
	`ifdef NDS_IO_BIU_X2
		`define ATCBMC300_MST1_SUPPORT	// Dual BIU IF for i
		`define ATCBMC300_MST2_SUPPORT	// Dual BIU IF for d
	`else
		`define ATCBMC300_MST0_SUPPORT	// Single BIU IF
	`endif
`endif


`ifdef AE350_DMA_SUPPORT
	`define ATCBMC300_MST5_SUPPORT
	`ifdef ATCDMAC300_DUAL_MASTER_IF_SUPPORT
		`define ATCBMC300_MST6_SUPPORT
	`endif // ATCDMAC300_DUAL_MASTER_IF_SUPPORT
`endif
`ifdef AE350_MAC_SUPPORT
	`define ATCBMC300_MST7_SUPPORT
`endif
`ifdef AE350_LCDC_SUPPORT
	`define ATCBMC300_MST8_SUPPORT
`endif

`ifdef NDS_TRACE_TILELINK
	`define ATCBMC300_MST9_SUPPORT
	`define ATCBMC300_SLV6_SUPPORT
`endif


`ifdef PLATFORM_DEBUG_PORT
	`ifdef PLATFORM_PLDM_SYS_BUS_ACCESS
	        `define ATCBMC300_MST10_SUPPORT
	`endif // PLATFORM_PLDM_SYS_BUS_ACCESS
`endif // PLATFORM_DEBUG_PORT

`define ATCBMC300_SLV0_SUPPORT
`define ATCBMC300_SLV1_SUPPORT
`define ATCBMC300_SLV2_SUPPORT
`ifdef NDS_IO_SLAVEPORT_COMMON_X1
	`define ATCBMC300_SLV3_SUPPORT
`endif
`define ATCBMC300_SLV4_SUPPORT
`ifdef NDS_IO_COHERENCE
	`define ATCBMC300_SLV5_SUPPORT
`endif // NDS_IO_COHERENCE

`ifdef NDS_IO_CORE_BRG_ASYNC
	`define ATCBMC300_SLV31_SUPPORT		
`endif // NDS_IO_CORE_BRG_ASYNC

`define ATCBMC300_MST0_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST0_DEFAULT_HIGH_PRIORITY   1
`define ATCBMC300_MST0_OUTSTANDING_DEPTH 32
`define ATCBMC300_MST1_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST1_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST2_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST2_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST3_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST3_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST4_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST4_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST5_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST5_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST6_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST6_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST7_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST7_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST8_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST8_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST9_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST9_OUTSTANDING_DEPTH 8
`define ATCBMC300_MST10_DEFAULT_PRIORITY_RELOAD 1
`define ATCBMC300_MST10_OUTSTANDING_DEPTH 8
//`define ATCBMC300_MST11_OUTSTANDING_DEPTH 4
//`define ATCBMC300_MST12_DEFAULT_PRIORITY_RELOAD 1
//`define ATCBMC300_MST12_OUTSTANDING_DEPTH 4
//`define ATCBMC300_MST13_DEFAULT_PRIORITY_RELOAD 1
//`define ATCBMC300_MST13_OUTSTANDING_DEPTH 4
//`define ATCBMC300_MST14_DEFAULT_PRIORITY_RELOAD 1
//`define ATCBMC300_MST14_OUTSTANDING_DEPTH 4
//`define ATCBMC300_MST15_DEFAULT_PRIORITY_RELOAD 1
//`define ATCBMC300_MST15_OUTSTANDING_DEPTH 4
//-------------------------------------------------
// AXI Slave Base Address
//-------------------------------------------------
`define ATCBMC300_SLV0_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hC0000000
`define ATCBMC300_SLV1_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hE0000000
`define ATCBMC300_SLV2_BASE_ADDR `ATCBMC300_ADDR_WIDTH'h0
`define ATCBMC300_SLV3_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hA0000000
`define ATCBMC300_SLV4_BASE_ADDR `ATCBMC300_ADDR_WIDTH'h80000000
`define ATCBMC300_SLV5_BASE_ADDR `ATCBMC300_ADDR_WIDTH'h0000_0000	//2G - IOCP
`define ATCBMC300_SLV6_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hd000_0000	//256M - Trace Tilelink
//`define ATCBMC300_SLV7_BASE_ADDR `ATCBMC300_ADDR_WIDTH'ha000_0000	//256M
//`define ATCBMC300_SLV8_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hb000_0000	//32M
//`define ATCBMC300_SLV9_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hb200_0000	//32M
//`define ATCBMC300_SLV10_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hb400_0000	//32M
//`define ATCBMC300_SLV11_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hb600_0000	//32M
//`define ATCBMC300_SLV12_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hb800_0000	//32M
//`define ATCBMC300_SLV13_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hba00_0000	//32M
//`define ATCBMC300_SLV14_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbc00_0000	//32M
//`define ATCBMC300_SLV15_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbe00_0000	//8M
//`define ATCBMC300_SLV16_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbe80_0000	//8M
//`define ATCBMC300_SLV17_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbf00_0000	//8M
//`define ATCBMC300_SLV18_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbf80_0000	//4M
//`define ATCBMC300_SLV19_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hbfc0_0000	//4M
//`define ATCBMC300_SLV20_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc030_0000	//1M
//`define ATCBMC300_SLV21_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc040_0000	//4M
//`define ATCBMC300_SLV22_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc080_0000	//8M
//`define ATCBMC300_SLV23_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc100_0000	//16
//`define ATCBMC300_SLV24_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc200_0000	//16
//`define ATCBMC300_SLV25_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc300_0000	//16
//`define ATCBMC300_SLV26_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc400_0000	//32
//`define ATCBMC300_SLV27_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hc800_0000	//32
//`define ATCBMC300_SLV28_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hcc00_0000	//32
//`define ATCBMC300_SLV29_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hd000_0000	//32
//`define ATCBMC300_SLV30_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hd400_0000	//32
`define ATCBMC300_SLV31_BASE_ADDR `ATCBMC300_ADDR_WIDTH'hC0200000

`define ATCBMC300_SLV1_SIZE 10
`define ATCBMC300_SLV2_SIZE 12
`ifdef NDS_IO_HART3
	`define ATCBMC300_SLV3_SIZE 3
`else
`ifdef NDS_IO_HART2
	`define ATCBMC300_SLV3_SIZE 3
`else
`ifdef NDS_IO_HART1
	`define ATCBMC300_SLV3_SIZE 3
`else
	`define ATCBMC300_SLV3_SIZE 3
`endif // NDS_IO_HART1
`endif // NDS_IO_HART2
`endif // NDS_IO_HART3
`define ATCBMC300_SLV4_SIZE 9
`define ATCBMC300_SLV5_SIZE 12
`define ATCBMC300_SLV6_SIZE 9
//`define ATCBMC300_SLV7_SIZE 9
//`define ATCBMC300_SLV8_SIZE 6
//`define ATCBMC300_SLV9_SIZE 6
//`define ATCBMC300_SLV10_SIZE 6
//`define ATCBMC300_SLV11_SIZE 6
//`define ATCBMC300_SLV12_SIZE 6
//`define ATCBMC300_SLV13_SIZE 6
//`define ATCBMC300_SLV14_SIZE 6
//`define ATCBMC300_SLV15_SIZE 4
//`define ATCBMC300_SLV16_SIZE 4
//`define ATCBMC300_SLV17_SIZE 4
//`define ATCBMC300_SLV18_SIZE 3
//`define ATCBMC300_SLV19_SIZE 3
//`define ATCBMC300_SLV20_SIZE 1
//`define ATCBMC300_SLV21_SIZE 3
//`define ATCBMC300_SLV22_SIZE 4
//`define ATCBMC300_SLV23_SIZE 5
//`define ATCBMC300_SLV24_SIZE 5
//`define ATCBMC300_SLV25_SIZE 5
//`define ATCBMC300_SLV26_SIZE 6
//`define ATCBMC300_SLV27_SIZE 6
//`define ATCBMC300_SLV28_SIZE 6
//`define ATCBMC300_SLV29_SIZE 6
//`define ATCBMC300_SLV30_SIZE 6
`define ATCBMC300_SLV31_SIZE 1
`define ATCBMC300_SLV1_FIFO_DEPTH 2
`define ATCBMC300_SLV2_FIFO_DEPTH 8
`define ATCBMC300_SLV3_FIFO_DEPTH 2
`define ATCBMC300_SLV4_FIFO_DEPTH 8
`define ATCBMC300_SLV5_FIFO_DEPTH 4
`define ATCBMC300_SLV6_FIFO_DEPTH 4
//`define ATCBMC300_SLV7_FIFO_DEPTH 4
//`define ATCBMC300_SLV8_FIFO_DEPTH 4
//`define ATCBMC300_SLV9_FIFO_DEPTH 4
//`define ATCBMC300_SLV10_FIFO_DEPTH 4
//`define ATCBMC300_SLV11_FIFO_DEPTH 4
//`define ATCBMC300_SLV12_FIFO_DEPTH 4
//`define ATCBMC300_SLV13_FIFO_DEPTH 4
//`define ATCBMC300_SLV14_FIFO_DEPTH 4
//`define ATCBMC300_SLV15_FIFO_DEPTH 4
//`define ATCBMC300_SLV16_FIFO_DEPTH 4
//`define ATCBMC300_SLV17_FIFO_DEPTH 4
//`define ATCBMC300_SLV18_FIFO_DEPTH 4
//`define ATCBMC300_SLV19_FIFO_DEPTH 4
//`define ATCBMC300_SLV20_FIFO_DEPTH 4
//`define ATCBMC300_SLV21_FIFO_DEPTH 4
//`define ATCBMC300_SLV22_FIFO_DEPTH 4
//`define ATCBMC300_SLV23_FIFO_DEPTH 4
//`define ATCBMC300_SLV24_FIFO_DEPTH 4
//`define ATCBMC300_SLV25_FIFO_DEPTH 4
//`define ATCBMC300_SLV26_FIFO_DEPTH 4
//`define ATCBMC300_SLV27_FIFO_DEPTH 4
//`define ATCBMC300_SLV28_FIFO_DEPTH 4
//`define ATCBMC300_SLV29_FIFO_DEPTH 4
//`define ATCBMC300_SLV30_FIFO_DEPTH 4
`define ATCBMC300_SLV31_FIFO_DEPTH 2

//#VPERL_BEGIN
//#: //-------------------------------------------------
//#: // AXI Master & Slave Ports Connectivity
//#: //-------------------------------------------------
//# for($i = 0; $i < 16; ++$i) {
//#: `ifdef ATCBMC300_MST${i}_SUPPORT
//# for($j = 0; $j < 32; ++$j) {
//#:   %s`define ATCBMC300_MST${i}_SLV${j}	:: ((${j}>4) || (${i}>9))  ? "//" : "";
//# }
//#: `endif // ATCBMC300_MST${i}
//# }
//#VPERL_END

// VPERL_GENERATED_BEGIN
//-------------------------------------------------
// AXI Master & Slave Ports Connectivity
//-------------------------------------------------
`ifdef ATCBMC300_MST0_SUPPORT
  `define ATCBMC300_MST0_SLV0
  `define ATCBMC300_MST0_SLV1
  `define ATCBMC300_MST0_SLV2
  `define ATCBMC300_MST0_SLV3
  `define ATCBMC300_MST0_SLV4
  //`define ATCBMC300_MST0_SLV5
  `define ATCBMC300_MST0_SLV6
  //`define ATCBMC300_MST0_SLV7
  //`define ATCBMC300_MST0_SLV8
  //`define ATCBMC300_MST0_SLV9
  //`define ATCBMC300_MST0_SLV10
  //`define ATCBMC300_MST0_SLV11
  //`define ATCBMC300_MST0_SLV12
  //`define ATCBMC300_MST0_SLV13
  //`define ATCBMC300_MST0_SLV14
  //`define ATCBMC300_MST0_SLV15
  //`define ATCBMC300_MST0_SLV16
  //`define ATCBMC300_MST0_SLV17
  //`define ATCBMC300_MST0_SLV18
  //`define ATCBMC300_MST0_SLV19
  //`define ATCBMC300_MST0_SLV20
  //`define ATCBMC300_MST0_SLV21
  //`define ATCBMC300_MST0_SLV22
  //`define ATCBMC300_MST0_SLV23
  //`define ATCBMC300_MST0_SLV24
  //`define ATCBMC300_MST0_SLV25
  //`define ATCBMC300_MST0_SLV26
  //`define ATCBMC300_MST0_SLV27
  //`define ATCBMC300_MST0_SLV28
  //`define ATCBMC300_MST0_SLV29
  //`define ATCBMC300_MST0_SLV30
  //`define ATCBMC300_MST0_SLV31
`endif // ATCBMC300_MST0
`ifdef ATCBMC300_MST1_SUPPORT
  `define ATCBMC300_MST1_SLV0
  `define ATCBMC300_MST1_SLV1
  `define ATCBMC300_MST1_SLV2
  `define ATCBMC300_MST1_SLV3
  `define ATCBMC300_MST1_SLV4
  //`define ATCBMC300_MST1_SLV5
  `define ATCBMC300_MST1_SLV6
  //`define ATCBMC300_MST1_SLV7
  //`define ATCBMC300_MST1_SLV8
  //`define ATCBMC300_MST1_SLV9
  //`define ATCBMC300_MST1_SLV10
  //`define ATCBMC300_MST1_SLV11
  //`define ATCBMC300_MST1_SLV12
  //`define ATCBMC300_MST1_SLV13
  //`define ATCBMC300_MST1_SLV14
  //`define ATCBMC300_MST1_SLV15
  //`define ATCBMC300_MST1_SLV16
  //`define ATCBMC300_MST1_SLV17
  //`define ATCBMC300_MST1_SLV18
  //`define ATCBMC300_MST1_SLV19
  //`define ATCBMC300_MST1_SLV20
  //`define ATCBMC300_MST1_SLV21
  //`define ATCBMC300_MST1_SLV22
  //`define ATCBMC300_MST1_SLV23
  //`define ATCBMC300_MST1_SLV24
  //`define ATCBMC300_MST1_SLV25
  //`define ATCBMC300_MST1_SLV26
  //`define ATCBMC300_MST1_SLV27
  //`define ATCBMC300_MST1_SLV28
  //`define ATCBMC300_MST1_SLV29
  //`define ATCBMC300_MST1_SLV30
  //`define ATCBMC300_MST1_SLV31
`endif // ATCBMC300_MST1
`ifdef ATCBMC300_MST2_SUPPORT
  `define ATCBMC300_MST2_SLV0
  `define ATCBMC300_MST2_SLV1
  `define ATCBMC300_MST2_SLV2
  `define ATCBMC300_MST2_SLV3
  `define ATCBMC300_MST2_SLV4
  //`define ATCBMC300_MST2_SLV5
  `define ATCBMC300_MST2_SLV6
  //`define ATCBMC300_MST2_SLV7
  //`define ATCBMC300_MST2_SLV8
  //`define ATCBMC300_MST2_SLV9
  //`define ATCBMC300_MST2_SLV10
  //`define ATCBMC300_MST2_SLV11
  //`define ATCBMC300_MST2_SLV12
  //`define ATCBMC300_MST2_SLV13
  //`define ATCBMC300_MST2_SLV14
  //`define ATCBMC300_MST2_SLV15
  //`define ATCBMC300_MST2_SLV16
  //`define ATCBMC300_MST2_SLV17
  //`define ATCBMC300_MST2_SLV18
  //`define ATCBMC300_MST2_SLV19
  //`define ATCBMC300_MST2_SLV20
  //`define ATCBMC300_MST2_SLV21
  //`define ATCBMC300_MST2_SLV22
  //`define ATCBMC300_MST2_SLV23
  //`define ATCBMC300_MST2_SLV24
  //`define ATCBMC300_MST2_SLV25
  //`define ATCBMC300_MST2_SLV26
  //`define ATCBMC300_MST2_SLV27
  //`define ATCBMC300_MST2_SLV28
  //`define ATCBMC300_MST2_SLV29
  //`define ATCBMC300_MST2_SLV30
  //`define ATCBMC300_MST2_SLV31
`endif // ATCBMC300_MST2
`ifdef ATCBMC300_MST3_SUPPORT
  `define ATCBMC300_MST3_SLV0
  `define ATCBMC300_MST3_SLV1
  `define ATCBMC300_MST3_SLV2
  `define ATCBMC300_MST3_SLV3
  `define ATCBMC300_MST3_SLV4
  //`define ATCBMC300_MST3_SLV5
  `define ATCBMC300_MST3_SLV6
  //`define ATCBMC300_MST3_SLV7
  //`define ATCBMC300_MST3_SLV8
  //`define ATCBMC300_MST3_SLV9
  //`define ATCBMC300_MST3_SLV10
  //`define ATCBMC300_MST3_SLV11
  //`define ATCBMC300_MST3_SLV12
  //`define ATCBMC300_MST3_SLV13
  //`define ATCBMC300_MST3_SLV14
  //`define ATCBMC300_MST3_SLV15
  //`define ATCBMC300_MST3_SLV16
  //`define ATCBMC300_MST3_SLV17
  //`define ATCBMC300_MST3_SLV18
  //`define ATCBMC300_MST3_SLV19
  //`define ATCBMC300_MST3_SLV20
  //`define ATCBMC300_MST3_SLV21
  //`define ATCBMC300_MST3_SLV22
  //`define ATCBMC300_MST3_SLV23
  //`define ATCBMC300_MST3_SLV24
  //`define ATCBMC300_MST3_SLV25
  //`define ATCBMC300_MST3_SLV26
  //`define ATCBMC300_MST3_SLV27
  //`define ATCBMC300_MST3_SLV28
  //`define ATCBMC300_MST3_SLV29
  //`define ATCBMC300_MST3_SLV30
  //`define ATCBMC300_MST3_SLV31
`endif // ATCBMC300_MST3
`ifdef ATCBMC300_MST4_SUPPORT
  `define ATCBMC300_MST4_SLV0
  `define ATCBMC300_MST4_SLV1
  `define ATCBMC300_MST4_SLV2
  `define ATCBMC300_MST4_SLV3
  `define ATCBMC300_MST4_SLV4
  //`define ATCBMC300_MST4_SLV5
  `define ATCBMC300_MST4_SLV6
  //`define ATCBMC300_MST4_SLV7
  //`define ATCBMC300_MST4_SLV8
  //`define ATCBMC300_MST4_SLV9
  //`define ATCBMC300_MST4_SLV10
  //`define ATCBMC300_MST4_SLV11
  //`define ATCBMC300_MST4_SLV12
  //`define ATCBMC300_MST4_SLV13
  //`define ATCBMC300_MST4_SLV14
  //`define ATCBMC300_MST4_SLV15
  //`define ATCBMC300_MST4_SLV16
  //`define ATCBMC300_MST4_SLV17
  //`define ATCBMC300_MST4_SLV18
  //`define ATCBMC300_MST4_SLV19
  //`define ATCBMC300_MST4_SLV20
  //`define ATCBMC300_MST4_SLV21
  //`define ATCBMC300_MST4_SLV22
  //`define ATCBMC300_MST4_SLV23
  //`define ATCBMC300_MST4_SLV24
  //`define ATCBMC300_MST4_SLV25
  //`define ATCBMC300_MST4_SLV26
  //`define ATCBMC300_MST4_SLV27
  //`define ATCBMC300_MST4_SLV28
  //`define ATCBMC300_MST4_SLV29
  //`define ATCBMC300_MST4_SLV30

    `ifdef NDS_IO_CORE_BRG_ASYNC
      `define ATCBMC300_MST4_SLV31		
    `endif // NDS_IO_CORE_BRG_ASYNC

`endif // ATCBMC300_MST4
`ifdef ATCBMC300_MST5_SUPPORT
  `define ATCBMC300_MST5_SLV0
  `define ATCBMC300_MST5_SLV1
  `ifndef NDS_IO_COHERENCE
    `define ATCBMC300_MST5_SLV2
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST5_SLV3
  `define ATCBMC300_MST5_SLV4
  `ifdef NDS_IO_COHERENCE
    `define ATCBMC300_MST5_SLV5
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST5_SLV6
  //`define ATCBMC300_MST5_SLV7
  //`define ATCBMC300_MST5_SLV8
  //`define ATCBMC300_MST5_SLV9
  //`define ATCBMC300_MST5_SLV10
  //`define ATCBMC300_MST5_SLV11
  //`define ATCBMC300_MST5_SLV12
  //`define ATCBMC300_MST5_SLV13
  //`define ATCBMC300_MST5_SLV14
  //`define ATCBMC300_MST5_SLV15
  //`define ATCBMC300_MST5_SLV16
  //`define ATCBMC300_MST5_SLV17
  //`define ATCBMC300_MST5_SLV18
  //`define ATCBMC300_MST5_SLV19
  //`define ATCBMC300_MST5_SLV20
  //`define ATCBMC300_MST5_SLV21
  //`define ATCBMC300_MST5_SLV22
  //`define ATCBMC300_MST5_SLV23
  //`define ATCBMC300_MST5_SLV24
  //`define ATCBMC300_MST5_SLV25
  //`define ATCBMC300_MST5_SLV26
  //`define ATCBMC300_MST5_SLV27
  //`define ATCBMC300_MST5_SLV28
  //`define ATCBMC300_MST5_SLV29
  //`define ATCBMC300_MST5_SLV30
  //`define ATCBMC300_MST5_SLV31
`endif // ATCBMC300_MST5
`ifdef ATCBMC300_MST6_SUPPORT
  `define ATCBMC300_MST6_SLV0
  `define ATCBMC300_MST6_SLV1
  `ifndef NDS_IO_COHERENCE
    `define ATCBMC300_MST6_SLV2
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST6_SLV3
  `define ATCBMC300_MST6_SLV4
  `ifdef NDS_IO_COHERENCE
    `define ATCBMC300_MST6_SLV5
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST6_SLV6
  //`define ATCBMC300_MST6_SLV7
  //`define ATCBMC300_MST6_SLV8
  //`define ATCBMC300_MST6_SLV9
  //`define ATCBMC300_MST6_SLV10
  //`define ATCBMC300_MST6_SLV11
  //`define ATCBMC300_MST6_SLV12
  //`define ATCBMC300_MST6_SLV13
  //`define ATCBMC300_MST6_SLV14
  //`define ATCBMC300_MST6_SLV15
  //`define ATCBMC300_MST6_SLV16
  //`define ATCBMC300_MST6_SLV17
  //`define ATCBMC300_MST6_SLV18
  //`define ATCBMC300_MST6_SLV19
  //`define ATCBMC300_MST6_SLV20
  //`define ATCBMC300_MST6_SLV21
  //`define ATCBMC300_MST6_SLV22
  //`define ATCBMC300_MST6_SLV23
  //`define ATCBMC300_MST6_SLV24
  //`define ATCBMC300_MST6_SLV25
  //`define ATCBMC300_MST6_SLV26
  //`define ATCBMC300_MST6_SLV27
  //`define ATCBMC300_MST6_SLV28
  //`define ATCBMC300_MST6_SLV29
  //`define ATCBMC300_MST6_SLV30
  //`define ATCBMC300_MST6_SLV31
`endif // ATCBMC300_MST6
`ifdef ATCBMC300_MST7_SUPPORT
  `define ATCBMC300_MST7_SLV0
  `define ATCBMC300_MST7_SLV1
  `ifndef NDS_IO_COHERENCE
    `define ATCBMC300_MST7_SLV2
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST7_SLV3
  `define ATCBMC300_MST7_SLV4
  `ifdef NDS_IO_COHERENCE
    `define ATCBMC300_MST7_SLV5
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST7_SLV6
  //`define ATCBMC300_MST7_SLV7
  //`define ATCBMC300_MST7_SLV8
  //`define ATCBMC300_MST7_SLV9
  //`define ATCBMC300_MST7_SLV10
  //`define ATCBMC300_MST7_SLV11
  //`define ATCBMC300_MST7_SLV12
  //`define ATCBMC300_MST7_SLV13
  //`define ATCBMC300_MST7_SLV14
  //`define ATCBMC300_MST7_SLV15
  //`define ATCBMC300_MST7_SLV16
  //`define ATCBMC300_MST7_SLV17
  //`define ATCBMC300_MST7_SLV18
  //`define ATCBMC300_MST7_SLV19
  //`define ATCBMC300_MST7_SLV20
  //`define ATCBMC300_MST7_SLV21
  //`define ATCBMC300_MST7_SLV22
  //`define ATCBMC300_MST7_SLV23
  //`define ATCBMC300_MST7_SLV24
  //`define ATCBMC300_MST7_SLV25
  //`define ATCBMC300_MST7_SLV26
  //`define ATCBMC300_MST7_SLV27
  //`define ATCBMC300_MST7_SLV28
  //`define ATCBMC300_MST7_SLV29
  //`define ATCBMC300_MST7_SLV30
  //`define ATCBMC300_MST7_SLV31
`endif // ATCBMC300_MST7
`ifdef ATCBMC300_MST8_SUPPORT
  `define ATCBMC300_MST8_SLV0
  `define ATCBMC300_MST8_SLV1
  `ifndef NDS_IO_COHERENCE
    `define ATCBMC300_MST8_SLV2
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST8_SLV3
  `define ATCBMC300_MST8_SLV4
  `ifdef NDS_IO_COHERENCE
    `define ATCBMC300_MST8_SLV5
  `endif // NDS_IO_COHERENCE
  `define ATCBMC300_MST8_SLV6
  //`define ATCBMC300_MST8_SLV7
  //`define ATCBMC300_MST8_SLV8
  //`define ATCBMC300_MST8_SLV9
  //`define ATCBMC300_MST8_SLV10
  //`define ATCBMC300_MST8_SLV11
  //`define ATCBMC300_MST8_SLV12
  //`define ATCBMC300_MST8_SLV13
  //`define ATCBMC300_MST8_SLV14
  //`define ATCBMC300_MST8_SLV15
  //`define ATCBMC300_MST8_SLV16
  //`define ATCBMC300_MST8_SLV17
  //`define ATCBMC300_MST8_SLV18
  //`define ATCBMC300_MST8_SLV19
  //`define ATCBMC300_MST8_SLV20
  //`define ATCBMC300_MST8_SLV21
  //`define ATCBMC300_MST8_SLV22
  //`define ATCBMC300_MST8_SLV23
  //`define ATCBMC300_MST8_SLV24
  //`define ATCBMC300_MST8_SLV25
  //`define ATCBMC300_MST8_SLV26
  //`define ATCBMC300_MST8_SLV27
  //`define ATCBMC300_MST8_SLV28
  //`define ATCBMC300_MST8_SLV29
  //`define ATCBMC300_MST8_SLV30
  //`define ATCBMC300_MST8_SLV31
`endif // ATCBMC300_MST8
`ifdef ATCBMC300_MST9_SUPPORT
  `define ATCBMC300_MST9_SLV0
  `define ATCBMC300_MST9_SLV1
  `define ATCBMC300_MST9_SLV2
  `define ATCBMC300_MST9_SLV3
  `define ATCBMC300_MST9_SLV4
  //`define ATCBMC300_MST9_SLV5
  `define ATCBMC300_MST9_SLV6
  //`define ATCBMC300_MST9_SLV7
  //`define ATCBMC300_MST9_SLV8
  //`define ATCBMC300_MST9_SLV9
  //`define ATCBMC300_MST9_SLV10
  //`define ATCBMC300_MST9_SLV11
  //`define ATCBMC300_MST9_SLV12
  //`define ATCBMC300_MST9_SLV13
  //`define ATCBMC300_MST9_SLV14
  //`define ATCBMC300_MST9_SLV15
  //`define ATCBMC300_MST9_SLV16
  //`define ATCBMC300_MST9_SLV17
  //`define ATCBMC300_MST9_SLV18
  //`define ATCBMC300_MST9_SLV19
  //`define ATCBMC300_MST9_SLV20
  //`define ATCBMC300_MST9_SLV21
  //`define ATCBMC300_MST9_SLV22
  //`define ATCBMC300_MST9_SLV23
  //`define ATCBMC300_MST9_SLV24
  //`define ATCBMC300_MST9_SLV25
  //`define ATCBMC300_MST9_SLV26
  //`define ATCBMC300_MST9_SLV27
  //`define ATCBMC300_MST9_SLV28
  //`define ATCBMC300_MST9_SLV29
  //`define ATCBMC300_MST9_SLV30
  //`define ATCBMC300_MST9_SLV31
`endif // ATCBMC300_MST9
`ifdef ATCBMC300_MST10_SUPPORT
  `define ATCBMC300_MST10_SLV0
  `define ATCBMC300_MST10_SLV1
  `define ATCBMC300_MST10_SLV2
  `define ATCBMC300_MST10_SLV3
  `define ATCBMC300_MST10_SLV4
  //`define ATCBMC300_MST10_SLV5
  `define ATCBMC300_MST10_SLV6
  //`define ATCBMC300_MST10_SLV7
  //`define ATCBMC300_MST10_SLV8
  //`define ATCBMC300_MST10_SLV9
  //`define ATCBMC300_MST10_SLV10
  //`define ATCBMC300_MST10_SLV11
  //`define ATCBMC300_MST10_SLV12
  //`define ATCBMC300_MST10_SLV13
  //`define ATCBMC300_MST10_SLV14
  //`define ATCBMC300_MST10_SLV15
  //`define ATCBMC300_MST10_SLV16
  //`define ATCBMC300_MST10_SLV17
  //`define ATCBMC300_MST10_SLV18
  //`define ATCBMC300_MST10_SLV19
  //`define ATCBMC300_MST10_SLV20
  //`define ATCBMC300_MST10_SLV21
  //`define ATCBMC300_MST10_SLV22
  //`define ATCBMC300_MST10_SLV23
  //`define ATCBMC300_MST10_SLV24
  //`define ATCBMC300_MST10_SLV25
  //`define ATCBMC300_MST10_SLV26
  //`define ATCBMC300_MST10_SLV27
  //`define ATCBMC300_MST10_SLV28
  //`define ATCBMC300_MST10_SLV29
  //`define ATCBMC300_MST10_SLV30
  //`define ATCBMC300_MST10_SLV31
`endif // ATCBMC300_MST10
`ifdef ATCBMC300_MST11_SUPPORT
  //`define ATCBMC300_MST11_SLV0
  //`define ATCBMC300_MST11_SLV1
  //`define ATCBMC300_MST11_SLV2
  //`define ATCBMC300_MST11_SLV3
  //`define ATCBMC300_MST11_SLV4
  //`define ATCBMC300_MST11_SLV5
  //`define ATCBMC300_MST11_SLV6
  //`define ATCBMC300_MST11_SLV7
  //`define ATCBMC300_MST11_SLV8
  //`define ATCBMC300_MST11_SLV9
  //`define ATCBMC300_MST11_SLV10
  //`define ATCBMC300_MST11_SLV11
  //`define ATCBMC300_MST11_SLV12
  //`define ATCBMC300_MST11_SLV13
  //`define ATCBMC300_MST11_SLV14
  //`define ATCBMC300_MST11_SLV15
  //`define ATCBMC300_MST11_SLV16
  //`define ATCBMC300_MST11_SLV17
  //`define ATCBMC300_MST11_SLV18
  //`define ATCBMC300_MST11_SLV19
  //`define ATCBMC300_MST11_SLV20
  //`define ATCBMC300_MST11_SLV21
  //`define ATCBMC300_MST11_SLV22
  //`define ATCBMC300_MST11_SLV23
  //`define ATCBMC300_MST11_SLV24
  //`define ATCBMC300_MST11_SLV25
  //`define ATCBMC300_MST11_SLV26
  //`define ATCBMC300_MST11_SLV27
  //`define ATCBMC300_MST11_SLV28
  //`define ATCBMC300_MST11_SLV29
  //`define ATCBMC300_MST11_SLV30
  //`define ATCBMC300_MST11_SLV31
`endif // ATCBMC300_MST11
`ifdef ATCBMC300_MST12_SUPPORT
  //`define ATCBMC300_MST12_SLV0
  //`define ATCBMC300_MST12_SLV1
  //`define ATCBMC300_MST12_SLV2
  //`define ATCBMC300_MST12_SLV3
  //`define ATCBMC300_MST12_SLV4
  //`define ATCBMC300_MST12_SLV5
  //`define ATCBMC300_MST12_SLV6
  //`define ATCBMC300_MST12_SLV7
  //`define ATCBMC300_MST12_SLV8
  //`define ATCBMC300_MST12_SLV9
  //`define ATCBMC300_MST12_SLV10
  //`define ATCBMC300_MST12_SLV11
  //`define ATCBMC300_MST12_SLV12
  //`define ATCBMC300_MST12_SLV13
  //`define ATCBMC300_MST12_SLV14
  //`define ATCBMC300_MST12_SLV15
  //`define ATCBMC300_MST12_SLV16
  //`define ATCBMC300_MST12_SLV17
  //`define ATCBMC300_MST12_SLV18
  //`define ATCBMC300_MST12_SLV19
  //`define ATCBMC300_MST12_SLV20
  //`define ATCBMC300_MST12_SLV21
  //`define ATCBMC300_MST12_SLV22
  //`define ATCBMC300_MST12_SLV23
  //`define ATCBMC300_MST12_SLV24
  //`define ATCBMC300_MST12_SLV25
  //`define ATCBMC300_MST12_SLV26
  //`define ATCBMC300_MST12_SLV27
  //`define ATCBMC300_MST12_SLV28
  //`define ATCBMC300_MST12_SLV29
  //`define ATCBMC300_MST12_SLV30
  //`define ATCBMC300_MST12_SLV31
`endif // ATCBMC300_MST12
`ifdef ATCBMC300_MST13_SUPPORT
  //`define ATCBMC300_MST13_SLV0
  //`define ATCBMC300_MST13_SLV1
  //`define ATCBMC300_MST13_SLV2
  //`define ATCBMC300_MST13_SLV3
  //`define ATCBMC300_MST13_SLV4
  //`define ATCBMC300_MST13_SLV5
  //`define ATCBMC300_MST13_SLV6
  //`define ATCBMC300_MST13_SLV7
  //`define ATCBMC300_MST13_SLV8
  //`define ATCBMC300_MST13_SLV9
  //`define ATCBMC300_MST13_SLV10
  //`define ATCBMC300_MST13_SLV11
  //`define ATCBMC300_MST13_SLV12
  //`define ATCBMC300_MST13_SLV13
  //`define ATCBMC300_MST13_SLV14
  //`define ATCBMC300_MST13_SLV15
  //`define ATCBMC300_MST13_SLV16
  //`define ATCBMC300_MST13_SLV17
  //`define ATCBMC300_MST13_SLV18
  //`define ATCBMC300_MST13_SLV19
  //`define ATCBMC300_MST13_SLV20
  //`define ATCBMC300_MST13_SLV21
  //`define ATCBMC300_MST13_SLV22
  //`define ATCBMC300_MST13_SLV23
  //`define ATCBMC300_MST13_SLV24
  //`define ATCBMC300_MST13_SLV25
  //`define ATCBMC300_MST13_SLV26
  //`define ATCBMC300_MST13_SLV27
  //`define ATCBMC300_MST13_SLV28
  //`define ATCBMC300_MST13_SLV29
  //`define ATCBMC300_MST13_SLV30
  //`define ATCBMC300_MST13_SLV31
`endif // ATCBMC300_MST13
`ifdef ATCBMC300_MST14_SUPPORT
  //`define ATCBMC300_MST14_SLV0
  //`define ATCBMC300_MST14_SLV1
  //`define ATCBMC300_MST14_SLV2
  //`define ATCBMC300_MST14_SLV3
  //`define ATCBMC300_MST14_SLV4
  //`define ATCBMC300_MST14_SLV5
  //`define ATCBMC300_MST14_SLV6
  //`define ATCBMC300_MST14_SLV7
  //`define ATCBMC300_MST14_SLV8
  //`define ATCBMC300_MST14_SLV9
  //`define ATCBMC300_MST14_SLV10
  //`define ATCBMC300_MST14_SLV11
  //`define ATCBMC300_MST14_SLV12
  //`define ATCBMC300_MST14_SLV13
  //`define ATCBMC300_MST14_SLV14
  //`define ATCBMC300_MST14_SLV15
  //`define ATCBMC300_MST14_SLV16
  //`define ATCBMC300_MST14_SLV17
  //`define ATCBMC300_MST14_SLV18
  //`define ATCBMC300_MST14_SLV19
  //`define ATCBMC300_MST14_SLV20
  //`define ATCBMC300_MST14_SLV21
  //`define ATCBMC300_MST14_SLV22
  //`define ATCBMC300_MST14_SLV23
  //`define ATCBMC300_MST14_SLV24
  //`define ATCBMC300_MST14_SLV25
  //`define ATCBMC300_MST14_SLV26
  //`define ATCBMC300_MST14_SLV27
  //`define ATCBMC300_MST14_SLV28
  //`define ATCBMC300_MST14_SLV29
  //`define ATCBMC300_MST14_SLV30
  //`define ATCBMC300_MST14_SLV31
`endif // ATCBMC300_MST14
`ifdef ATCBMC300_MST15_SUPPORT
  //`define ATCBMC300_MST15_SLV0
  //`define ATCBMC300_MST15_SLV1
  //`define ATCBMC300_MST15_SLV2
  //`define ATCBMC300_MST15_SLV3
  //`define ATCBMC300_MST15_SLV4
  //`define ATCBMC300_MST15_SLV5
  //`define ATCBMC300_MST15_SLV6
  //`define ATCBMC300_MST15_SLV7
  //`define ATCBMC300_MST15_SLV8
  //`define ATCBMC300_MST15_SLV9
  //`define ATCBMC300_MST15_SLV10
  //`define ATCBMC300_MST15_SLV11
  //`define ATCBMC300_MST15_SLV12
  //`define ATCBMC300_MST15_SLV13
  //`define ATCBMC300_MST15_SLV14
  //`define ATCBMC300_MST15_SLV15
  //`define ATCBMC300_MST15_SLV16
  //`define ATCBMC300_MST15_SLV17
  //`define ATCBMC300_MST15_SLV18
  //`define ATCBMC300_MST15_SLV19
  //`define ATCBMC300_MST15_SLV20
  //`define ATCBMC300_MST15_SLV21
  //`define ATCBMC300_MST15_SLV22
  //`define ATCBMC300_MST15_SLV23
  //`define ATCBMC300_MST15_SLV24
  //`define ATCBMC300_MST15_SLV25
  //`define ATCBMC300_MST15_SLV26
  //`define ATCBMC300_MST15_SLV27
  //`define ATCBMC300_MST15_SLV28
  //`define ATCBMC300_MST15_SLV29
  //`define ATCBMC300_MST15_SLV30
  //`define ATCBMC300_MST15_SLV31
`endif // ATCBMC300_MST15
// VPERL_GENERATED_END


`endif // ATCBMC300_CONFIG_VH


