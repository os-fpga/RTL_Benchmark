module top ( 
    \totalcoeffs[0] , \totalcoeffs[1] , \totalcoeffs[2] , \totalcoeffs[3] ,
    \totalcoeffs[4] , \ctable[0] , \ctable[1] , \ctable[2] ,
    \trailingones[0] , \trailingones[1] ,
    \coeff_token[0] , \coeff_token[1] , \coeff_token[2] , \coeff_token[3] ,
    \coeff_token[4] , \coeff_token[5] , \ctoken_len[0] , \ctoken_len[1] ,
    \ctoken_len[2] , \ctoken_len[3] , \ctoken_len[4]   );
  input  \totalcoeffs[0] , \totalcoeffs[1] , \totalcoeffs[2] ,
    \totalcoeffs[3] , \totalcoeffs[4] , \ctable[0] , \ctable[1] ,
    \ctable[2] , \trailingones[0] , \trailingones[1] ;
  output \coeff_token[0] , \coeff_token[1] , \coeff_token[2] ,
    \coeff_token[3] , \coeff_token[4] , \coeff_token[5] , \ctoken_len[0] ,
    \ctoken_len[1] , \ctoken_len[2] , \ctoken_len[3] , \ctoken_len[4] ;
  wire n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
    n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
    n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n422, n423, n424, n425, n426, n427, n428, n430, n431, n432, n433,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n708, n709, n710, n711, n712, n713;
  assign n22 = ~\totalcoeffs[3]  & ~\ctable[0] ;
  assign n23 = ~\totalcoeffs[1]  & \trailingones[1] ;
  assign n24 = ~\totalcoeffs[0]  & \trailingones[1] ;
  assign n25 = \totalcoeffs[1]  & ~n24;
  assign n26 = ~n23 & ~n25;
  assign n27 = n22 & n26;
  assign n28 = \totalcoeffs[0]  & ~\trailingones[1] ;
  assign n29 = ~\totalcoeffs[1]  & ~n28;
  assign n30 = \totalcoeffs[1]  & ~\trailingones[1] ;
  assign n31 = ~\ctable[2]  & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~\totalcoeffs[2]  & ~n33;
  assign n35 = ~\totalcoeffs[2]  & ~\ctable[0] ;
  assign n36 = ~\totalcoeffs[0]  & ~n35;
  assign n37 = \totalcoeffs[1]  & \totalcoeffs[2] ;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~\trailingones[1]  & ~n38;
  assign n40 = ~\totalcoeffs[2]  & ~\totalcoeffs[3] ;
  assign n41 = \trailingones[1]  & ~n40;
  assign n42 = \totalcoeffs[0]  & \totalcoeffs[3] ;
  assign n43 = ~n41 & ~n42;
  assign n44 = ~\totalcoeffs[1]  & ~n43;
  assign n45 = \totalcoeffs[1]  & ~\totalcoeffs[3] ;
  assign n46 = ~n44 & ~n45;
  assign n47 = ~n39 & n46;
  assign n48 = ~\ctable[2]  & ~n47;
  assign n49 = ~n34 & ~n48;
  assign n50 = ~\trailingones[0]  & ~n49;
  assign n51 = \ctable[2]  & \trailingones[0] ;
  assign n52 = ~\ctable[0]  & n51;
  assign n53 = ~\ctable[2]  & \trailingones[1] ;
  assign n54 = ~n52 & ~n53;
  assign n55 = \totalcoeffs[1]  & ~n54;
  assign n56 = \totalcoeffs[1]  & ~\ctable[2] ;
  assign n57 = ~\ctable[0]  & ~\trailingones[1] ;
  assign n58 = ~n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = \totalcoeffs[0]  & ~\totalcoeffs[2] ;
  assign n61 = ~n59 & n60;
  assign n62 = \totalcoeffs[2]  & ~\trailingones[1] ;
  assign n63 = ~\totalcoeffs[0]  & ~\totalcoeffs[1] ;
  assign n64 = n62 & n63;
  assign n65 = n52 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~\totalcoeffs[3]  & ~n66;
  assign n68 = ~n50 & ~n67;
  assign n69 = ~\ctable[1]  & ~n68;
  assign n70 = ~\totalcoeffs[0]  & ~\totalcoeffs[2] ;
  assign n71 = n23 & n70;
  assign n72 = ~\ctable[0]  & ~n71;
  assign n73 = \ctable[1]  & ~n72;
  assign n74 = ~\totalcoeffs[0]  & ~\trailingones[1] ;
  assign n75 = \totalcoeffs[0]  & \trailingones[1] ;
  assign n76 = ~n74 & ~n75;
  assign n77 = \totalcoeffs[1]  & ~n76;
  assign n78 = \totalcoeffs[2]  & n77;
  assign n79 = \ctable[0]  & n78;
  assign n80 = ~n73 & ~n79;
  assign n81 = \trailingones[0]  & ~n80;
  assign n82 = ~\totalcoeffs[1]  & ~n24;
  assign n83 = ~\trailingones[0]  & ~n82;
  assign n84 = ~\totalcoeffs[1]  & \totalcoeffs[2] ;
  assign n85 = n28 & n84;
  assign n86 = ~n83 & ~n85;
  assign n87 = ~\ctable[0]  & ~n86;
  assign n88 = ~n81 & ~n87;
  assign n89 = \totalcoeffs[3]  & ~n88;
  assign n90 = ~\totalcoeffs[2]  & ~n28;
  assign n91 = \ctable[1]  & ~n90;
  assign n92 = n40 & n77;
  assign n93 = ~n91 & ~n92;
  assign n94 = \ctable[0]  & ~n93;
  assign n95 = \totalcoeffs[2]  & \trailingones[1] ;
  assign n96 = ~\totalcoeffs[2]  & n30;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~\totalcoeffs[0]  & ~\totalcoeffs[3] ;
  assign n99 = ~n97 & n98;
  assign n100 = \ctable[1]  & n99;
  assign n101 = ~n94 & ~n100;
  assign n102 = \trailingones[0]  & ~n101;
  assign n103 = \totalcoeffs[2]  & ~\totalcoeffs[3] ;
  assign n104 = n23 & n103;
  assign n105 = \totalcoeffs[1]  & ~\trailingones[0] ;
  assign n106 = ~n104 & ~n105;
  assign n107 = ~\totalcoeffs[0]  & ~n106;
  assign n108 = ~\totalcoeffs[1]  & ~\trailingones[1] ;
  assign n109 = ~\totalcoeffs[2]  & \ctable[1] ;
  assign n110 = \totalcoeffs[3]  & ~n109;
  assign n111 = n108 & ~n110;
  assign n112 = ~n95 & ~n111;
  assign n113 = ~\trailingones[0]  & ~n112;
  assign n114 = ~n107 & ~n113;
  assign n115 = ~\ctable[0]  & ~n114;
  assign n116 = ~\totalcoeffs[0]  & n40;
  assign n117 = ~\trailingones[0]  & n108;
  assign n118 = n116 & n117;
  assign n119 = ~n115 & ~n118;
  assign n120 = ~n102 & n119;
  assign n121 = ~n89 & n120;
  assign n122 = ~\ctable[2]  & ~n121;
  assign n123 = ~n69 & ~n122;
  assign n124 = ~\totalcoeffs[4]  & ~n123;
  assign n125 = ~\trailingones[0]  & ~\trailingones[1] ;
  assign n126 = ~\ctable[1]  & n125;
  assign n127 = \totalcoeffs[4]  & \trailingones[0] ;
  assign n128 = \ctable[1]  & n127;
  assign n129 = ~n126 & ~n128;
  assign n130 = \ctable[0]  & ~n129;
  assign n131 = \ctable[1]  & ~\trailingones[1] ;
  assign n132 = \totalcoeffs[4]  & \trailingones[1] ;
  assign n133 = ~n131 & ~n132;
  assign n134 = \ctable[0]  & \ctable[1] ;
  assign n135 = ~n133 & ~n134;
  assign n136 = ~\trailingones[0]  & n135;
  assign n137 = ~n130 & ~n136;
  assign n138 = ~\ctable[2]  & ~n137;
  assign n139 = ~\totalcoeffs[1]  & ~\totalcoeffs[3] ;
  assign n140 = ~\totalcoeffs[2]  & n139;
  assign n141 = n138 & n140;
  assign n142 = ~\totalcoeffs[0]  & n141;
  assign \coeff_token[0]  = n124 | n142;
  assign n144 = \totalcoeffs[0]  & \trailingones[0] ;
  assign n145 = n95 & n144;
  assign n146 = ~\totalcoeffs[2]  & ~\trailingones[0] ;
  assign n147 = n74 & n146;
  assign n148 = ~n145 & ~n147;
  assign n149 = \ctable[0]  & ~n148;
  assign n150 = ~\ctable[0]  & \trailingones[0] ;
  assign n151 = \ctable[1]  & \trailingones[1] ;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~\totalcoeffs[0]  & ~n152;
  assign n154 = \trailingones[0]  & n151;
  assign n155 = ~\trailingones[0]  & n57;
  assign n156 = ~n154 & ~n155;
  assign n157 = ~n153 & n156;
  assign n158 = \totalcoeffs[2]  & ~n157;
  assign n159 = ~n149 & ~n158;
  assign n160 = ~\totalcoeffs[4]  & ~n159;
  assign n161 = ~\ctable[1]  & \trailingones[1] ;
  assign n162 = \ctable[0]  & ~\trailingones[0] ;
  assign n163 = ~n127 & ~n162;
  assign n164 = ~\ctable[1]  & ~n163;
  assign n165 = ~n132 & ~n164;
  assign n166 = ~n161 & ~n165;
  assign n167 = n70 & n166;
  assign n168 = ~n160 & ~n167;
  assign n169 = ~\totalcoeffs[1]  & ~n168;
  assign n170 = \ctable[1]  & \trailingones[0] ;
  assign n171 = ~n152 & ~n170;
  assign n172 = \totalcoeffs[0]  & n171;
  assign n173 = ~\totalcoeffs[0]  & \ctable[0] ;
  assign n174 = ~\trailingones[0]  & \trailingones[1] ;
  assign n175 = n173 & n174;
  assign n176 = ~n172 & ~n175;
  assign n177 = ~\totalcoeffs[2]  & ~n176;
  assign n178 = ~\ctable[1]  & ~\trailingones[0] ;
  assign n179 = ~\totalcoeffs[0]  & \ctable[1] ;
  assign n180 = ~\totalcoeffs[2]  & ~n179;
  assign n181 = n150 & ~n180;
  assign n182 = ~n178 & ~n181;
  assign n183 = ~\trailingones[1]  & ~n182;
  assign n184 = ~n177 & ~n183;
  assign n185 = \totalcoeffs[1]  & ~n184;
  assign n186 = ~\ctable[1]  & \trailingones[0] ;
  assign n187 = n62 & n186;
  assign n188 = ~n185 & ~n187;
  assign n189 = ~\totalcoeffs[4]  & ~n188;
  assign n190 = ~n169 & ~n189;
  assign n191 = ~\totalcoeffs[3]  & ~n190;
  assign n192 = \ctable[0]  & n146;
  assign n193 = ~\totalcoeffs[3]  & ~\trailingones[0] ;
  assign n194 = ~n150 & ~n193;
  assign n195 = \totalcoeffs[0]  & n194;
  assign n196 = ~n192 & ~n195;
  assign n197 = ~\totalcoeffs[1]  & ~n196;
  assign n198 = \totalcoeffs[3]  & \trailingones[0] ;
  assign n199 = ~\totalcoeffs[2]  & ~n198;
  assign n200 = ~\totalcoeffs[0]  & ~n199;
  assign n201 = ~\totalcoeffs[2]  & \trailingones[0] ;
  assign n202 = \totalcoeffs[0]  & n201;
  assign n203 = \totalcoeffs[0]  & ~\ctable[0] ;
  assign n204 = ~n173 & ~n203;
  assign n205 = ~n202 & n204;
  assign n206 = \totalcoeffs[1]  & ~n205;
  assign n207 = ~n200 & ~n206;
  assign n208 = ~n197 & n207;
  assign n209 = ~\ctable[1]  & ~n208;
  assign n210 = ~\totalcoeffs[1]  & \ctable[1] ;
  assign n211 = \totalcoeffs[2]  & ~n210;
  assign n212 = ~\totalcoeffs[1]  & ~\trailingones[0] ;
  assign n213 = ~n211 & ~n212;
  assign n214 = \totalcoeffs[3]  & n213;
  assign n215 = ~\totalcoeffs[0]  & \trailingones[0] ;
  assign n216 = ~\totalcoeffs[1]  & ~\ctable[1] ;
  assign n217 = \totalcoeffs[0]  & \totalcoeffs[1] ;
  assign n218 = ~n216 & ~n217;
  assign n219 = ~n215 & n218;
  assign n220 = ~\totalcoeffs[2]  & n219;
  assign n221 = ~n214 & ~n220;
  assign n222 = ~\ctable[0]  & ~n221;
  assign n223 = ~n209 & ~n222;
  assign n224 = ~\trailingones[1]  & ~n223;
  assign n225 = \totalcoeffs[1]  & \ctable[0] ;
  assign n226 = \totalcoeffs[3]  & ~\trailingones[0] ;
  assign n227 = ~\totalcoeffs[1]  & ~\totalcoeffs[2] ;
  assign n228 = n226 & n227;
  assign n229 = ~n225 & ~n228;
  assign n230 = \totalcoeffs[0]  & ~n229;
  assign n231 = \ctable[0]  & ~n40;
  assign n232 = \totalcoeffs[3]  & n37;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n230 & n233;
  assign n235 = \ctable[1]  & ~n234;
  assign n236 = n162 & n232;
  assign n237 = ~n235 & ~n236;
  assign n238 = \trailingones[1]  & ~n237;
  assign n239 = ~n224 & ~n238;
  assign n240 = ~\totalcoeffs[4]  & ~n239;
  assign n241 = ~n191 & ~n240;
  assign n242 = ~\ctable[2]  & ~n241;
  assign n243 = \totalcoeffs[2]  & ~n63;
  assign n244 = n90 & ~n217;
  assign n245 = ~n243 & ~n244;
  assign n246 = ~\trailingones[0]  & n245;
  assign n247 = n30 & n201;
  assign n248 = ~n246 & ~n247;
  assign n249 = \ctable[2]  & ~n248;
  assign n250 = ~n64 & ~n249;
  assign n251 = ~\totalcoeffs[4]  & ~n250;
  assign n252 = ~\ctable[1]  & n251;
  assign n253 = n22 & n252;
  assign \coeff_token[1]  = n242 | n253;
  assign n255 = ~\totalcoeffs[3]  & \trailingones[1] ;
  assign n256 = ~n45 & ~n174;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~\ctable[1]  & n257;
  assign n259 = \totalcoeffs[3]  & ~n201;
  assign n260 = \ctable[0]  & ~n259;
  assign n261 = \totalcoeffs[2]  & ~\ctable[0] ;
  assign n262 = \totalcoeffs[3]  & ~n261;
  assign n263 = \trailingones[0]  & ~n262;
  assign n264 = ~n260 & ~n263;
  assign n265 = \totalcoeffs[1]  & ~n264;
  assign n266 = ~\ctable[0]  & \ctable[1] ;
  assign n267 = ~\trailingones[0]  & n266;
  assign n268 = n139 & n267;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~\trailingones[1]  & ~n269;
  assign n271 = ~\totalcoeffs[1]  & ~n199;
  assign n272 = \totalcoeffs[2]  & ~n186;
  assign n273 = ~n271 & ~n272;
  assign n274 = \ctable[0]  & ~n273;
  assign n275 = \totalcoeffs[1]  & \trailingones[0] ;
  assign n276 = \ctable[1]  & ~n275;
  assign n277 = ~\trailingones[1]  & ~n276;
  assign n278 = ~\totalcoeffs[2]  & ~n277;
  assign n279 = ~\totalcoeffs[1]  & n174;
  assign n280 = ~n278 & ~n279;
  assign n281 = \totalcoeffs[3]  & ~n280;
  assign n282 = \ctable[1]  & ~\trailingones[0] ;
  assign n283 = \totalcoeffs[1]  & n255;
  assign n284 = n282 & n283;
  assign n285 = ~n281 & ~n284;
  assign n286 = ~n274 & n285;
  assign n287 = ~n270 & n286;
  assign n288 = ~n258 & n287;
  assign n289 = ~\totalcoeffs[4]  & ~n288;
  assign n290 = \trailingones[0]  & ~\trailingones[1] ;
  assign n291 = ~n178 & ~n290;
  assign n292 = ~\ctable[0]  & n291;
  assign n293 = ~\totalcoeffs[3]  & \totalcoeffs[4] ;
  assign n294 = ~\totalcoeffs[1]  & n293;
  assign n295 = ~n292 & n294;
  assign n296 = ~\totalcoeffs[2]  & n295;
  assign n297 = ~n289 & ~n296;
  assign n298 = ~\totalcoeffs[0]  & ~n297;
  assign n299 = \trailingones[0]  & n75;
  assign n300 = ~n125 & ~n299;
  assign n301 = \ctable[0]  & ~n300;
  assign n302 = ~\ctable[0]  & n95;
  assign n303 = ~n301 & ~n302;
  assign n304 = \totalcoeffs[1]  & ~n303;
  assign n305 = ~n174 & ~n290;
  assign n306 = ~n108 & n305;
  assign n307 = \totalcoeffs[2]  & ~n306;
  assign n308 = ~n304 & ~n307;
  assign n309 = ~\totalcoeffs[3]  & ~n308;
  assign n310 = ~\totalcoeffs[1]  & \totalcoeffs[3] ;
  assign n311 = \ctable[0]  & ~n310;
  assign n312 = ~\totalcoeffs[2]  & n125;
  assign n313 = ~n311 & n312;
  assign n314 = ~\totalcoeffs[1]  & \trailingones[0] ;
  assign n315 = n41 & n314;
  assign n316 = ~n313 & ~n315;
  assign n317 = \totalcoeffs[0]  & ~n316;
  assign n318 = ~n309 & ~n317;
  assign n319 = ~\ctable[1]  & ~n318;
  assign n320 = \totalcoeffs[1]  & \trailingones[1] ;
  assign n321 = \totalcoeffs[2]  & n320;
  assign n322 = ~n314 & ~n321;
  assign n323 = \ctable[1]  & ~n322;
  assign n324 = \trailingones[0]  & ~n62;
  assign n325 = \totalcoeffs[2]  & n125;
  assign n326 = ~n324 & ~n325;
  assign n327 = ~n323 & n326;
  assign n328 = \totalcoeffs[3]  & ~n327;
  assign n329 = \ctable[1]  & ~n23;
  assign n330 = ~n30 & ~n329;
  assign n331 = \trailingones[0]  & ~n330;
  assign n332 = ~n108 & ~n320;
  assign n333 = n193 & ~n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~\totalcoeffs[2]  & ~n334;
  assign n336 = ~n328 & ~n335;
  assign n337 = n203 & ~n336;
  assign n338 = ~n319 & ~n337;
  assign n339 = ~\totalcoeffs[4]  & ~n338;
  assign n340 = ~n298 & ~n339;
  assign n341 = ~\ctable[2]  & ~n340;
  assign n342 = ~\ctable[0]  & ~\ctable[1] ;
  assign n343 = n51 & n75;
  assign n344 = ~n74 & ~n343;
  assign n345 = \totalcoeffs[1]  & ~n344;
  assign n346 = n28 & n212;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~\totalcoeffs[4]  & ~n347;
  assign n349 = n40 & n348;
  assign n350 = n342 & n349;
  assign \coeff_token[2]  = n341 | n350;
  assign n352 = \totalcoeffs[3]  & ~n161;
  assign n353 = \totalcoeffs[2]  & \ctable[1] ;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~\totalcoeffs[4]  & ~n354;
  assign n356 = \trailingones[0]  & \trailingones[1] ;
  assign n357 = n342 & n356;
  assign n358 = ~n134 & ~n357;
  assign n359 = ~\totalcoeffs[2]  & n293;
  assign n360 = ~n358 & n359;
  assign n361 = ~n355 & ~n360;
  assign n362 = ~\totalcoeffs[1]  & ~n361;
  assign n363 = \ctable[0]  & \trailingones[0] ;
  assign n364 = n161 & n363;
  assign n365 = ~n155 & ~n364;
  assign n366 = \totalcoeffs[2]  & ~n365;
  assign n367 = \ctable[0]  & ~n186;
  assign n368 = \totalcoeffs[3]  & ~n367;
  assign n369 = ~n267 & ~n368;
  assign n370 = ~n366 & n369;
  assign n371 = \totalcoeffs[1]  & ~n370;
  assign n372 = \totalcoeffs[2]  & n266;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~\totalcoeffs[4]  & ~n373;
  assign n375 = ~n362 & ~n374;
  assign n376 = ~\totalcoeffs[0]  & ~n375;
  assign n377 = \totalcoeffs[2]  & ~n194;
  assign n378 = ~\totalcoeffs[2]  & n363;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~\trailingones[1]  & ~n379;
  assign n381 = \ctable[0]  & \trailingones[1] ;
  assign n382 = ~\trailingones[0]  & n381;
  assign n383 = ~\totalcoeffs[3]  & ~n382;
  assign n384 = ~\totalcoeffs[2]  & ~n383;
  assign n385 = ~\ctable[1]  & ~n226;
  assign n386 = \totalcoeffs[3]  & ~\ctable[0] ;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~n384 & ~n387;
  assign n389 = ~n380 & n388;
  assign n390 = \totalcoeffs[1]  & ~n389;
  assign n391 = ~\totalcoeffs[3]  & n266;
  assign n392 = n192 & n216;
  assign n393 = ~n391 & ~n392;
  assign n394 = ~\trailingones[1]  & ~n393;
  assign n395 = ~n390 & ~n394;
  assign n396 = \totalcoeffs[0]  & ~n395;
  assign n397 = ~n40 & n266;
  assign n398 = \totalcoeffs[3]  & ~\ctable[1] ;
  assign n399 = \totalcoeffs[2]  & n398;
  assign n400 = ~n397 & ~n399;
  assign n401 = \trailingones[1]  & ~n400;
  assign n402 = ~\trailingones[1]  & n266;
  assign n403 = ~n398 & ~n402;
  assign n404 = ~\trailingones[0]  & ~n403;
  assign n405 = ~n401 & ~n404;
  assign n406 = ~\totalcoeffs[1]  & ~n405;
  assign n407 = ~n57 & ~n178;
  assign n408 = ~\totalcoeffs[2]  & ~n407;
  assign n409 = ~\ctable[1]  & ~n381;
  assign n410 = ~n320 & ~n363;
  assign n411 = n409 & ~n410;
  assign n412 = ~n408 & ~n411;
  assign n413 = \totalcoeffs[3]  & ~n412;
  assign n414 = \totalcoeffs[1]  & n290;
  assign n415 = n266 & n414;
  assign n416 = ~n413 & ~n415;
  assign n417 = ~n406 & n416;
  assign n418 = ~n396 & n417;
  assign n419 = ~\totalcoeffs[4]  & ~n418;
  assign n420 = ~n376 & ~n419;
  assign \coeff_token[3]  = ~\ctable[2]  & ~n420;
  assign n422 = ~\totalcoeffs[4]  & n243;
  assign n423 = \totalcoeffs[3]  & ~\totalcoeffs[4] ;
  assign n424 = ~n293 & ~n423;
  assign n425 = ~\totalcoeffs[0]  & n227;
  assign n426 = ~n424 & n425;
  assign n427 = ~n422 & ~n426;
  assign n428 = ~\ctable[2]  & ~n427;
  assign \coeff_token[4]  = n134 & n428;
  assign n430 = n63 & n359;
  assign n431 = n423 & ~n425;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~\ctable[2]  & ~n432;
  assign \coeff_token[5]  = n134 & n433;
  assign n435 = ~\totalcoeffs[1]  & ~\ctable[0] ;
  assign n436 = \totalcoeffs[2]  & ~n435;
  assign n437 = ~\trailingones[1]  & ~n436;
  assign n438 = ~\ctable[1]  & n437;
  assign n439 = \ctable[0]  & n320;
  assign n440 = ~n438 & ~n439;
  assign n441 = \totalcoeffs[0]  & ~n440;
  assign n442 = ~\totalcoeffs[0]  & ~n57;
  assign n443 = \totalcoeffs[2]  & n442;
  assign n444 = ~n441 & ~n443;
  assign n445 = \trailingones[0]  & ~n444;
  assign n446 = \totalcoeffs[2]  & n24;
  assign n447 = ~n117 & ~n446;
  assign n448 = \ctable[0]  & ~n447;
  assign n449 = ~n445 & ~n448;
  assign n450 = ~n125 & ~n356;
  assign n451 = \ctable[1]  & ~n450;
  assign n452 = ~\totalcoeffs[2]  & \trailingones[1] ;
  assign n453 = ~n62 & ~n452;
  assign n454 = n451 & n453;
  assign n455 = n449 & ~n454;
  assign n456 = ~\ctable[2]  & ~n455;
  assign n457 = \ctable[2]  & ~\trailingones[1] ;
  assign n458 = \trailingones[0]  & ~n457;
  assign n459 = n84 & ~n458;
  assign n460 = ~n96 & ~n459;
  assign n461 = ~\totalcoeffs[0]  & ~n460;
  assign n462 = n144 & n320;
  assign n463 = ~n125 & ~n462;
  assign n464 = \ctable[2]  & ~n463;
  assign n465 = ~\totalcoeffs[2]  & n464;
  assign n466 = ~n461 & ~n465;
  assign n467 = n342 & ~n466;
  assign n468 = ~n456 & ~n467;
  assign n469 = ~\totalcoeffs[3]  & ~n468;
  assign n470 = ~n117 & ~n320;
  assign n471 = \totalcoeffs[0]  & ~n470;
  assign n472 = \totalcoeffs[2]  & n30;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~\totalcoeffs[0]  & ~\ctable[1] ;
  assign n475 = ~n212 & n332;
  assign n476 = n474 & n475;
  assign n477 = n473 & ~n476;
  assign n478 = ~\ctable[0]  & ~n477;
  assign n479 = ~\trailingones[0]  & n217;
  assign n480 = \totalcoeffs[0]  & n170;
  assign n481 = ~n105 & ~n480;
  assign n482 = ~\totalcoeffs[2]  & ~n481;
  assign n483 = ~n479 & ~n482;
  assign n484 = \trailingones[1]  & ~n483;
  assign n485 = ~\totalcoeffs[0]  & ~\trailingones[0] ;
  assign n486 = ~n203 & ~n485;
  assign n487 = n30 & n486;
  assign n488 = ~n484 & ~n487;
  assign n489 = ~n478 & n488;
  assign n490 = \totalcoeffs[3]  & ~n489;
  assign n491 = ~\totalcoeffs[2]  & \ctable[0] ;
  assign n492 = ~n76 & n491;
  assign n493 = ~\ctable[1]  & ~n261;
  assign n494 = n24 & ~n493;
  assign n495 = ~n492 & ~n494;
  assign n496 = ~\trailingones[0]  & ~n495;
  assign n497 = \totalcoeffs[2]  & ~n125;
  assign n498 = ~n299 & ~n497;
  assign n499 = \ctable[1]  & ~n498;
  assign n500 = ~n496 & ~n499;
  assign n501 = \totalcoeffs[1]  & ~n500;
  assign n502 = ~\trailingones[0]  & ~n474;
  assign n503 = ~n203 & ~n502;
  assign n504 = ~\trailingones[1]  & ~n503;
  assign n505 = ~\totalcoeffs[2]  & n504;
  assign n506 = \totalcoeffs[2]  & \trailingones[0] ;
  assign n507 = n24 & n506;
  assign n508 = ~n505 & ~n507;
  assign n509 = ~\totalcoeffs[1]  & ~n508;
  assign n510 = ~n501 & ~n509;
  assign n511 = ~n490 & n510;
  assign n512 = ~\ctable[2]  & ~n511;
  assign n513 = ~n469 & ~n512;
  assign n514 = ~\totalcoeffs[4]  & ~n513;
  assign n515 = ~\totalcoeffs[1]  & \totalcoeffs[4] ;
  assign n516 = n116 & n515;
  assign n517 = ~n134 & ~n516;
  assign n518 = ~\ctable[2]  & ~n517;
  assign \ctoken_len[0]  = ~n514 & ~n518;
  assign n520 = ~\totalcoeffs[3]  & \trailingones[0] ;
  assign n521 = ~n151 & ~n520;
  assign n522 = \totalcoeffs[0]  & ~n521;
  assign n523 = n215 & n398;
  assign n524 = ~n282 & ~n523;
  assign n525 = \trailingones[1]  & ~n524;
  assign n526 = ~\trailingones[1]  & n170;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~n522 & n527;
  assign n529 = ~\totalcoeffs[2]  & ~n528;
  assign n530 = ~\totalcoeffs[3]  & n356;
  assign n531 = \totalcoeffs[3]  & ~n356;
  assign n532 = ~n144 & ~n531;
  assign n533 = ~\ctable[1]  & ~n532;
  assign n534 = ~n530 & ~n533;
  assign n535 = \totalcoeffs[2]  & ~n534;
  assign n536 = ~\totalcoeffs[3]  & n126;
  assign n537 = ~n535 & ~n536;
  assign n538 = ~n529 & n537;
  assign n539 = \totalcoeffs[1]  & ~n538;
  assign n540 = ~n74 & ~n174;
  assign n541 = ~\ctable[1]  & ~n540;
  assign n542 = ~\totalcoeffs[2]  & n541;
  assign n543 = ~\totalcoeffs[0]  & n451;
  assign n544 = ~n542 & ~n543;
  assign n545 = \totalcoeffs[3]  & ~n544;
  assign n546 = ~\totalcoeffs[0]  & n146;
  assign n547 = ~n480 & ~n546;
  assign n548 = ~\trailingones[1]  & ~n547;
  assign n549 = ~\ctable[1]  & ~n193;
  assign n550 = n497 & ~n549;
  assign n551 = ~n548 & ~n550;
  assign n552 = ~n545 & n551;
  assign n553 = ~\totalcoeffs[1]  & ~n552;
  assign n554 = ~\totalcoeffs[2]  & \totalcoeffs[3] ;
  assign n555 = ~\trailingones[1]  & n282;
  assign n556 = n554 & n555;
  assign n557 = ~n553 & ~n556;
  assign n558 = ~n539 & n557;
  assign n559 = ~\ctable[0]  & ~n558;
  assign n560 = \totalcoeffs[0]  & ~n453;
  assign n561 = \ctable[0]  & ~\trailingones[1] ;
  assign n562 = ~\totalcoeffs[0]  & n561;
  assign n563 = ~n560 & ~n562;
  assign n564 = \trailingones[0]  & ~n563;
  assign n565 = n95 & n162;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~\totalcoeffs[3]  & ~n566;
  assign n568 = \totalcoeffs[3]  & \ctable[0] ;
  assign n569 = ~n62 & ~n568;
  assign n570 = ~\totalcoeffs[0]  & ~n569;
  assign n571 = \totalcoeffs[3]  & n491;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~\trailingones[0]  & ~n572;
  assign n574 = n554 & n561;
  assign n575 = ~n573 & ~n574;
  assign n576 = ~n567 & n575;
  assign n577 = \totalcoeffs[1]  & ~n576;
  assign n578 = \totalcoeffs[2]  & \totalcoeffs[3] ;
  assign n579 = ~\totalcoeffs[2]  & ~n42;
  assign n580 = ~n450 & ~n579;
  assign n581 = ~n578 & ~n580;
  assign n582 = \ctable[0]  & ~n581;
  assign n583 = n42 & n325;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~\totalcoeffs[1]  & ~n584;
  assign n586 = \trailingones[0]  & n381;
  assign n587 = n578 & n586;
  assign n588 = ~n585 & ~n587;
  assign n589 = ~n577 & n588;
  assign n590 = ~\ctable[1]  & ~n589;
  assign n591 = ~n559 & ~n590;
  assign n592 = ~\ctable[2]  & ~n591;
  assign n593 = \totalcoeffs[2]  & ~n305;
  assign n594 = ~\totalcoeffs[0]  & n593;
  assign n595 = ~\trailingones[1]  & n51;
  assign n596 = n60 & n595;
  assign n597 = ~n594 & ~n596;
  assign n598 = n216 & ~n597;
  assign n599 = n22 & n598;
  assign n600 = ~n592 & ~n599;
  assign n601 = ~\totalcoeffs[4]  & ~n600;
  assign n602 = n35 & n98;
  assign n603 = \totalcoeffs[4]  & ~\ctable[2] ;
  assign n604 = n216 & n603;
  assign n605 = n602 & n604;
  assign \ctoken_len[1]  = ~n601 & ~n605;
  assign n607 = n227 & n561;
  assign n608 = ~n283 & ~n607;
  assign n609 = ~\totalcoeffs[0]  & ~n608;
  assign n610 = ~\totalcoeffs[1]  & \ctable[0] ;
  assign n611 = ~n22 & ~n610;
  assign n612 = ~n108 & ~n255;
  assign n613 = ~n611 & n612;
  assign n614 = ~\totalcoeffs[2]  & n613;
  assign n615 = n332 & ~n435;
  assign n616 = n103 & ~n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = ~n609 & n617;
  assign n619 = ~\trailingones[0]  & ~n618;
  assign n620 = ~n98 & ~n611;
  assign n621 = ~\totalcoeffs[2]  & n620;
  assign n622 = n139 & n203;
  assign n623 = ~n621 & ~n622;
  assign n624 = \trailingones[0]  & ~n623;
  assign n625 = ~\ctable[0]  & ~n215;
  assign n626 = ~n568 & ~n625;
  assign n627 = n37 & n626;
  assign n628 = ~n624 & ~n627;
  assign n629 = ~\trailingones[1]  & ~n628;
  assign n630 = ~n261 & ~n568;
  assign n631 = ~n259 & ~n630;
  assign n632 = \totalcoeffs[1]  & n631;
  assign n633 = ~n173 & n310;
  assign n634 = n201 & n633;
  assign n635 = ~n632 & ~n634;
  assign n636 = \trailingones[1]  & ~n635;
  assign n637 = ~n629 & ~n636;
  assign n638 = ~n619 & n637;
  assign n639 = ~\ctable[1]  & ~n638;
  assign n640 = ~\totalcoeffs[1]  & ~n125;
  assign n641 = \totalcoeffs[2]  & ~n640;
  assign n642 = ~n329 & ~n641;
  assign n643 = \totalcoeffs[0]  & ~n642;
  assign n644 = ~\ctable[1]  & ~n105;
  assign n645 = \totalcoeffs[2]  & ~n644;
  assign n646 = \trailingones[0]  & ~n30;
  assign n647 = n329 & ~n646;
  assign n648 = ~n645 & ~n647;
  assign n649 = ~n643 & n648;
  assign n650 = n386 & ~n649;
  assign n651 = ~n639 & ~n650;
  assign n652 = ~\ctable[2]  & ~n651;
  assign n653 = ~n146 & ~n506;
  assign n654 = ~\totalcoeffs[0]  & ~n653;
  assign n655 = ~n202 & ~n654;
  assign n656 = ~\trailingones[1]  & ~n655;
  assign n657 = n95 & n485;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~\totalcoeffs[1]  & ~n658;
  assign n660 = n320 & n546;
  assign n661 = ~n659 & ~n660;
  assign n662 = n22 & ~n661;
  assign n663 = ~\ctable[1]  & n662;
  assign n664 = ~n652 & ~n663;
  assign n665 = ~\totalcoeffs[4]  & ~n664;
  assign n666 = n22 & n603;
  assign n667 = n425 & n666;
  assign \ctoken_len[2]  = ~n665 & ~n667;
  assign n669 = \totalcoeffs[4]  & ~n140;
  assign n670 = n203 & n399;
  assign n671 = ~\ctable[2]  & ~n670;
  assign n672 = ~n640 & ~n671;
  assign n673 = ~\ctable[2]  & ~n140;
  assign n674 = \totalcoeffs[0]  & ~n673;
  assign n675 = \ctable[2]  & ~n103;
  assign n676 = ~\totalcoeffs[3]  & ~n57;
  assign n677 = \totalcoeffs[3]  & ~n151;
  assign n678 = n215 & ~n677;
  assign n679 = ~n676 & ~n678;
  assign n680 = ~\totalcoeffs[2]  & ~n679;
  assign n681 = ~n356 & n399;
  assign n682 = ~\ctable[0]  & n681;
  assign n683 = ~\ctable[1]  & ~n586;
  assign n684 = ~\totalcoeffs[3]  & ~n683;
  assign n685 = ~n682 & ~n684;
  assign n686 = ~n680 & n685;
  assign n687 = \totalcoeffs[1]  & ~n686;
  assign n688 = n215 & ~n409;
  assign n689 = ~n151 & ~n688;
  assign n690 = \totalcoeffs[3]  & ~n689;
  assign n691 = \totalcoeffs[4]  & ~n342;
  assign n692 = ~\totalcoeffs[3]  & ~n691;
  assign n693 = ~n690 & ~n692;
  assign n694 = ~\totalcoeffs[2]  & ~n693;
  assign n695 = ~\trailingones[0]  & ~n381;
  assign n696 = n676 & ~n695;
  assign n697 = \totalcoeffs[2]  & n696;
  assign n698 = ~n694 & ~n697;
  assign n699 = ~\totalcoeffs[1]  & ~n698;
  assign n700 = ~\ctable[0]  & ~n103;
  assign n701 = \ctable[1]  & ~n700;
  assign n702 = ~n699 & ~n701;
  assign n703 = ~n687 & n702;
  assign n704 = ~n675 & n703;
  assign n705 = ~n674 & n704;
  assign n706 = ~n672 & n705;
  assign \ctoken_len[3]  = ~n669 & n706;
  assign n708 = ~\trailingones[0]  & ~n29;
  assign n709 = ~n25 & ~n708;
  assign n710 = n423 & ~n709;
  assign n711 = \totalcoeffs[2]  & n710;
  assign n712 = ~n430 & ~n711;
  assign n713 = ~\ctable[2]  & ~n712;
  assign \ctoken_len[4]  = n342 & n713;
endmodule

