//------------------------------------------------------------------------
// Filename     : ae350p_config.inc
// Description  : Add for peripheral IP configurations
//------------------------------------------------------------------------
`ifdef AE350_CONFIG_VH
`else
`define AE350_CONFIG_VH

// `define AE350_GPIO_SUPPORT
// `define AE350_DMA_SUPPORT
`define	AE350_SPI1_SUPPORT
// `define	AE350_SPI2_SUPPORT
// `define	AE350_I2C_SUPPORT
// `define	AE350_UART1_SUPPORT
// `define	AE350_UART2_SUPPORT
// `define AE350_PIT_SUPPORT
// `define AE350_WDT_SUPPORT
// `define AE350_RTC_SUPPORT

//------------------------------------------------------------------------
// Debug configs
//------------------------------------------------------------------------
// Generated by config tool
//`define PLATFORM_NO_DEBUG_SUPPORT
//
//--- minor configurations
//`define PLATFORM_JTAG_TWOWIRE
`define PLATFORM_PLDM_SYS_BUS_ACCESS
`define PLATFORM_PLDM_PROGBUF_SIZE      8
`define PLATFORM_PLDM_HALTGROUP_COUNT   0
 `define PLATFORM_VECTOR_PLIC_SUPPORT
//------------------------------------------------------------------------
// Unconfigurable
//------------------------------------------------------------------------
`define AE350_AXI_SUPPORT

`ifndef PLATFORM_NO_DEBUG_SUPPORT
`define PLATFORM_DEBUG_PORT
`define PLATFORM_DEBUG_SUBSYSTEM
`endif // PLATFORM_NO_DEBUG_SUPPORT

`define PLATFORM_RESET_VECTOR 64'h0000000080000000
`define PLATFORM_PLDM_REGS_BASE 64'h00000000E6800000
`define PLATFORM_DEBUG_VECTOR 64'h00000000E6800000
`define PLATFORM_SLVPORT_DLM_SEL_BIT 21
`define PLATFORM_SPI_MEM_BASE 64'h0000000080000000
`endif //AE350_CONFIG_VH
