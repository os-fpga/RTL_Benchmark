library ieee;
use ieee.std_logic_1164.all;

entity top is
port( a, b: in std_logic_vector(63 downto 0);
f: out std_logic_vector(127 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061: std_logic;

begin

w0 <= a(0) and b(0);
w1 <= a(2) and not w0;
w2 <= not a(2) and not w0;
w3 <= not w1 and not w2;
w4 <= not a(0) and a(1);
w5 <= b(0) and w4;
w6 <= not a(1) and a(2);
w7 <= a(1) and not a(2);
w8 <= not w6 and not w7;
w9 <= a(0) and w8;
w10 <= b(1) and w9;
w11 <= not w5 and not w10;
w12 <= a(0) and not w8;
w13 <= b(0) and not b(1);
w14 <= not b(0) and b(1);
w15 <= not w13 and not w14;
w16 <= w12 and not w15;
w17 <= w11 and not w16;
w18 <= a(2) and not w17;
w19 <= a(2) and not w18;
w20 <= not w17 and not w18;
w21 <= not w19 and not w20;
w22 <= w1 and not w21;
w23 <= not w1 and w21;
w24 <= not w22 and not w23;
w25 <= b(2) and w9;
w26 <= not a(0) and not w8;
w27 <= not a(1) and w26;
w28 <= b(0) and w27;
w29 <= b(1) and w4;
w30 <= not w28 and not w29;
w31 <= not w25 and w30;
w32 <= b(0) and not b(2);
w33 <= b(1) and w32;
w34 <= b(1) and not b(2);
w35 <= not b(1) and b(2);
w36 <= not w34 and not w35;
w37 <= b(0) and b(1);
w38 <= w36 and not w37;
w39 <= not w33 and not w38;
w40 <= w12 and w39;
w41 <= w31 and not w40;
w42 <= a(2) and not w41;
w43 <= a(2) and not w42;
w44 <= not w41 and not w42;
w45 <= not w43 and not w44;
w46 <= w22 and not w45;
w47 <= not w22 and w45;
w48 <= not w46 and not w47;
w49 <= b(3) and w9;
w50 <= b(1) and w27;
w51 <= b(2) and w4;
w52 <= not w50 and not w51;
w53 <= not w49 and w52;
w54 <= b(1) and b(2);
w55 <= not w33 and not w54;
w56 <= not b(2) and not b(3);
w57 <= b(2) and b(3);
w58 <= not w56 and not w57;
w59 <= not w55 and w58;
w60 <= w55 and not w58;
w61 <= not w59 and not w60;
w62 <= w12 and w61;
w63 <= w53 and not w62;
w64 <= a(2) and not w63;
w65 <= a(2) and not w64;
w66 <= not w63 and not w64;
w67 <= not w65 and not w66;
w68 <= a(2) and not a(3);
w69 <= not a(2) and a(3);
w70 <= not w68 and not w69;
w71 <= b(0) and not w70;
w72 <= not w67 and w71;
w73 <= w67 and not w71;
w74 <= not w72 and not w73;
w75 <= w46 and w74;
w76 <= not w46 and not w74;
w77 <= not w75 and not w76;
w78 <= b(4) and w9;
w79 <= b(2) and w27;
w80 <= b(3) and w4;
w81 <= not w79 and not w80;
w82 <= not w78 and w81;
w83 <= not w57 and not w59;
w84 <= not b(3) and not b(4);
w85 <= b(3) and b(4);
w86 <= not w84 and not w85;
w87 <= not w83 and w86;
w88 <= w83 and not w86;
w89 <= not w87 and not w88;
w90 <= w12 and w89;
w91 <= w82 and not w90;
w92 <= a(2) and not w91;
w93 <= a(2) and not w92;
w94 <= not w91 and not w92;
w95 <= not w93 and not w94;
w96 <= a(5) and not w71;
w97 <= not a(3) and a(4);
w98 <= a(3) and not a(4);
w99 <= not w97 and not w98;
w100 <= w70 and not w99;
w101 <= b(0) and w100;
w102 <= not a(4) and a(5);
w103 <= a(4) and not a(5);
w104 <= not w102 and not w103;
w105 <= not w70 and w104;
w106 <= b(1) and w105;
w107 <= not w101 and not w106;
w108 <= not w70 and not w104;
w109 <= not w15 and w108;
w110 <= w107 and not w109;
w111 <= a(5) and not w110;
w112 <= a(5) and not w111;
w113 <= not w110 and not w111;
w114 <= not w112 and not w113;
w115 <= w96 and not w114;
w116 <= not w96 and w114;
w117 <= not w115 and not w116;
w118 <= not w95 and w117;
w119 <= w117 and not w118;
w120 <= not w95 and not w118;
w121 <= not w119 and not w120;
w122 <= not w72 and not w75;
w123 <= not w121 and not w122;
w124 <= w121 and w122;
w125 <= not w123 and not w124;
w126 <= b(5) and w9;
w127 <= b(3) and w27;
w128 <= b(4) and w4;
w129 <= not w127 and not w128;
w130 <= not w126 and w129;
w131 <= not w85 and not w87;
w132 <= not b(4) and not b(5);
w133 <= b(4) and b(5);
w134 <= not w132 and not w133;
w135 <= not w131 and w134;
w136 <= w131 and not w134;
w137 <= not w135 and not w136;
w138 <= w12 and w137;
w139 <= w130 and not w138;
w140 <= a(2) and not w139;
w141 <= a(2) and not w140;
w142 <= not w139 and not w140;
w143 <= not w141 and not w142;
w144 <= b(2) and w105;
w145 <= w70 and not w104;
w146 <= w99 and w145;
w147 <= b(0) and w146;
w148 <= b(1) and w100;
w149 <= not w147 and not w148;
w150 <= not w144 and w149;
w151 <= not w108 and w150;
w152 <= not w39 and w150;
w153 <= not w151 and not w152;
w154 <= a(5) and not w153;
w155 <= not a(5) and w153;
w156 <= not w154 and not w155;
w157 <= w115 and not w156;
w158 <= not w115 and w156;
w159 <= not w157 and not w158;
w160 <= not w143 and w159;
w161 <= w159 and not w160;
w162 <= not w143 and not w160;
w163 <= not w161 and not w162;
w164 <= not w118 and not w123;
w165 <= not w163 and not w164;
w166 <= w163 and w164;
w167 <= not w165 and not w166;
w168 <= not w160 and not w165;
w169 <= a(5) and not a(6);
w170 <= not a(5) and a(6);
w171 <= not w169 and not w170;
w172 <= b(0) and not w171;
w173 <= w157 and w172;
w174 <= w157 and not w173;
w175 <= w172 and not w173;
w176 <= not w174 and not w175;
w177 <= b(3) and w105;
w178 <= b(1) and w146;
w179 <= b(2) and w100;
w180 <= not w178 and not w179;
w181 <= not w177 and w180;
w182 <= w61 and w108;
w183 <= w181 and not w182;
w184 <= a(5) and not w183;
w185 <= a(5) and not w184;
w186 <= not w183 and not w184;
w187 <= not w185 and not w186;
w188 <= not w176 and w187;
w189 <= w176 and not w187;
w190 <= not w188 and not w189;
w191 <= b(6) and w9;
w192 <= b(4) and w27;
w193 <= b(5) and w4;
w194 <= not w192 and not w193;
w195 <= not w191 and w194;
w196 <= not w133 and not w135;
w197 <= not b(5) and not b(6);
w198 <= b(5) and b(6);
w199 <= not w197 and not w198;
w200 <= not w196 and w199;
w201 <= w196 and not w199;
w202 <= not w200 and not w201;
w203 <= w12 and w202;
w204 <= w195 and not w203;
w205 <= a(2) and not w204;
w206 <= a(2) and not w205;
w207 <= not w204 and not w205;
w208 <= not w206 and not w207;
w209 <= not w190 and not w208;
w210 <= w190 and w208;
w211 <= not w209 and not w210;
w212 <= not w168 and w211;
w213 <= w168 and not w211;
w214 <= not w212 and not w213;
w215 <= not w209 and not w212;
w216 <= b(7) and w9;
w217 <= b(5) and w27;
w218 <= b(6) and w4;
w219 <= not w217 and not w218;
w220 <= not w216 and w219;
w221 <= not w198 and not w200;
w222 <= not b(6) and not b(7);
w223 <= b(6) and b(7);
w224 <= not w222 and not w223;
w225 <= not w221 and w224;
w226 <= w221 and not w224;
w227 <= not w225 and not w226;
w228 <= w12 and w227;
w229 <= w220 and not w228;
w230 <= a(2) and not w229;
w231 <= a(2) and not w230;
w232 <= not w229 and not w230;
w233 <= not w231 and not w232;
w234 <= b(4) and w105;
w235 <= b(2) and w146;
w236 <= b(3) and w100;
w237 <= not w235 and not w236;
w238 <= not w234 and w237;
w239 <= w89 and w108;
w240 <= w238 and not w239;
w241 <= a(5) and not w240;
w242 <= a(5) and not w241;
w243 <= not w240 and not w241;
w244 <= not w242 and not w243;
w245 <= a(8) and not w172;
w246 <= not a(6) and a(7);
w247 <= a(6) and not a(7);
w248 <= not w246 and not w247;
w249 <= w171 and not w248;
w250 <= b(0) and w249;
w251 <= not a(7) and a(8);
w252 <= a(7) and not a(8);
w253 <= not w251 and not w252;
w254 <= not w171 and w253;
w255 <= b(1) and w254;
w256 <= not w250 and not w255;
w257 <= not w171 and not w253;
w258 <= not w15 and w257;
w259 <= w256 and not w258;
w260 <= a(8) and not w259;
w261 <= a(8) and not w260;
w262 <= not w259 and not w260;
w263 <= not w261 and not w262;
w264 <= w245 and not w263;
w265 <= not w245 and w263;
w266 <= not w264 and not w265;
w267 <= not w244 and w266;
w268 <= w266 and not w267;
w269 <= not w244 and not w267;
w270 <= not w268 and not w269;
w271 <= not w176 and not w187;
w272 <= not w173 and not w271;
w273 <= not w270 and not w272;
w274 <= w270 and w272;
w275 <= not w273 and not w274;
w276 <= not w233 and w275;
w277 <= w233 and not w275;
w278 <= not w276 and not w277;
w279 <= not w215 and w278;
w280 <= w215 and not w278;
w281 <= not w279 and not w280;
w282 <= b(2) and w254;
w283 <= w171 and not w253;
w284 <= w248 and w283;
w285 <= b(0) and w284;
w286 <= b(1) and w249;
w287 <= not w285 and not w286;
w288 <= not w282 and w287;
w289 <= w39 and w257;
w290 <= w288 and not w289;
w291 <= a(8) and not w290;
w292 <= a(8) and not w291;
w293 <= not w290 and not w291;
w294 <= not w292 and not w293;
w295 <= not w264 and w294;
w296 <= w264 and not w294;
w297 <= not w295 and not w296;
w298 <= b(5) and w105;
w299 <= b(3) and w146;
w300 <= b(4) and w100;
w301 <= not w299 and not w300;
w302 <= not w298 and w301;
w303 <= w108 and w137;
w304 <= w302 and not w303;
w305 <= a(5) and not w304;
w306 <= a(5) and not w305;
w307 <= not w304 and not w305;
w308 <= not w306 and not w307;
w309 <= w297 and not w308;
w310 <= w297 and not w309;
w311 <= not w308 and not w309;
w312 <= not w310 and not w311;
w313 <= not w267 and not w273;
w314 <= w312 and w313;
w315 <= not w312 and not w313;
w316 <= not w314 and not w315;
w317 <= b(8) and w9;
w318 <= b(6) and w27;
w319 <= b(7) and w4;
w320 <= not w318 and not w319;
w321 <= not w317 and w320;
w322 <= not w223 and not w225;
w323 <= not b(7) and not b(8);
w324 <= b(7) and b(8);
w325 <= not w323 and not w324;
w326 <= not w322 and w325;
w327 <= w322 and not w325;
w328 <= not w326 and not w327;
w329 <= w12 and w328;
w330 <= w321 and not w329;
w331 <= a(2) and not w330;
w332 <= a(2) and not w331;
w333 <= not w330 and not w331;
w334 <= not w332 and not w333;
w335 <= w316 and not w334;
w336 <= w316 and not w335;
w337 <= not w334 and not w335;
w338 <= not w336 and not w337;
w339 <= not w276 and not w279;
w340 <= not w338 and not w339;
w341 <= w338 and w339;
w342 <= not w340 and not w341;
w343 <= b(6) and w105;
w344 <= b(4) and w146;
w345 <= b(5) and w100;
w346 <= not w344 and not w345;
w347 <= not w343 and w346;
w348 <= w108 and w202;
w349 <= w347 and not w348;
w350 <= a(5) and not w349;
w351 <= a(5) and not w350;
w352 <= not w349 and not w350;
w353 <= not w351 and not w352;
w354 <= a(8) and not a(9);
w355 <= not a(8) and a(9);
w356 <= not w354 and not w355;
w357 <= b(0) and not w356;
w358 <= not w296 and w357;
w359 <= w296 and not w357;
w360 <= not w358 and not w359;
w361 <= b(3) and w254;
w362 <= b(1) and w284;
w363 <= b(2) and w249;
w364 <= not w362 and not w363;
w365 <= not w361 and w364;
w366 <= w61 and w257;
w367 <= w365 and not w366;
w368 <= a(8) and not w367;
w369 <= a(8) and not w368;
w370 <= not w367 and not w368;
w371 <= not w369 and not w370;
w372 <= not w360 and not w371;
w373 <= w360 and w371;
w374 <= not w372 and not w373;
w375 <= not w353 and w374;
w376 <= w374 and not w375;
w377 <= not w353 and not w375;
w378 <= not w376 and not w377;
w379 <= not w309 and not w315;
w380 <= w378 and w379;
w381 <= not w378 and not w379;
w382 <= not w380 and not w381;
w383 <= b(9) and w9;
w384 <= b(7) and w27;
w385 <= b(8) and w4;
w386 <= not w384 and not w385;
w387 <= not w383 and w386;
w388 <= not w324 and not w326;
w389 <= not b(8) and not b(9);
w390 <= b(8) and b(9);
w391 <= not w389 and not w390;
w392 <= not w388 and w391;
w393 <= w388 and not w391;
w394 <= not w392 and not w393;
w395 <= w12 and w394;
w396 <= w387 and not w395;
w397 <= a(2) and not w396;
w398 <= a(2) and not w397;
w399 <= not w396 and not w397;
w400 <= not w398 and not w399;
w401 <= w382 and not w400;
w402 <= w382 and not w401;
w403 <= not w400 and not w401;
w404 <= not w402 and not w403;
w405 <= not w335 and not w340;
w406 <= not w404 and not w405;
w407 <= w404 and w405;
w408 <= not w406 and not w407;
w409 <= not w401 and not w406;
w410 <= b(7) and w105;
w411 <= b(5) and w146;
w412 <= b(6) and w100;
w413 <= not w411 and not w412;
w414 <= not w410 and w413;
w415 <= w108 and w227;
w416 <= w414 and not w415;
w417 <= a(5) and not w416;
w418 <= a(5) and not w417;
w419 <= not w416 and not w417;
w420 <= not w418 and not w419;
w421 <= w296 and w357;
w422 <= not w372 and not w421;
w423 <= b(4) and w254;
w424 <= b(2) and w284;
w425 <= b(3) and w249;
w426 <= not w424 and not w425;
w427 <= not w423 and w426;
w428 <= w89 and w257;
w429 <= w427 and not w428;
w430 <= a(8) and not w429;
w431 <= a(8) and not w430;
w432 <= not w429 and not w430;
w433 <= not w431 and not w432;
w434 <= a(11) and not w357;
w435 <= not a(9) and a(10);
w436 <= a(9) and not a(10);
w437 <= not w435 and not w436;
w438 <= w356 and not w437;
w439 <= b(0) and w438;
w440 <= not a(10) and a(11);
w441 <= a(10) and not a(11);
w442 <= not w440 and not w441;
w443 <= not w356 and w442;
w444 <= b(1) and w443;
w445 <= not w439 and not w444;
w446 <= not w356 and not w442;
w447 <= not w15 and w446;
w448 <= w445 and not w447;
w449 <= a(11) and not w448;
w450 <= a(11) and not w449;
w451 <= not w448 and not w449;
w452 <= not w450 and not w451;
w453 <= w434 and not w452;
w454 <= not w434 and w452;
w455 <= not w453 and not w454;
w456 <= w433 and not w455;
w457 <= not w433 and w455;
w458 <= not w456 and not w457;
w459 <= not w422 and w458;
w460 <= w422 and not w458;
w461 <= not w459 and not w460;
w462 <= not w420 and w461;
w463 <= w461 and not w462;
w464 <= not w420 and not w462;
w465 <= not w463 and not w464;
w466 <= not w375 and not w381;
w467 <= w465 and w466;
w468 <= not w465 and not w466;
w469 <= not w467 and not w468;
w470 <= b(10) and w9;
w471 <= b(8) and w27;
w472 <= b(9) and w4;
w473 <= not w471 and not w472;
w474 <= not w470 and w473;
w475 <= not w390 and not w392;
w476 <= not b(9) and not b(10);
w477 <= b(9) and b(10);
w478 <= not w476 and not w477;
w479 <= not w475 and w478;
w480 <= w475 and not w478;
w481 <= not w479 and not w480;
w482 <= w12 and w481;
w483 <= w474 and not w482;
w484 <= a(2) and not w483;
w485 <= a(2) and not w484;
w486 <= not w483 and not w484;
w487 <= not w485 and not w486;
w488 <= not w469 and w487;
w489 <= w469 and not w487;
w490 <= not w488 and not w489;
w491 <= not w409 and w490;
w492 <= w409 and not w490;
w493 <= not w491 and not w492;
w494 <= not w489 and not w491;
w495 <= not w462 and not w468;
w496 <= b(8) and w105;
w497 <= b(6) and w146;
w498 <= b(7) and w100;
w499 <= not w497 and not w498;
w500 <= not w496 and w499;
w501 <= w108 and w328;
w502 <= w500 and not w501;
w503 <= a(5) and not w502;
w504 <= a(5) and not w503;
w505 <= not w502 and not w503;
w506 <= not w504 and not w505;
w507 <= not w457 and not w459;
w508 <= b(2) and w443;
w509 <= w356 and not w442;
w510 <= w437 and w509;
w511 <= b(0) and w510;
w512 <= b(1) and w438;
w513 <= not w511 and not w512;
w514 <= not w508 and w513;
w515 <= w39 and w446;
w516 <= w514 and not w515;
w517 <= a(11) and not w516;
w518 <= a(11) and not w517;
w519 <= not w516 and not w517;
w520 <= not w518 and not w519;
w521 <= not w453 and w520;
w522 <= w453 and not w520;
w523 <= not w521 and not w522;
w524 <= b(5) and w254;
w525 <= b(3) and w284;
w526 <= b(4) and w249;
w527 <= not w525 and not w526;
w528 <= not w524 and w527;
w529 <= w137 and w257;
w530 <= w528 and not w529;
w531 <= a(8) and not w530;
w532 <= a(8) and not w531;
w533 <= not w530 and not w531;
w534 <= not w532 and not w533;
w535 <= w523 and not w534;
w536 <= w523 and not w535;
w537 <= not w534 and not w535;
w538 <= not w536 and not w537;
w539 <= not w507 and not w538;
w540 <= w507 and w538;
w541 <= not w539 and not w540;
w542 <= not w506 and w541;
w543 <= not w506 and not w542;
w544 <= w541 and not w542;
w545 <= not w543 and not w544;
w546 <= not w495 and not w545;
w547 <= not w495 and not w546;
w548 <= not w545 and not w546;
w549 <= not w547 and not w548;
w550 <= b(11) and w9;
w551 <= b(9) and w27;
w552 <= b(10) and w4;
w553 <= not w551 and not w552;
w554 <= not w550 and w553;
w555 <= not w477 and not w479;
w556 <= not b(10) and not b(11);
w557 <= b(10) and b(11);
w558 <= not w556 and not w557;
w559 <= not w555 and w558;
w560 <= w555 and not w558;
w561 <= not w559 and not w560;
w562 <= w12 and w561;
w563 <= w554 and not w562;
w564 <= a(2) and not w563;
w565 <= a(2) and not w564;
w566 <= not w563 and not w564;
w567 <= not w565 and not w566;
w568 <= not w549 and w567;
w569 <= w549 and not w567;
w570 <= not w568 and not w569;
w571 <= not w494 and not w570;
w572 <= w494 and w570;
w573 <= not w571 and not w572;
w574 <= b(12) and w9;
w575 <= b(10) and w27;
w576 <= b(11) and w4;
w577 <= not w575 and not w576;
w578 <= not w574 and w577;
w579 <= not w557 and not w559;
w580 <= not b(11) and not b(12);
w581 <= b(11) and b(12);
w582 <= not w580 and not w581;
w583 <= not w579 and w582;
w584 <= w579 and not w582;
w585 <= not w583 and not w584;
w586 <= w12 and w585;
w587 <= w578 and not w586;
w588 <= a(2) and not w587;
w589 <= a(2) and not w588;
w590 <= not w587 and not w588;
w591 <= not w589 and not w590;
w592 <= b(6) and w254;
w593 <= b(4) and w284;
w594 <= b(5) and w249;
w595 <= not w593 and not w594;
w596 <= not w592 and w595;
w597 <= w202 and w257;
w598 <= w596 and not w597;
w599 <= a(8) and not w598;
w600 <= a(8) and not w599;
w601 <= not w598 and not w599;
w602 <= not w600 and not w601;
w603 <= a(11) and not a(12);
w604 <= not a(11) and a(12);
w605 <= not w603 and not w604;
w606 <= b(0) and not w605;
w607 <= not w522 and w606;
w608 <= w522 and not w606;
w609 <= not w607 and not w608;
w610 <= b(3) and w443;
w611 <= b(1) and w510;
w612 <= b(2) and w438;
w613 <= not w611 and not w612;
w614 <= not w610 and w613;
w615 <= w61 and w446;
w616 <= w614 and not w615;
w617 <= a(11) and not w616;
w618 <= a(11) and not w617;
w619 <= not w616 and not w617;
w620 <= not w618 and not w619;
w621 <= not w609 and not w620;
w622 <= w609 and w620;
w623 <= not w621 and not w622;
w624 <= not w602 and w623;
w625 <= w623 and not w624;
w626 <= not w602 and not w624;
w627 <= not w625 and not w626;
w628 <= not w535 and not w539;
w629 <= w627 and w628;
w630 <= not w627 and not w628;
w631 <= not w629 and not w630;
w632 <= b(9) and w105;
w633 <= b(7) and w146;
w634 <= b(8) and w100;
w635 <= not w633 and not w634;
w636 <= not w632 and w635;
w637 <= w108 and w394;
w638 <= w636 and not w637;
w639 <= a(5) and not w638;
w640 <= a(5) and not w639;
w641 <= not w638 and not w639;
w642 <= not w640 and not w641;
w643 <= not w631 and w642;
w644 <= w631 and not w642;
w645 <= not w643 and not w644;
w646 <= not w542 and not w546;
w647 <= w645 and not w646;
w648 <= not w645 and w646;
w649 <= not w647 and not w648;
w650 <= not w591 and w649;
w651 <= w649 and not w650;
w652 <= not w591 and not w650;
w653 <= not w651 and not w652;
w654 <= not w549 and not w567;
w655 <= not w571 and not w654;
w656 <= not w653 and not w655;
w657 <= w653 and w655;
w658 <= not w656 and not w657;
w659 <= not w650 and not w656;
w660 <= not w644 and not w647;
w661 <= b(7) and w254;
w662 <= b(5) and w284;
w663 <= b(6) and w249;
w664 <= not w662 and not w663;
w665 <= not w661 and w664;
w666 <= w227 and w257;
w667 <= w665 and not w666;
w668 <= a(8) and not w667;
w669 <= a(8) and not w668;
w670 <= not w667 and not w668;
w671 <= not w669 and not w670;
w672 <= w522 and w606;
w673 <= not w621 and not w672;
w674 <= b(4) and w443;
w675 <= b(2) and w510;
w676 <= b(3) and w438;
w677 <= not w675 and not w676;
w678 <= not w674 and w677;
w679 <= w89 and w446;
w680 <= w678 and not w679;
w681 <= a(11) and not w680;
w682 <= a(11) and not w681;
w683 <= not w680 and not w681;
w684 <= not w682 and not w683;
w685 <= a(14) and not w606;
w686 <= not a(12) and a(13);
w687 <= a(12) and not a(13);
w688 <= not w686 and not w687;
w689 <= w605 and not w688;
w690 <= b(0) and w689;
w691 <= not a(13) and a(14);
w692 <= a(13) and not a(14);
w693 <= not w691 and not w692;
w694 <= not w605 and w693;
w695 <= b(1) and w694;
w696 <= not w690 and not w695;
w697 <= not w605 and not w693;
w698 <= not w15 and w697;
w699 <= w696 and not w698;
w700 <= a(14) and not w699;
w701 <= a(14) and not w700;
w702 <= not w699 and not w700;
w703 <= not w701 and not w702;
w704 <= w685 and not w703;
w705 <= not w685 and w703;
w706 <= not w704 and not w705;
w707 <= w684 and not w706;
w708 <= not w684 and w706;
w709 <= not w707 and not w708;
w710 <= not w673 and w709;
w711 <= w673 and not w709;
w712 <= not w710 and not w711;
w713 <= not w671 and w712;
w714 <= w712 and not w713;
w715 <= not w671 and not w713;
w716 <= not w714 and not w715;
w717 <= not w624 and not w630;
w718 <= w716 and w717;
w719 <= not w716 and not w717;
w720 <= not w718 and not w719;
w721 <= b(10) and w105;
w722 <= b(8) and w146;
w723 <= b(9) and w100;
w724 <= not w722 and not w723;
w725 <= not w721 and w724;
w726 <= w108 and w481;
w727 <= w725 and not w726;
w728 <= a(5) and not w727;
w729 <= a(5) and not w728;
w730 <= not w727 and not w728;
w731 <= not w729 and not w730;
w732 <= w720 and not w731;
w733 <= not w720 and w731;
w734 <= not w660 and not w733;
w735 <= not w732 and w734;
w736 <= not w660 and not w735;
w737 <= not w732 and not w735;
w738 <= not w733 and w737;
w739 <= not w736 and not w738;
w740 <= b(13) and w9;
w741 <= b(11) and w27;
w742 <= b(12) and w4;
w743 <= not w741 and not w742;
w744 <= not w740 and w743;
w745 <= not w581 and not w583;
w746 <= not b(12) and not b(13);
w747 <= b(12) and b(13);
w748 <= not w746 and not w747;
w749 <= not w745 and w748;
w750 <= w745 and not w748;
w751 <= not w749 and not w750;
w752 <= w12 and w751;
w753 <= w744 and not w752;
w754 <= a(2) and not w753;
w755 <= a(2) and not w754;
w756 <= not w753 and not w754;
w757 <= not w755 and not w756;
w758 <= not w739 and w757;
w759 <= w739 and not w757;
w760 <= not w758 and not w759;
w761 <= not w659 and not w760;
w762 <= w659 and w760;
w763 <= not w761 and not w762;
w764 <= not w739 and not w757;
w765 <= not w761 and not w764;
w766 <= b(14) and w9;
w767 <= b(12) and w27;
w768 <= b(13) and w4;
w769 <= not w767 and not w768;
w770 <= not w766 and w769;
w771 <= not w747 and not w749;
w772 <= not b(13) and not b(14);
w773 <= b(13) and b(14);
w774 <= not w772 and not w773;
w775 <= not w771 and w774;
w776 <= w771 and not w774;
w777 <= not w775 and not w776;
w778 <= w12 and w777;
w779 <= w770 and not w778;
w780 <= a(2) and not w779;
w781 <= a(2) and not w780;
w782 <= not w779 and not w780;
w783 <= not w781 and not w782;
w784 <= b(11) and w105;
w785 <= b(9) and w146;
w786 <= b(10) and w100;
w787 <= not w785 and not w786;
w788 <= not w784 and w787;
w789 <= w108 and w561;
w790 <= w788 and not w789;
w791 <= a(5) and not w790;
w792 <= a(5) and not w791;
w793 <= not w790 and not w791;
w794 <= not w792 and not w793;
w795 <= not w713 and not w719;
w796 <= not w708 and not w710;
w797 <= b(2) and w694;
w798 <= w605 and not w693;
w799 <= w688 and w798;
w800 <= b(0) and w799;
w801 <= b(1) and w689;
w802 <= not w800 and not w801;
w803 <= not w797 and w802;
w804 <= w39 and w697;
w805 <= w803 and not w804;
w806 <= a(14) and not w805;
w807 <= a(14) and not w806;
w808 <= not w805 and not w806;
w809 <= not w807 and not w808;
w810 <= not w704 and w809;
w811 <= w704 and not w809;
w812 <= not w810 and not w811;
w813 <= b(5) and w443;
w814 <= b(3) and w510;
w815 <= b(4) and w438;
w816 <= not w814 and not w815;
w817 <= not w813 and w816;
w818 <= w137 and w446;
w819 <= w817 and not w818;
w820 <= a(11) and not w819;
w821 <= a(11) and not w820;
w822 <= not w819 and not w820;
w823 <= not w821 and not w822;
w824 <= w812 and not w823;
w825 <= not w812 and w823;
w826 <= not w796 and not w825;
w827 <= not w824 and w826;
w828 <= not w796 and not w827;
w829 <= not w824 and not w827;
w830 <= not w825 and w829;
w831 <= not w828 and not w830;
w832 <= b(8) and w254;
w833 <= b(6) and w284;
w834 <= b(7) and w249;
w835 <= not w833 and not w834;
w836 <= not w832 and w835;
w837 <= w257 and w328;
w838 <= w836 and not w837;
w839 <= a(8) and not w838;
w840 <= a(8) and not w839;
w841 <= not w838 and not w839;
w842 <= not w840 and not w841;
w843 <= w831 and w842;
w844 <= not w831 and not w842;
w845 <= not w843 and not w844;
w846 <= not w795 and w845;
w847 <= w795 and not w845;
w848 <= not w846 and not w847;
w849 <= w794 and not w848;
w850 <= not w794 and w848;
w851 <= not w849 and not w850;
w852 <= not w737 and w851;
w853 <= w737 and not w851;
w854 <= not w852 and not w853;
w855 <= w783 and w854;
w856 <= not w783 and not w854;
w857 <= not w855 and not w856;
w858 <= not w765 and not w857;
w859 <= w765 and w857;
w860 <= not w858 and not w859;
w861 <= not w783 and w854;
w862 <= not w858 and not w861;
w863 <= b(15) and w9;
w864 <= b(13) and w27;
w865 <= b(14) and w4;
w866 <= not w864 and not w865;
w867 <= not w863 and w866;
w868 <= not w773 and not w775;
w869 <= not b(14) and not b(15);
w870 <= b(14) and b(15);
w871 <= not w869 and not w870;
w872 <= not w868 and w871;
w873 <= w868 and not w871;
w874 <= not w872 and not w873;
w875 <= w12 and w874;
w876 <= w867 and not w875;
w877 <= a(2) and not w876;
w878 <= a(2) and not w877;
w879 <= not w876 and not w877;
w880 <= not w878 and not w879;
w881 <= not w850 and not w852;
w882 <= b(12) and w105;
w883 <= b(10) and w146;
w884 <= b(11) and w100;
w885 <= not w883 and not w884;
w886 <= not w882 and w885;
w887 <= w108 and w585;
w888 <= w886 and not w887;
w889 <= a(5) and not w888;
w890 <= a(5) and not w889;
w891 <= not w888 and not w889;
w892 <= not w890 and not w891;
w893 <= not w844 and not w846;
w894 <= b(9) and w254;
w895 <= b(7) and w284;
w896 <= b(8) and w249;
w897 <= not w895 and not w896;
w898 <= not w894 and w897;
w899 <= w257 and w394;
w900 <= w898 and not w899;
w901 <= a(8) and not w900;
w902 <= a(8) and not w901;
w903 <= not w900 and not w901;
w904 <= not w902 and not w903;
w905 <= b(6) and w443;
w906 <= b(4) and w510;
w907 <= b(5) and w438;
w908 <= not w906 and not w907;
w909 <= not w905 and w908;
w910 <= w202 and w446;
w911 <= w909 and not w910;
w912 <= a(11) and not w911;
w913 <= a(11) and not w912;
w914 <= not w911 and not w912;
w915 <= not w913 and not w914;
w916 <= a(14) and not a(15);
w917 <= not a(14) and a(15);
w918 <= not w916 and not w917;
w919 <= b(0) and not w918;
w920 <= not w811 and w919;
w921 <= w811 and not w919;
w922 <= not w920 and not w921;
w923 <= b(3) and w694;
w924 <= b(1) and w799;
w925 <= b(2) and w689;
w926 <= not w924 and not w925;
w927 <= not w923 and w926;
w928 <= w61 and w697;
w929 <= w927 and not w928;
w930 <= a(14) and not w929;
w931 <= a(14) and not w930;
w932 <= not w929 and not w930;
w933 <= not w931 and not w932;
w934 <= not w922 and not w933;
w935 <= w922 and w933;
w936 <= not w934 and not w935;
w937 <= not w915 and w936;
w938 <= w936 and not w937;
w939 <= not w915 and not w937;
w940 <= not w938 and not w939;
w941 <= not w829 and not w940;
w942 <= w829 and w940;
w943 <= not w941 and not w942;
w944 <= not w904 and w943;
w945 <= not w904 and not w944;
w946 <= w943 and not w944;
w947 <= not w945 and not w946;
w948 <= not w893 and not w947;
w949 <= w893 and not w946;
w950 <= not w945 and w949;
w951 <= not w948 and not w950;
w952 <= not w892 and w951;
w953 <= not w892 and not w952;
w954 <= w951 and not w952;
w955 <= not w953 and not w954;
w956 <= not w881 and not w955;
w957 <= w881 and not w954;
w958 <= not w953 and w957;
w959 <= not w956 and not w958;
w960 <= not w880 and w959;
w961 <= not w880 and not w960;
w962 <= w959 and not w960;
w963 <= not w961 and not w962;
w964 <= not w862 and not w963;
w965 <= w862 and not w962;
w966 <= not w961 and w965;
w967 <= not w964 and not w966;
w968 <= not w960 and not w964;
w969 <= b(16) and w9;
w970 <= b(14) and w27;
w971 <= b(15) and w4;
w972 <= not w970 and not w971;
w973 <= not w969 and w972;
w974 <= not w870 and not w872;
w975 <= not b(15) and not b(16);
w976 <= b(15) and b(16);
w977 <= not w975 and not w976;
w978 <= not w974 and w977;
w979 <= w974 and not w977;
w980 <= not w978 and not w979;
w981 <= w12 and w980;
w982 <= w973 and not w981;
w983 <= a(2) and not w982;
w984 <= a(2) and not w983;
w985 <= not w982 and not w983;
w986 <= not w984 and not w985;
w987 <= not w952 and not w956;
w988 <= b(13) and w105;
w989 <= b(11) and w146;
w990 <= b(12) and w100;
w991 <= not w989 and not w990;
w992 <= not w988 and w991;
w993 <= w108 and w751;
w994 <= w992 and not w993;
w995 <= a(5) and not w994;
w996 <= a(5) and not w995;
w997 <= not w994 and not w995;
w998 <= not w996 and not w997;
w999 <= not w944 and not w948;
w1000 <= b(10) and w254;
w1001 <= b(8) and w284;
w1002 <= b(9) and w249;
w1003 <= not w1001 and not w1002;
w1004 <= not w1000 and w1003;
w1005 <= w257 and w481;
w1006 <= w1004 and not w1005;
w1007 <= a(8) and not w1006;
w1008 <= a(8) and not w1007;
w1009 <= not w1006 and not w1007;
w1010 <= not w1008 and not w1009;
w1011 <= not w937 and not w941;
w1012 <= b(7) and w443;
w1013 <= b(5) and w510;
w1014 <= b(6) and w438;
w1015 <= not w1013 and not w1014;
w1016 <= not w1012 and w1015;
w1017 <= w227 and w446;
w1018 <= w1016 and not w1017;
w1019 <= a(11) and not w1018;
w1020 <= a(11) and not w1019;
w1021 <= not w1018 and not w1019;
w1022 <= not w1020 and not w1021;
w1023 <= w811 and w919;
w1024 <= not w934 and not w1023;
w1025 <= b(4) and w694;
w1026 <= b(2) and w799;
w1027 <= b(3) and w689;
w1028 <= not w1026 and not w1027;
w1029 <= not w1025 and w1028;
w1030 <= w89 and w697;
w1031 <= w1029 and not w1030;
w1032 <= a(14) and not w1031;
w1033 <= a(14) and not w1032;
w1034 <= not w1031 and not w1032;
w1035 <= not w1033 and not w1034;
w1036 <= a(17) and not w919;
w1037 <= not a(15) and a(16);
w1038 <= a(15) and not a(16);
w1039 <= not w1037 and not w1038;
w1040 <= w918 and not w1039;
w1041 <= b(0) and w1040;
w1042 <= not a(16) and a(17);
w1043 <= a(16) and not a(17);
w1044 <= not w1042 and not w1043;
w1045 <= not w918 and w1044;
w1046 <= b(1) and w1045;
w1047 <= not w1041 and not w1046;
w1048 <= not w918 and not w1044;
w1049 <= not w15 and w1048;
w1050 <= w1047 and not w1049;
w1051 <= a(17) and not w1050;
w1052 <= a(17) and not w1051;
w1053 <= not w1050 and not w1051;
w1054 <= not w1052 and not w1053;
w1055 <= w1036 and not w1054;
w1056 <= not w1036 and w1054;
w1057 <= not w1055 and not w1056;
w1058 <= w1035 and not w1057;
w1059 <= not w1035 and w1057;
w1060 <= not w1058 and not w1059;
w1061 <= not w1024 and w1060;
w1062 <= w1024 and not w1060;
w1063 <= not w1061 and not w1062;
w1064 <= w1022 and not w1063;
w1065 <= not w1022 and w1063;
w1066 <= not w1064 and not w1065;
w1067 <= not w1011 and w1066;
w1068 <= w1011 and not w1066;
w1069 <= not w1067 and not w1068;
w1070 <= w1010 and not w1069;
w1071 <= not w1010 and w1069;
w1072 <= not w1070 and not w1071;
w1073 <= not w999 and w1072;
w1074 <= w999 and not w1072;
w1075 <= not w1073 and not w1074;
w1076 <= w998 and not w1075;
w1077 <= not w998 and w1075;
w1078 <= not w1076 and not w1077;
w1079 <= not w987 and w1078;
w1080 <= w987 and not w1078;
w1081 <= not w1079 and not w1080;
w1082 <= w986 and w1081;
w1083 <= not w986 and not w1081;
w1084 <= not w1082 and not w1083;
w1085 <= not w968 and not w1084;
w1086 <= w968 and w1084;
w1087 <= not w1085 and not w1086;
w1088 <= b(17) and w9;
w1089 <= b(15) and w27;
w1090 <= b(16) and w4;
w1091 <= not w1089 and not w1090;
w1092 <= not w1088 and w1091;
w1093 <= not w976 and not w978;
w1094 <= not b(16) and not b(17);
w1095 <= b(16) and b(17);
w1096 <= not w1094 and not w1095;
w1097 <= not w1093 and w1096;
w1098 <= w1093 and not w1096;
w1099 <= not w1097 and not w1098;
w1100 <= w12 and w1099;
w1101 <= w1092 and not w1100;
w1102 <= a(2) and not w1101;
w1103 <= a(2) and not w1102;
w1104 <= not w1101 and not w1102;
w1105 <= not w1103 and not w1104;
w1106 <= not w1077 and not w1079;
w1107 <= b(14) and w105;
w1108 <= b(12) and w146;
w1109 <= b(13) and w100;
w1110 <= not w1108 and not w1109;
w1111 <= not w1107 and w1110;
w1112 <= w108 and w777;
w1113 <= w1111 and not w1112;
w1114 <= a(5) and not w1113;
w1115 <= a(5) and not w1114;
w1116 <= not w1113 and not w1114;
w1117 <= not w1115 and not w1116;
w1118 <= not w1071 and not w1073;
w1119 <= b(11) and w254;
w1120 <= b(9) and w284;
w1121 <= b(10) and w249;
w1122 <= not w1120 and not w1121;
w1123 <= not w1119 and w1122;
w1124 <= w257 and w561;
w1125 <= w1123 and not w1124;
w1126 <= a(8) and not w1125;
w1127 <= a(8) and not w1126;
w1128 <= not w1125 and not w1126;
w1129 <= not w1127 and not w1128;
w1130 <= not w1065 and not w1067;
w1131 <= not w1059 and not w1061;
w1132 <= b(2) and w1045;
w1133 <= w918 and not w1044;
w1134 <= w1039 and w1133;
w1135 <= b(0) and w1134;
w1136 <= b(1) and w1040;
w1137 <= not w1135 and not w1136;
w1138 <= not w1132 and w1137;
w1139 <= w39 and w1048;
w1140 <= w1138 and not w1139;
w1141 <= a(17) and not w1140;
w1142 <= a(17) and not w1141;
w1143 <= not w1140 and not w1141;
w1144 <= not w1142 and not w1143;
w1145 <= not w1055 and w1144;
w1146 <= w1055 and not w1144;
w1147 <= not w1145 and not w1146;
w1148 <= b(5) and w694;
w1149 <= b(3) and w799;
w1150 <= b(4) and w689;
w1151 <= not w1149 and not w1150;
w1152 <= not w1148 and w1151;
w1153 <= w137 and w697;
w1154 <= w1152 and not w1153;
w1155 <= a(14) and not w1154;
w1156 <= a(14) and not w1155;
w1157 <= not w1154 and not w1155;
w1158 <= not w1156 and not w1157;
w1159 <= w1147 and not w1158;
w1160 <= not w1147 and w1158;
w1161 <= not w1131 and not w1160;
w1162 <= not w1159 and w1161;
w1163 <= not w1131 and not w1162;
w1164 <= not w1159 and not w1162;
w1165 <= not w1160 and w1164;
w1166 <= not w1163 and not w1165;
w1167 <= b(8) and w443;
w1168 <= b(6) and w510;
w1169 <= b(7) and w438;
w1170 <= not w1168 and not w1169;
w1171 <= not w1167 and w1170;
w1172 <= w328 and w446;
w1173 <= w1171 and not w1172;
w1174 <= a(11) and not w1173;
w1175 <= a(11) and not w1174;
w1176 <= not w1173 and not w1174;
w1177 <= not w1175 and not w1176;
w1178 <= w1166 and w1177;
w1179 <= not w1166 and not w1177;
w1180 <= not w1178 and not w1179;
w1181 <= not w1130 and w1180;
w1182 <= w1130 and not w1180;
w1183 <= not w1181 and not w1182;
w1184 <= w1129 and not w1183;
w1185 <= not w1129 and w1183;
w1186 <= not w1184 and not w1185;
w1187 <= not w1118 and w1186;
w1188 <= w1118 and not w1186;
w1189 <= not w1187 and not w1188;
w1190 <= w1117 and not w1189;
w1191 <= not w1117 and w1189;
w1192 <= not w1190 and not w1191;
w1193 <= not w1106 and w1192;
w1194 <= w1106 and not w1192;
w1195 <= not w1193 and not w1194;
w1196 <= not w1105 and w1195;
w1197 <= w1195 and not w1196;
w1198 <= not w1105 and not w1196;
w1199 <= not w1197 and not w1198;
w1200 <= not w986 and w1081;
w1201 <= not w1085 and not w1200;
w1202 <= not w1199 and not w1201;
w1203 <= w1199 and w1201;
w1204 <= not w1202 and not w1203;
w1205 <= not w1191 and not w1193;
w1206 <= b(15) and w105;
w1207 <= b(13) and w146;
w1208 <= b(14) and w100;
w1209 <= not w1207 and not w1208;
w1210 <= not w1206 and w1209;
w1211 <= w108 and w874;
w1212 <= w1210 and not w1211;
w1213 <= a(5) and not w1212;
w1214 <= a(5) and not w1213;
w1215 <= not w1212 and not w1213;
w1216 <= not w1214 and not w1215;
w1217 <= not w1185 and not w1187;
w1218 <= b(12) and w254;
w1219 <= b(10) and w284;
w1220 <= b(11) and w249;
w1221 <= not w1219 and not w1220;
w1222 <= not w1218 and w1221;
w1223 <= w257 and w585;
w1224 <= w1222 and not w1223;
w1225 <= a(8) and not w1224;
w1226 <= a(8) and not w1225;
w1227 <= not w1224 and not w1225;
w1228 <= not w1226 and not w1227;
w1229 <= not w1179 and not w1181;
w1230 <= b(6) and w694;
w1231 <= b(4) and w799;
w1232 <= b(5) and w689;
w1233 <= not w1231 and not w1232;
w1234 <= not w1230 and w1233;
w1235 <= w202 and w697;
w1236 <= w1234 and not w1235;
w1237 <= a(14) and not w1236;
w1238 <= a(14) and not w1237;
w1239 <= not w1236 and not w1237;
w1240 <= not w1238 and not w1239;
w1241 <= a(17) and not a(18);
w1242 <= not a(17) and a(18);
w1243 <= not w1241 and not w1242;
w1244 <= b(0) and not w1243;
w1245 <= not w1146 and w1244;
w1246 <= w1146 and not w1244;
w1247 <= not w1245 and not w1246;
w1248 <= b(3) and w1045;
w1249 <= b(1) and w1134;
w1250 <= b(2) and w1040;
w1251 <= not w1249 and not w1250;
w1252 <= not w1248 and w1251;
w1253 <= w61 and w1048;
w1254 <= w1252 and not w1253;
w1255 <= a(17) and not w1254;
w1256 <= a(17) and not w1255;
w1257 <= not w1254 and not w1255;
w1258 <= not w1256 and not w1257;
w1259 <= not w1247 and not w1258;
w1260 <= w1247 and w1258;
w1261 <= not w1259 and not w1260;
w1262 <= not w1240 and w1261;
w1263 <= w1261 and not w1262;
w1264 <= not w1240 and not w1262;
w1265 <= not w1263 and not w1264;
w1266 <= not w1164 and w1265;
w1267 <= w1164 and not w1265;
w1268 <= not w1266 and not w1267;
w1269 <= b(9) and w443;
w1270 <= b(7) and w510;
w1271 <= b(8) and w438;
w1272 <= not w1270 and not w1271;
w1273 <= not w1269 and w1272;
w1274 <= w394 and w446;
w1275 <= w1273 and not w1274;
w1276 <= a(11) and not w1275;
w1277 <= a(11) and not w1276;
w1278 <= not w1275 and not w1276;
w1279 <= not w1277 and not w1278;
w1280 <= not w1268 and not w1279;
w1281 <= w1268 and w1279;
w1282 <= not w1280 and not w1281;
w1283 <= not w1229 and w1282;
w1284 <= w1229 and not w1282;
w1285 <= not w1283 and not w1284;
w1286 <= w1228 and not w1285;
w1287 <= not w1228 and w1285;
w1288 <= not w1286 and not w1287;
w1289 <= not w1217 and w1288;
w1290 <= w1217 and not w1288;
w1291 <= not w1289 and not w1290;
w1292 <= not w1216 and w1291;
w1293 <= w1216 and not w1291;
w1294 <= not w1292 and not w1293;
w1295 <= not w1205 and w1294;
w1296 <= w1205 and not w1294;
w1297 <= not w1295 and not w1296;
w1298 <= b(18) and w9;
w1299 <= b(16) and w27;
w1300 <= b(17) and w4;
w1301 <= not w1299 and not w1300;
w1302 <= not w1298 and w1301;
w1303 <= not w1095 and not w1097;
w1304 <= not b(17) and not b(18);
w1305 <= b(17) and b(18);
w1306 <= not w1304 and not w1305;
w1307 <= not w1303 and w1306;
w1308 <= w1303 and not w1306;
w1309 <= not w1307 and not w1308;
w1310 <= w12 and w1309;
w1311 <= w1302 and not w1310;
w1312 <= a(2) and not w1311;
w1313 <= a(2) and not w1312;
w1314 <= not w1311 and not w1312;
w1315 <= not w1313 and not w1314;
w1316 <= w1297 and not w1315;
w1317 <= w1297 and not w1316;
w1318 <= not w1315 and not w1316;
w1319 <= not w1317 and not w1318;
w1320 <= not w1196 and not w1202;
w1321 <= not w1319 and not w1320;
w1322 <= w1319 and w1320;
w1323 <= not w1321 and not w1322;
w1324 <= b(16) and w105;
w1325 <= b(14) and w146;
w1326 <= b(15) and w100;
w1327 <= not w1325 and not w1326;
w1328 <= not w1324 and w1327;
w1329 <= w108 and w980;
w1330 <= w1328 and not w1329;
w1331 <= a(5) and not w1330;
w1332 <= a(5) and not w1331;
w1333 <= not w1330 and not w1331;
w1334 <= not w1332 and not w1333;
w1335 <= not w1164 and not w1265;
w1336 <= not w1262 and not w1335;
w1337 <= b(7) and w694;
w1338 <= b(5) and w799;
w1339 <= b(6) and w689;
w1340 <= not w1338 and not w1339;
w1341 <= not w1337 and w1340;
w1342 <= w227 and w697;
w1343 <= w1341 and not w1342;
w1344 <= a(14) and not w1343;
w1345 <= a(14) and not w1344;
w1346 <= not w1343 and not w1344;
w1347 <= not w1345 and not w1346;
w1348 <= w1146 and w1244;
w1349 <= not w1259 and not w1348;
w1350 <= b(4) and w1045;
w1351 <= b(2) and w1134;
w1352 <= b(3) and w1040;
w1353 <= not w1351 and not w1352;
w1354 <= not w1350 and w1353;
w1355 <= w89 and w1048;
w1356 <= w1354 and not w1355;
w1357 <= a(17) and not w1356;
w1358 <= a(17) and not w1357;
w1359 <= not w1356 and not w1357;
w1360 <= not w1358 and not w1359;
w1361 <= a(20) and not w1244;
w1362 <= not a(18) and a(19);
w1363 <= a(18) and not a(19);
w1364 <= not w1362 and not w1363;
w1365 <= w1243 and not w1364;
w1366 <= b(0) and w1365;
w1367 <= not a(19) and a(20);
w1368 <= a(19) and not a(20);
w1369 <= not w1367 and not w1368;
w1370 <= not w1243 and w1369;
w1371 <= b(1) and w1370;
w1372 <= not w1366 and not w1371;
w1373 <= not w1243 and not w1369;
w1374 <= not w15 and w1373;
w1375 <= w1372 and not w1374;
w1376 <= a(20) and not w1375;
w1377 <= a(20) and not w1376;
w1378 <= not w1375 and not w1376;
w1379 <= not w1377 and not w1378;
w1380 <= w1361 and not w1379;
w1381 <= not w1361 and w1379;
w1382 <= not w1380 and not w1381;
w1383 <= w1360 and w1382;
w1384 <= not w1360 and not w1382;
w1385 <= not w1383 and not w1384;
w1386 <= not w1349 and not w1385;
w1387 <= w1349 and w1385;
w1388 <= not w1386 and not w1387;
w1389 <= not w1347 and w1388;
w1390 <= w1347 and not w1388;
w1391 <= not w1389 and not w1390;
w1392 <= not w1336 and w1391;
w1393 <= w1336 and not w1391;
w1394 <= not w1392 and not w1393;
w1395 <= b(10) and w443;
w1396 <= b(8) and w510;
w1397 <= b(9) and w438;
w1398 <= not w1396 and not w1397;
w1399 <= not w1395 and w1398;
w1400 <= w446 and w481;
w1401 <= w1399 and not w1400;
w1402 <= a(11) and not w1401;
w1403 <= a(11) and not w1402;
w1404 <= not w1401 and not w1402;
w1405 <= not w1403 and not w1404;
w1406 <= w1394 and not w1405;
w1407 <= w1394 and not w1406;
w1408 <= not w1405 and not w1406;
w1409 <= not w1407 and not w1408;
w1410 <= not w1280 and not w1283;
w1411 <= w1409 and w1410;
w1412 <= not w1409 and not w1410;
w1413 <= not w1411 and not w1412;
w1414 <= b(13) and w254;
w1415 <= b(11) and w284;
w1416 <= b(12) and w249;
w1417 <= not w1415 and not w1416;
w1418 <= not w1414 and w1417;
w1419 <= w257 and w751;
w1420 <= w1418 and not w1419;
w1421 <= a(8) and not w1420;
w1422 <= a(8) and not w1421;
w1423 <= not w1420 and not w1421;
w1424 <= not w1422 and not w1423;
w1425 <= not w1413 and w1424;
w1426 <= w1413 and not w1424;
w1427 <= not w1425 and not w1426;
w1428 <= not w1287 and not w1289;
w1429 <= w1427 and not w1428;
w1430 <= not w1427 and w1428;
w1431 <= not w1429 and not w1430;
w1432 <= not w1334 and w1431;
w1433 <= w1431 and not w1432;
w1434 <= not w1334 and not w1432;
w1435 <= not w1433 and not w1434;
w1436 <= not w1292 and not w1295;
w1437 <= w1435 and w1436;
w1438 <= not w1435 and not w1436;
w1439 <= not w1437 and not w1438;
w1440 <= b(19) and w9;
w1441 <= b(17) and w27;
w1442 <= b(18) and w4;
w1443 <= not w1441 and not w1442;
w1444 <= not w1440 and w1443;
w1445 <= not w1305 and not w1307;
w1446 <= not b(18) and not b(19);
w1447 <= b(18) and b(19);
w1448 <= not w1446 and not w1447;
w1449 <= not w1445 and w1448;
w1450 <= w1445 and not w1448;
w1451 <= not w1449 and not w1450;
w1452 <= w12 and w1451;
w1453 <= w1444 and not w1452;
w1454 <= a(2) and not w1453;
w1455 <= a(2) and not w1454;
w1456 <= not w1453 and not w1454;
w1457 <= not w1455 and not w1456;
w1458 <= w1439 and not w1457;
w1459 <= w1439 and not w1458;
w1460 <= not w1457 and not w1458;
w1461 <= not w1459 and not w1460;
w1462 <= not w1316 and not w1321;
w1463 <= not w1461 and not w1462;
w1464 <= w1461 and w1462;
w1465 <= not w1463 and not w1464;
w1466 <= not w1432 and not w1438;
w1467 <= b(17) and w105;
w1468 <= b(15) and w146;
w1469 <= b(16) and w100;
w1470 <= not w1468 and not w1469;
w1471 <= not w1467 and w1470;
w1472 <= w108 and w1099;
w1473 <= w1471 and not w1472;
w1474 <= a(5) and not w1473;
w1475 <= a(5) and not w1474;
w1476 <= not w1473 and not w1474;
w1477 <= not w1475 and not w1476;
w1478 <= b(14) and w254;
w1479 <= b(12) and w284;
w1480 <= b(13) and w249;
w1481 <= not w1479 and not w1480;
w1482 <= not w1478 and w1481;
w1483 <= w257 and w777;
w1484 <= w1482 and not w1483;
w1485 <= a(8) and not w1484;
w1486 <= a(8) and not w1485;
w1487 <= not w1484 and not w1485;
w1488 <= not w1486 and not w1487;
w1489 <= not w1406 and not w1412;
w1490 <= b(11) and w443;
w1491 <= b(9) and w510;
w1492 <= b(10) and w438;
w1493 <= not w1491 and not w1492;
w1494 <= not w1490 and w1493;
w1495 <= w446 and w561;
w1496 <= w1494 and not w1495;
w1497 <= a(11) and not w1496;
w1498 <= a(11) and not w1497;
w1499 <= not w1496 and not w1497;
w1500 <= not w1498 and not w1499;
w1501 <= not w1389 and not w1392;
w1502 <= not w1360 and w1382;
w1503 <= not w1386 and not w1502;
w1504 <= b(2) and w1370;
w1505 <= w1243 and not w1369;
w1506 <= w1364 and w1505;
w1507 <= b(0) and w1506;
w1508 <= b(1) and w1365;
w1509 <= not w1507 and not w1508;
w1510 <= not w1504 and w1509;
w1511 <= w39 and w1373;
w1512 <= w1510 and not w1511;
w1513 <= a(20) and not w1512;
w1514 <= a(20) and not w1513;
w1515 <= not w1512 and not w1513;
w1516 <= not w1514 and not w1515;
w1517 <= not w1380 and w1516;
w1518 <= w1380 and not w1516;
w1519 <= not w1517 and not w1518;
w1520 <= b(5) and w1045;
w1521 <= b(3) and w1134;
w1522 <= b(4) and w1040;
w1523 <= not w1521 and not w1522;
w1524 <= not w1520 and w1523;
w1525 <= w137 and w1048;
w1526 <= w1524 and not w1525;
w1527 <= a(17) and not w1526;
w1528 <= a(17) and not w1527;
w1529 <= not w1526 and not w1527;
w1530 <= not w1528 and not w1529;
w1531 <= w1519 and not w1530;
w1532 <= not w1519 and w1530;
w1533 <= not w1503 and not w1532;
w1534 <= not w1531 and w1533;
w1535 <= not w1503 and not w1534;
w1536 <= not w1531 and not w1534;
w1537 <= not w1532 and w1536;
w1538 <= not w1535 and not w1537;
w1539 <= b(8) and w694;
w1540 <= b(6) and w799;
w1541 <= b(7) and w689;
w1542 <= not w1540 and not w1541;
w1543 <= not w1539 and w1542;
w1544 <= w328 and w697;
w1545 <= w1543 and not w1544;
w1546 <= a(14) and not w1545;
w1547 <= a(14) and not w1546;
w1548 <= not w1545 and not w1546;
w1549 <= not w1547 and not w1548;
w1550 <= w1538 and w1549;
w1551 <= not w1538 and not w1549;
w1552 <= not w1550 and not w1551;
w1553 <= not w1501 and w1552;
w1554 <= w1501 and not w1552;
w1555 <= not w1553 and not w1554;
w1556 <= w1500 and not w1555;
w1557 <= not w1500 and w1555;
w1558 <= not w1556 and not w1557;
w1559 <= not w1489 and w1558;
w1560 <= w1489 and not w1558;
w1561 <= not w1559 and not w1560;
w1562 <= not w1488 and w1561;
w1563 <= w1561 and not w1562;
w1564 <= not w1488 and not w1562;
w1565 <= not w1563 and not w1564;
w1566 <= not w1426 and not w1429;
w1567 <= not w1565 and not w1566;
w1568 <= w1565 and w1566;
w1569 <= not w1567 and not w1568;
w1570 <= not w1477 and w1569;
w1571 <= not w1477 and not w1570;
w1572 <= w1569 and not w1570;
w1573 <= not w1571 and not w1572;
w1574 <= not w1466 and not w1573;
w1575 <= not w1466 and not w1574;
w1576 <= not w1573 and not w1574;
w1577 <= not w1575 and not w1576;
w1578 <= b(20) and w9;
w1579 <= b(18) and w27;
w1580 <= b(19) and w4;
w1581 <= not w1579 and not w1580;
w1582 <= not w1578 and w1581;
w1583 <= not w1447 and not w1449;
w1584 <= not b(19) and not b(20);
w1585 <= b(19) and b(20);
w1586 <= not w1584 and not w1585;
w1587 <= not w1583 and w1586;
w1588 <= w1583 and not w1586;
w1589 <= not w1587 and not w1588;
w1590 <= w12 and w1589;
w1591 <= w1582 and not w1590;
w1592 <= a(2) and not w1591;
w1593 <= a(2) and not w1592;
w1594 <= not w1591 and not w1592;
w1595 <= not w1593 and not w1594;
w1596 <= not w1577 and not w1595;
w1597 <= not w1577 and not w1596;
w1598 <= not w1595 and not w1596;
w1599 <= not w1597 and not w1598;
w1600 <= not w1458 and not w1463;
w1601 <= not w1599 and not w1600;
w1602 <= w1599 and w1600;
w1603 <= not w1601 and not w1602;
w1604 <= not w1562 and not w1567;
w1605 <= b(15) and w254;
w1606 <= b(13) and w284;
w1607 <= b(14) and w249;
w1608 <= not w1606 and not w1607;
w1609 <= not w1605 and w1608;
w1610 <= w257 and w874;
w1611 <= w1609 and not w1610;
w1612 <= a(8) and not w1611;
w1613 <= a(8) and not w1612;
w1614 <= not w1611 and not w1612;
w1615 <= not w1613 and not w1614;
w1616 <= not w1557 and not w1559;
w1617 <= b(12) and w443;
w1618 <= b(10) and w510;
w1619 <= b(11) and w438;
w1620 <= not w1618 and not w1619;
w1621 <= not w1617 and w1620;
w1622 <= w446 and w585;
w1623 <= w1621 and not w1622;
w1624 <= a(11) and not w1623;
w1625 <= a(11) and not w1624;
w1626 <= not w1623 and not w1624;
w1627 <= not w1625 and not w1626;
w1628 <= not w1551 and not w1553;
w1629 <= b(6) and w1045;
w1630 <= b(4) and w1134;
w1631 <= b(5) and w1040;
w1632 <= not w1630 and not w1631;
w1633 <= not w1629 and w1632;
w1634 <= w202 and w1048;
w1635 <= w1633 and not w1634;
w1636 <= a(17) and not w1635;
w1637 <= a(17) and not w1636;
w1638 <= not w1635 and not w1636;
w1639 <= not w1637 and not w1638;
w1640 <= a(20) and not a(21);
w1641 <= not a(20) and a(21);
w1642 <= not w1640 and not w1641;
w1643 <= b(0) and not w1642;
w1644 <= not w1518 and w1643;
w1645 <= w1518 and not w1643;
w1646 <= not w1644 and not w1645;
w1647 <= b(3) and w1370;
w1648 <= b(1) and w1506;
w1649 <= b(2) and w1365;
w1650 <= not w1648 and not w1649;
w1651 <= not w1647 and w1650;
w1652 <= w61 and w1373;
w1653 <= w1651 and not w1652;
w1654 <= a(20) and not w1653;
w1655 <= a(20) and not w1654;
w1656 <= not w1653 and not w1654;
w1657 <= not w1655 and not w1656;
w1658 <= not w1646 and not w1657;
w1659 <= w1646 and w1657;
w1660 <= not w1658 and not w1659;
w1661 <= not w1639 and w1660;
w1662 <= w1660 and not w1661;
w1663 <= not w1639 and not w1661;
w1664 <= not w1662 and not w1663;
w1665 <= not w1536 and w1664;
w1666 <= w1536 and not w1664;
w1667 <= not w1665 and not w1666;
w1668 <= b(9) and w694;
w1669 <= b(7) and w799;
w1670 <= b(8) and w689;
w1671 <= not w1669 and not w1670;
w1672 <= not w1668 and w1671;
w1673 <= w394 and w697;
w1674 <= w1672 and not w1673;
w1675 <= a(14) and not w1674;
w1676 <= a(14) and not w1675;
w1677 <= not w1674 and not w1675;
w1678 <= not w1676 and not w1677;
w1679 <= not w1667 and not w1678;
w1680 <= w1667 and w1678;
w1681 <= not w1679 and not w1680;
w1682 <= not w1628 and w1681;
w1683 <= w1628 and not w1681;
w1684 <= not w1682 and not w1683;
w1685 <= w1627 and not w1684;
w1686 <= not w1627 and w1684;
w1687 <= not w1685 and not w1686;
w1688 <= not w1616 and w1687;
w1689 <= w1616 and not w1687;
w1690 <= not w1688 and not w1689;
w1691 <= not w1615 and w1690;
w1692 <= w1615 and not w1690;
w1693 <= not w1691 and not w1692;
w1694 <= not w1604 and w1693;
w1695 <= w1604 and not w1693;
w1696 <= not w1694 and not w1695;
w1697 <= b(18) and w105;
w1698 <= b(16) and w146;
w1699 <= b(17) and w100;
w1700 <= not w1698 and not w1699;
w1701 <= not w1697 and w1700;
w1702 <= w108 and w1309;
w1703 <= w1701 and not w1702;
w1704 <= a(5) and not w1703;
w1705 <= a(5) and not w1704;
w1706 <= not w1703 and not w1704;
w1707 <= not w1705 and not w1706;
w1708 <= w1696 and not w1707;
w1709 <= w1696 and not w1708;
w1710 <= not w1707 and not w1708;
w1711 <= not w1709 and not w1710;
w1712 <= not w1570 and not w1574;
w1713 <= w1711 and w1712;
w1714 <= not w1711 and not w1712;
w1715 <= not w1713 and not w1714;
w1716 <= b(21) and w9;
w1717 <= b(19) and w27;
w1718 <= b(20) and w4;
w1719 <= not w1717 and not w1718;
w1720 <= not w1716 and w1719;
w1721 <= not w1585 and not w1587;
w1722 <= not b(20) and not b(21);
w1723 <= b(20) and b(21);
w1724 <= not w1722 and not w1723;
w1725 <= not w1721 and w1724;
w1726 <= w1721 and not w1724;
w1727 <= not w1725 and not w1726;
w1728 <= w12 and w1727;
w1729 <= w1720 and not w1728;
w1730 <= a(2) and not w1729;
w1731 <= a(2) and not w1730;
w1732 <= not w1729 and not w1730;
w1733 <= not w1731 and not w1732;
w1734 <= w1715 and not w1733;
w1735 <= w1715 and not w1734;
w1736 <= not w1733 and not w1734;
w1737 <= not w1735 and not w1736;
w1738 <= not w1596 and not w1601;
w1739 <= not w1737 and not w1738;
w1740 <= w1737 and w1738;
w1741 <= not w1739 and not w1740;
w1742 <= not w1734 and not w1739;
w1743 <= not w1691 and not w1694;
w1744 <= b(16) and w254;
w1745 <= b(14) and w284;
w1746 <= b(15) and w249;
w1747 <= not w1745 and not w1746;
w1748 <= not w1744 and w1747;
w1749 <= w257 and w980;
w1750 <= w1748 and not w1749;
w1751 <= a(8) and not w1750;
w1752 <= a(8) and not w1751;
w1753 <= not w1750 and not w1751;
w1754 <= not w1752 and not w1753;
w1755 <= not w1686 and not w1688;
w1756 <= not w1536 and not w1664;
w1757 <= not w1661 and not w1756;
w1758 <= b(7) and w1045;
w1759 <= b(5) and w1134;
w1760 <= b(6) and w1040;
w1761 <= not w1759 and not w1760;
w1762 <= not w1758 and w1761;
w1763 <= w227 and w1048;
w1764 <= w1762 and not w1763;
w1765 <= a(17) and not w1764;
w1766 <= a(17) and not w1765;
w1767 <= not w1764 and not w1765;
w1768 <= not w1766 and not w1767;
w1769 <= w1518 and w1643;
w1770 <= not w1658 and not w1769;
w1771 <= b(4) and w1370;
w1772 <= b(2) and w1506;
w1773 <= b(3) and w1365;
w1774 <= not w1772 and not w1773;
w1775 <= not w1771 and w1774;
w1776 <= w89 and w1373;
w1777 <= w1775 and not w1776;
w1778 <= a(20) and not w1777;
w1779 <= a(20) and not w1778;
w1780 <= not w1777 and not w1778;
w1781 <= not w1779 and not w1780;
w1782 <= a(23) and not w1643;
w1783 <= not a(21) and a(22);
w1784 <= a(21) and not a(22);
w1785 <= not w1783 and not w1784;
w1786 <= w1642 and not w1785;
w1787 <= b(0) and w1786;
w1788 <= not a(22) and a(23);
w1789 <= a(22) and not a(23);
w1790 <= not w1788 and not w1789;
w1791 <= not w1642 and w1790;
w1792 <= b(1) and w1791;
w1793 <= not w1787 and not w1792;
w1794 <= not w1642 and not w1790;
w1795 <= not w15 and w1794;
w1796 <= w1793 and not w1795;
w1797 <= a(23) and not w1796;
w1798 <= a(23) and not w1797;
w1799 <= not w1796 and not w1797;
w1800 <= not w1798 and not w1799;
w1801 <= w1782 and not w1800;
w1802 <= not w1782 and w1800;
w1803 <= not w1801 and not w1802;
w1804 <= w1781 and w1803;
w1805 <= not w1781 and not w1803;
w1806 <= not w1804 and not w1805;
w1807 <= not w1770 and not w1806;
w1808 <= w1770 and w1806;
w1809 <= not w1807 and not w1808;
w1810 <= not w1768 and w1809;
w1811 <= w1768 and not w1809;
w1812 <= not w1810 and not w1811;
w1813 <= not w1757 and w1812;
w1814 <= w1757 and not w1812;
w1815 <= not w1813 and not w1814;
w1816 <= b(10) and w694;
w1817 <= b(8) and w799;
w1818 <= b(9) and w689;
w1819 <= not w1817 and not w1818;
w1820 <= not w1816 and w1819;
w1821 <= w481 and w697;
w1822 <= w1820 and not w1821;
w1823 <= a(14) and not w1822;
w1824 <= a(14) and not w1823;
w1825 <= not w1822 and not w1823;
w1826 <= not w1824 and not w1825;
w1827 <= w1815 and not w1826;
w1828 <= w1815 and not w1827;
w1829 <= not w1826 and not w1827;
w1830 <= not w1828 and not w1829;
w1831 <= not w1679 and not w1682;
w1832 <= w1830 and w1831;
w1833 <= not w1830 and not w1831;
w1834 <= not w1832 and not w1833;
w1835 <= b(13) and w443;
w1836 <= b(11) and w510;
w1837 <= b(12) and w438;
w1838 <= not w1836 and not w1837;
w1839 <= not w1835 and w1838;
w1840 <= w446 and w751;
w1841 <= w1839 and not w1840;
w1842 <= a(11) and not w1841;
w1843 <= a(11) and not w1842;
w1844 <= not w1841 and not w1842;
w1845 <= not w1843 and not w1844;
w1846 <= not w1834 and w1845;
w1847 <= w1834 and not w1845;
w1848 <= not w1846 and not w1847;
w1849 <= not w1755 and w1848;
w1850 <= w1755 and not w1848;
w1851 <= not w1849 and not w1850;
w1852 <= not w1754 and w1851;
w1853 <= w1754 and not w1851;
w1854 <= not w1852 and not w1853;
w1855 <= not w1743 and w1854;
w1856 <= w1743 and not w1854;
w1857 <= not w1855 and not w1856;
w1858 <= b(19) and w105;
w1859 <= b(17) and w146;
w1860 <= b(18) and w100;
w1861 <= not w1859 and not w1860;
w1862 <= not w1858 and w1861;
w1863 <= w108 and w1451;
w1864 <= w1862 and not w1863;
w1865 <= a(5) and not w1864;
w1866 <= a(5) and not w1865;
w1867 <= not w1864 and not w1865;
w1868 <= not w1866 and not w1867;
w1869 <= w1857 and not w1868;
w1870 <= w1857 and not w1869;
w1871 <= not w1868 and not w1869;
w1872 <= not w1870 and not w1871;
w1873 <= not w1708 and not w1714;
w1874 <= w1872 and w1873;
w1875 <= not w1872 and not w1873;
w1876 <= not w1874 and not w1875;
w1877 <= b(22) and w9;
w1878 <= b(20) and w27;
w1879 <= b(21) and w4;
w1880 <= not w1878 and not w1879;
w1881 <= not w1877 and w1880;
w1882 <= not w1723 and not w1725;
w1883 <= not b(21) and not b(22);
w1884 <= b(21) and b(22);
w1885 <= not w1883 and not w1884;
w1886 <= not w1882 and w1885;
w1887 <= w1882 and not w1885;
w1888 <= not w1886 and not w1887;
w1889 <= w12 and w1888;
w1890 <= w1881 and not w1889;
w1891 <= a(2) and not w1890;
w1892 <= a(2) and not w1891;
w1893 <= not w1890 and not w1891;
w1894 <= not w1892 and not w1893;
w1895 <= not w1876 and w1894;
w1896 <= w1876 and not w1894;
w1897 <= not w1895 and not w1896;
w1898 <= not w1742 and w1897;
w1899 <= w1742 and not w1897;
w1900 <= not w1898 and not w1899;
w1901 <= not w1852 and not w1855;
w1902 <= b(17) and w254;
w1903 <= b(15) and w284;
w1904 <= b(16) and w249;
w1905 <= not w1903 and not w1904;
w1906 <= not w1902 and w1905;
w1907 <= w257 and w1099;
w1908 <= w1906 and not w1907;
w1909 <= a(8) and not w1908;
w1910 <= a(8) and not w1909;
w1911 <= not w1908 and not w1909;
w1912 <= not w1910 and not w1911;
w1913 <= b(14) and w443;
w1914 <= b(12) and w510;
w1915 <= b(13) and w438;
w1916 <= not w1914 and not w1915;
w1917 <= not w1913 and w1916;
w1918 <= w446 and w777;
w1919 <= w1917 and not w1918;
w1920 <= a(11) and not w1919;
w1921 <= a(11) and not w1920;
w1922 <= not w1919 and not w1920;
w1923 <= not w1921 and not w1922;
w1924 <= not w1827 and not w1833;
w1925 <= b(11) and w694;
w1926 <= b(9) and w799;
w1927 <= b(10) and w689;
w1928 <= not w1926 and not w1927;
w1929 <= not w1925 and w1928;
w1930 <= w561 and w697;
w1931 <= w1929 and not w1930;
w1932 <= a(14) and not w1931;
w1933 <= a(14) and not w1932;
w1934 <= not w1931 and not w1932;
w1935 <= not w1933 and not w1934;
w1936 <= not w1810 and not w1813;
w1937 <= not w1781 and w1803;
w1938 <= not w1807 and not w1937;
w1939 <= b(2) and w1791;
w1940 <= w1642 and not w1790;
w1941 <= w1785 and w1940;
w1942 <= b(0) and w1941;
w1943 <= b(1) and w1786;
w1944 <= not w1942 and not w1943;
w1945 <= not w1939 and w1944;
w1946 <= w39 and w1794;
w1947 <= w1945 and not w1946;
w1948 <= a(23) and not w1947;
w1949 <= a(23) and not w1948;
w1950 <= not w1947 and not w1948;
w1951 <= not w1949 and not w1950;
w1952 <= not w1801 and w1951;
w1953 <= w1801 and not w1951;
w1954 <= not w1952 and not w1953;
w1955 <= b(5) and w1370;
w1956 <= b(3) and w1506;
w1957 <= b(4) and w1365;
w1958 <= not w1956 and not w1957;
w1959 <= not w1955 and w1958;
w1960 <= w137 and w1373;
w1961 <= w1959 and not w1960;
w1962 <= a(20) and not w1961;
w1963 <= a(20) and not w1962;
w1964 <= not w1961 and not w1962;
w1965 <= not w1963 and not w1964;
w1966 <= w1954 and not w1965;
w1967 <= not w1954 and w1965;
w1968 <= not w1938 and not w1967;
w1969 <= not w1966 and w1968;
w1970 <= not w1938 and not w1969;
w1971 <= not w1966 and not w1969;
w1972 <= not w1967 and w1971;
w1973 <= not w1970 and not w1972;
w1974 <= b(8) and w1045;
w1975 <= b(6) and w1134;
w1976 <= b(7) and w1040;
w1977 <= not w1975 and not w1976;
w1978 <= not w1974 and w1977;
w1979 <= w328 and w1048;
w1980 <= w1978 and not w1979;
w1981 <= a(17) and not w1980;
w1982 <= a(17) and not w1981;
w1983 <= not w1980 and not w1981;
w1984 <= not w1982 and not w1983;
w1985 <= w1973 and w1984;
w1986 <= not w1973 and not w1984;
w1987 <= not w1985 and not w1986;
w1988 <= not w1936 and w1987;
w1989 <= w1936 and not w1987;
w1990 <= not w1988 and not w1989;
w1991 <= w1935 and not w1990;
w1992 <= not w1935 and w1990;
w1993 <= not w1991 and not w1992;
w1994 <= not w1924 and w1993;
w1995 <= w1924 and not w1993;
w1996 <= not w1994 and not w1995;
w1997 <= not w1923 and w1996;
w1998 <= w1996 and not w1997;
w1999 <= not w1923 and not w1997;
w2000 <= not w1998 and not w1999;
w2001 <= not w1847 and not w1849;
w2002 <= not w2000 and not w2001;
w2003 <= w2000 and w2001;
w2004 <= not w2002 and not w2003;
w2005 <= not w1912 and w2004;
w2006 <= not w1912 and not w2005;
w2007 <= w2004 and not w2005;
w2008 <= not w2006 and not w2007;
w2009 <= not w1901 and not w2008;
w2010 <= not w1901 and not w2009;
w2011 <= not w2008 and not w2009;
w2012 <= not w2010 and not w2011;
w2013 <= b(20) and w105;
w2014 <= b(18) and w146;
w2015 <= b(19) and w100;
w2016 <= not w2014 and not w2015;
w2017 <= not w2013 and w2016;
w2018 <= w108 and w1589;
w2019 <= w2017 and not w2018;
w2020 <= a(5) and not w2019;
w2021 <= a(5) and not w2020;
w2022 <= not w2019 and not w2020;
w2023 <= not w2021 and not w2022;
w2024 <= not w2012 and not w2023;
w2025 <= not w2012 and not w2024;
w2026 <= not w2023 and not w2024;
w2027 <= not w2025 and not w2026;
w2028 <= not w1869 and not w1875;
w2029 <= w2027 and w2028;
w2030 <= not w2027 and not w2028;
w2031 <= not w2029 and not w2030;
w2032 <= b(23) and w9;
w2033 <= b(21) and w27;
w2034 <= b(22) and w4;
w2035 <= not w2033 and not w2034;
w2036 <= not w2032 and w2035;
w2037 <= not w1884 and not w1886;
w2038 <= not b(22) and not b(23);
w2039 <= b(22) and b(23);
w2040 <= not w2038 and not w2039;
w2041 <= not w2037 and w2040;
w2042 <= w2037 and not w2040;
w2043 <= not w2041 and not w2042;
w2044 <= w12 and w2043;
w2045 <= w2036 and not w2044;
w2046 <= a(2) and not w2045;
w2047 <= a(2) and not w2046;
w2048 <= not w2045 and not w2046;
w2049 <= not w2047 and not w2048;
w2050 <= w2031 and not w2049;
w2051 <= w2031 and not w2050;
w2052 <= not w2049 and not w2050;
w2053 <= not w2051 and not w2052;
w2054 <= not w1896 and not w1898;
w2055 <= not w2053 and not w2054;
w2056 <= w2053 and w2054;
w2057 <= not w2055 and not w2056;
w2058 <= not w2024 and not w2030;
w2059 <= b(21) and w105;
w2060 <= b(19) and w146;
w2061 <= b(20) and w100;
w2062 <= not w2060 and not w2061;
w2063 <= not w2059 and w2062;
w2064 <= w108 and w1727;
w2065 <= w2063 and not w2064;
w2066 <= a(5) and not w2065;
w2067 <= a(5) and not w2066;
w2068 <= not w2065 and not w2066;
w2069 <= not w2067 and not w2068;
w2070 <= not w2005 and not w2009;
w2071 <= b(15) and w443;
w2072 <= b(13) and w510;
w2073 <= b(14) and w438;
w2074 <= not w2072 and not w2073;
w2075 <= not w2071 and w2074;
w2076 <= w446 and w874;
w2077 <= w2075 and not w2076;
w2078 <= a(11) and not w2077;
w2079 <= a(11) and not w2078;
w2080 <= not w2077 and not w2078;
w2081 <= not w2079 and not w2080;
w2082 <= not w1992 and not w1994;
w2083 <= b(12) and w694;
w2084 <= b(10) and w799;
w2085 <= b(11) and w689;
w2086 <= not w2084 and not w2085;
w2087 <= not w2083 and w2086;
w2088 <= w585 and w697;
w2089 <= w2087 and not w2088;
w2090 <= a(14) and not w2089;
w2091 <= a(14) and not w2090;
w2092 <= not w2089 and not w2090;
w2093 <= not w2091 and not w2092;
w2094 <= not w1986 and not w1988;
w2095 <= b(6) and w1370;
w2096 <= b(4) and w1506;
w2097 <= b(5) and w1365;
w2098 <= not w2096 and not w2097;
w2099 <= not w2095 and w2098;
w2100 <= w202 and w1373;
w2101 <= w2099 and not w2100;
w2102 <= a(20) and not w2101;
w2103 <= a(20) and not w2102;
w2104 <= not w2101 and not w2102;
w2105 <= not w2103 and not w2104;
w2106 <= a(23) and not a(24);
w2107 <= not a(23) and a(24);
w2108 <= not w2106 and not w2107;
w2109 <= b(0) and not w2108;
w2110 <= not w1953 and w2109;
w2111 <= w1953 and not w2109;
w2112 <= not w2110 and not w2111;
w2113 <= b(3) and w1791;
w2114 <= b(1) and w1941;
w2115 <= b(2) and w1786;
w2116 <= not w2114 and not w2115;
w2117 <= not w2113 and w2116;
w2118 <= w61 and w1794;
w2119 <= w2117 and not w2118;
w2120 <= a(23) and not w2119;
w2121 <= a(23) and not w2120;
w2122 <= not w2119 and not w2120;
w2123 <= not w2121 and not w2122;
w2124 <= not w2112 and not w2123;
w2125 <= w2112 and w2123;
w2126 <= not w2124 and not w2125;
w2127 <= not w2105 and w2126;
w2128 <= w2126 and not w2127;
w2129 <= not w2105 and not w2127;
w2130 <= not w2128 and not w2129;
w2131 <= not w1971 and w2130;
w2132 <= w1971 and not w2130;
w2133 <= not w2131 and not w2132;
w2134 <= b(9) and w1045;
w2135 <= b(7) and w1134;
w2136 <= b(8) and w1040;
w2137 <= not w2135 and not w2136;
w2138 <= not w2134 and w2137;
w2139 <= w394 and w1048;
w2140 <= w2138 and not w2139;
w2141 <= a(17) and not w2140;
w2142 <= a(17) and not w2141;
w2143 <= not w2140 and not w2141;
w2144 <= not w2142 and not w2143;
w2145 <= not w2133 and not w2144;
w2146 <= w2133 and w2144;
w2147 <= not w2145 and not w2146;
w2148 <= not w2094 and w2147;
w2149 <= w2094 and not w2147;
w2150 <= not w2148 and not w2149;
w2151 <= w2093 and not w2150;
w2152 <= not w2093 and w2150;
w2153 <= not w2151 and not w2152;
w2154 <= not w2082 and w2153;
w2155 <= w2082 and not w2153;
w2156 <= not w2154 and not w2155;
w2157 <= not w2081 and w2156;
w2158 <= w2156 and not w2157;
w2159 <= not w2081 and not w2157;
w2160 <= not w2158 and not w2159;
w2161 <= not w1997 and not w2002;
w2162 <= w2160 and w2161;
w2163 <= not w2160 and not w2161;
w2164 <= not w2162 and not w2163;
w2165 <= b(18) and w254;
w2166 <= b(16) and w284;
w2167 <= b(17) and w249;
w2168 <= not w2166 and not w2167;
w2169 <= not w2165 and w2168;
w2170 <= w257 and w1309;
w2171 <= w2169 and not w2170;
w2172 <= a(8) and not w2171;
w2173 <= a(8) and not w2172;
w2174 <= not w2171 and not w2172;
w2175 <= not w2173 and not w2174;
w2176 <= not w2164 and w2175;
w2177 <= w2164 and not w2175;
w2178 <= not w2176 and not w2177;
w2179 <= not w2070 and w2178;
w2180 <= w2070 and not w2178;
w2181 <= not w2179 and not w2180;
w2182 <= not w2069 and w2181;
w2183 <= not w2069 and not w2182;
w2184 <= w2181 and not w2182;
w2185 <= not w2183 and not w2184;
w2186 <= not w2058 and not w2185;
w2187 <= not w2058 and not w2186;
w2188 <= not w2185 and not w2186;
w2189 <= not w2187 and not w2188;
w2190 <= b(24) and w9;
w2191 <= b(22) and w27;
w2192 <= b(23) and w4;
w2193 <= not w2191 and not w2192;
w2194 <= not w2190 and w2193;
w2195 <= not w2039 and not w2041;
w2196 <= not b(23) and not b(24);
w2197 <= b(23) and b(24);
w2198 <= not w2196 and not w2197;
w2199 <= not w2195 and w2198;
w2200 <= w2195 and not w2198;
w2201 <= not w2199 and not w2200;
w2202 <= w12 and w2201;
w2203 <= w2194 and not w2202;
w2204 <= a(2) and not w2203;
w2205 <= a(2) and not w2204;
w2206 <= not w2203 and not w2204;
w2207 <= not w2205 and not w2206;
w2208 <= not w2189 and not w2207;
w2209 <= not w2189 and not w2208;
w2210 <= not w2207 and not w2208;
w2211 <= not w2209 and not w2210;
w2212 <= not w2050 and not w2055;
w2213 <= not w2211 and not w2212;
w2214 <= w2211 and w2212;
w2215 <= not w2213 and not w2214;
w2216 <= not w2208 and not w2213;
w2217 <= b(25) and w9;
w2218 <= b(23) and w27;
w2219 <= b(24) and w4;
w2220 <= not w2218 and not w2219;
w2221 <= not w2217 and w2220;
w2222 <= not w2197 and not w2199;
w2223 <= not b(24) and not b(25);
w2224 <= b(24) and b(25);
w2225 <= not w2223 and not w2224;
w2226 <= not w2222 and w2225;
w2227 <= w2222 and not w2225;
w2228 <= not w2226 and not w2227;
w2229 <= w12 and w2228;
w2230 <= w2221 and not w2229;
w2231 <= a(2) and not w2230;
w2232 <= a(2) and not w2231;
w2233 <= not w2230 and not w2231;
w2234 <= not w2232 and not w2233;
w2235 <= not w2182 and not w2186;
w2236 <= b(16) and w443;
w2237 <= b(14) and w510;
w2238 <= b(15) and w438;
w2239 <= not w2237 and not w2238;
w2240 <= not w2236 and w2239;
w2241 <= w446 and w980;
w2242 <= w2240 and not w2241;
w2243 <= a(11) and not w2242;
w2244 <= a(11) and not w2243;
w2245 <= not w2242 and not w2243;
w2246 <= not w2244 and not w2245;
w2247 <= not w1971 and not w2130;
w2248 <= not w2127 and not w2247;
w2249 <= b(7) and w1370;
w2250 <= b(5) and w1506;
w2251 <= b(6) and w1365;
w2252 <= not w2250 and not w2251;
w2253 <= not w2249 and w2252;
w2254 <= w227 and w1373;
w2255 <= w2253 and not w2254;
w2256 <= a(20) and not w2255;
w2257 <= a(20) and not w2256;
w2258 <= not w2255 and not w2256;
w2259 <= not w2257 and not w2258;
w2260 <= w1953 and w2109;
w2261 <= not w2124 and not w2260;
w2262 <= b(4) and w1791;
w2263 <= b(2) and w1941;
w2264 <= b(3) and w1786;
w2265 <= not w2263 and not w2264;
w2266 <= not w2262 and w2265;
w2267 <= w89 and w1794;
w2268 <= w2266 and not w2267;
w2269 <= a(23) and not w2268;
w2270 <= a(23) and not w2269;
w2271 <= not w2268 and not w2269;
w2272 <= not w2270 and not w2271;
w2273 <= a(26) and not w2109;
w2274 <= not a(24) and a(25);
w2275 <= a(24) and not a(25);
w2276 <= not w2274 and not w2275;
w2277 <= w2108 and not w2276;
w2278 <= b(0) and w2277;
w2279 <= not a(25) and a(26);
w2280 <= a(25) and not a(26);
w2281 <= not w2279 and not w2280;
w2282 <= not w2108 and w2281;
w2283 <= b(1) and w2282;
w2284 <= not w2278 and not w2283;
w2285 <= not w2108 and not w2281;
w2286 <= not w15 and w2285;
w2287 <= w2284 and not w2286;
w2288 <= a(26) and not w2287;
w2289 <= a(26) and not w2288;
w2290 <= not w2287 and not w2288;
w2291 <= not w2289 and not w2290;
w2292 <= w2273 and not w2291;
w2293 <= not w2273 and w2291;
w2294 <= not w2292 and not w2293;
w2295 <= w2272 and w2294;
w2296 <= not w2272 and not w2294;
w2297 <= not w2295 and not w2296;
w2298 <= not w2261 and not w2297;
w2299 <= w2261 and w2297;
w2300 <= not w2298 and not w2299;
w2301 <= not w2259 and w2300;
w2302 <= w2259 and not w2300;
w2303 <= not w2301 and not w2302;
w2304 <= not w2248 and w2303;
w2305 <= w2248 and not w2303;
w2306 <= not w2304 and not w2305;
w2307 <= b(10) and w1045;
w2308 <= b(8) and w1134;
w2309 <= b(9) and w1040;
w2310 <= not w2308 and not w2309;
w2311 <= not w2307 and w2310;
w2312 <= w481 and w1048;
w2313 <= w2311 and not w2312;
w2314 <= a(17) and not w2313;
w2315 <= a(17) and not w2314;
w2316 <= not w2313 and not w2314;
w2317 <= not w2315 and not w2316;
w2318 <= w2306 and not w2317;
w2319 <= w2306 and not w2318;
w2320 <= not w2317 and not w2318;
w2321 <= not w2319 and not w2320;
w2322 <= not w2145 and not w2148;
w2323 <= w2321 and w2322;
w2324 <= not w2321 and not w2322;
w2325 <= not w2323 and not w2324;
w2326 <= b(13) and w694;
w2327 <= b(11) and w799;
w2328 <= b(12) and w689;
w2329 <= not w2327 and not w2328;
w2330 <= not w2326 and w2329;
w2331 <= w697 and w751;
w2332 <= w2330 and not w2331;
w2333 <= a(14) and not w2332;
w2334 <= a(14) and not w2333;
w2335 <= not w2332 and not w2333;
w2336 <= not w2334 and not w2335;
w2337 <= not w2325 and w2336;
w2338 <= w2325 and not w2336;
w2339 <= not w2337 and not w2338;
w2340 <= not w2152 and not w2154;
w2341 <= w2339 and not w2340;
w2342 <= not w2339 and w2340;
w2343 <= not w2341 and not w2342;
w2344 <= not w2246 and w2343;
w2345 <= w2343 and not w2344;
w2346 <= not w2246 and not w2344;
w2347 <= not w2345 and not w2346;
w2348 <= not w2157 and not w2163;
w2349 <= w2347 and w2348;
w2350 <= not w2347 and not w2348;
w2351 <= not w2349 and not w2350;
w2352 <= b(19) and w254;
w2353 <= b(17) and w284;
w2354 <= b(18) and w249;
w2355 <= not w2353 and not w2354;
w2356 <= not w2352 and w2355;
w2357 <= w257 and w1451;
w2358 <= w2356 and not w2357;
w2359 <= a(8) and not w2358;
w2360 <= a(8) and not w2359;
w2361 <= not w2358 and not w2359;
w2362 <= not w2360 and not w2361;
w2363 <= w2351 and not w2362;
w2364 <= w2351 and not w2363;
w2365 <= not w2362 and not w2363;
w2366 <= not w2364 and not w2365;
w2367 <= not w2177 and not w2179;
w2368 <= not w2366 and not w2367;
w2369 <= not w2366 and not w2368;
w2370 <= not w2367 and not w2368;
w2371 <= not w2369 and not w2370;
w2372 <= b(22) and w105;
w2373 <= b(20) and w146;
w2374 <= b(21) and w100;
w2375 <= not w2373 and not w2374;
w2376 <= not w2372 and w2375;
w2377 <= w108 and w1888;
w2378 <= w2376 and not w2377;
w2379 <= a(5) and not w2378;
w2380 <= a(5) and not w2379;
w2381 <= not w2378 and not w2379;
w2382 <= not w2380 and not w2381;
w2383 <= not w2371 and w2382;
w2384 <= w2371 and not w2382;
w2385 <= not w2383 and not w2384;
w2386 <= not w2235 and not w2385;
w2387 <= w2235 and w2385;
w2388 <= not w2386 and not w2387;
w2389 <= not w2234 and w2388;
w2390 <= w2234 and not w2388;
w2391 <= not w2389 and not w2390;
w2392 <= not w2216 and w2391;
w2393 <= w2216 and not w2391;
w2394 <= not w2392 and not w2393;
w2395 <= not w2389 and not w2392;
w2396 <= not w2371 and not w2382;
w2397 <= not w2386 and not w2396;
w2398 <= not w2344 and not w2350;
w2399 <= not w2338 and not w2341;
w2400 <= b(14) and w694;
w2401 <= b(12) and w799;
w2402 <= b(13) and w689;
w2403 <= not w2401 and not w2402;
w2404 <= not w2400 and w2403;
w2405 <= w697 and w777;
w2406 <= w2404 and not w2405;
w2407 <= a(14) and not w2406;
w2408 <= a(14) and not w2407;
w2409 <= not w2406 and not w2407;
w2410 <= not w2408 and not w2409;
w2411 <= not w2318 and not w2324;
w2412 <= b(11) and w1045;
w2413 <= b(9) and w1134;
w2414 <= b(10) and w1040;
w2415 <= not w2413 and not w2414;
w2416 <= not w2412 and w2415;
w2417 <= w561 and w1048;
w2418 <= w2416 and not w2417;
w2419 <= a(17) and not w2418;
w2420 <= a(17) and not w2419;
w2421 <= not w2418 and not w2419;
w2422 <= not w2420 and not w2421;
w2423 <= not w2301 and not w2304;
w2424 <= not w2272 and w2294;
w2425 <= not w2298 and not w2424;
w2426 <= b(2) and w2282;
w2427 <= w2108 and not w2281;
w2428 <= w2276 and w2427;
w2429 <= b(0) and w2428;
w2430 <= b(1) and w2277;
w2431 <= not w2429 and not w2430;
w2432 <= not w2426 and w2431;
w2433 <= w39 and w2285;
w2434 <= w2432 and not w2433;
w2435 <= a(26) and not w2434;
w2436 <= a(26) and not w2435;
w2437 <= not w2434 and not w2435;
w2438 <= not w2436 and not w2437;
w2439 <= not w2292 and w2438;
w2440 <= w2292 and not w2438;
w2441 <= not w2439 and not w2440;
w2442 <= b(5) and w1791;
w2443 <= b(3) and w1941;
w2444 <= b(4) and w1786;
w2445 <= not w2443 and not w2444;
w2446 <= not w2442 and w2445;
w2447 <= w137 and w1794;
w2448 <= w2446 and not w2447;
w2449 <= a(23) and not w2448;
w2450 <= a(23) and not w2449;
w2451 <= not w2448 and not w2449;
w2452 <= not w2450 and not w2451;
w2453 <= w2441 and not w2452;
w2454 <= not w2441 and w2452;
w2455 <= not w2425 and not w2454;
w2456 <= not w2453 and w2455;
w2457 <= not w2425 and not w2456;
w2458 <= not w2453 and not w2456;
w2459 <= not w2454 and w2458;
w2460 <= not w2457 and not w2459;
w2461 <= b(8) and w1370;
w2462 <= b(6) and w1506;
w2463 <= b(7) and w1365;
w2464 <= not w2462 and not w2463;
w2465 <= not w2461 and w2464;
w2466 <= w328 and w1373;
w2467 <= w2465 and not w2466;
w2468 <= a(20) and not w2467;
w2469 <= a(20) and not w2468;
w2470 <= not w2467 and not w2468;
w2471 <= not w2469 and not w2470;
w2472 <= w2460 and w2471;
w2473 <= not w2460 and not w2471;
w2474 <= not w2472 and not w2473;
w2475 <= not w2423 and w2474;
w2476 <= w2423 and not w2474;
w2477 <= not w2475 and not w2476;
w2478 <= w2422 and not w2477;
w2479 <= not w2422 and w2477;
w2480 <= not w2478 and not w2479;
w2481 <= not w2411 and w2480;
w2482 <= w2411 and not w2480;
w2483 <= not w2481 and not w2482;
w2484 <= not w2410 and w2483;
w2485 <= w2483 and not w2484;
w2486 <= not w2410 and not w2484;
w2487 <= not w2485 and not w2486;
w2488 <= not w2399 and w2487;
w2489 <= w2399 and not w2487;
w2490 <= not w2488 and not w2489;
w2491 <= b(17) and w443;
w2492 <= b(15) and w510;
w2493 <= b(16) and w438;
w2494 <= not w2492 and not w2493;
w2495 <= not w2491 and w2494;
w2496 <= w446 and w1099;
w2497 <= w2495 and not w2496;
w2498 <= a(11) and not w2497;
w2499 <= a(11) and not w2498;
w2500 <= not w2497 and not w2498;
w2501 <= not w2499 and not w2500;
w2502 <= not w2490 and not w2501;
w2503 <= w2490 and w2501;
w2504 <= not w2502 and not w2503;
w2505 <= w2398 and not w2504;
w2506 <= not w2398 and w2504;
w2507 <= not w2505 and not w2506;
w2508 <= b(20) and w254;
w2509 <= b(18) and w284;
w2510 <= b(19) and w249;
w2511 <= not w2509 and not w2510;
w2512 <= not w2508 and w2511;
w2513 <= w257 and w1589;
w2514 <= w2512 and not w2513;
w2515 <= a(8) and not w2514;
w2516 <= a(8) and not w2515;
w2517 <= not w2514 and not w2515;
w2518 <= not w2516 and not w2517;
w2519 <= w2507 and not w2518;
w2520 <= w2507 and not w2519;
w2521 <= not w2518 and not w2519;
w2522 <= not w2520 and not w2521;
w2523 <= not w2363 and not w2368;
w2524 <= w2522 and w2523;
w2525 <= not w2522 and not w2523;
w2526 <= not w2524 and not w2525;
w2527 <= b(23) and w105;
w2528 <= b(21) and w146;
w2529 <= b(22) and w100;
w2530 <= not w2528 and not w2529;
w2531 <= not w2527 and w2530;
w2532 <= w108 and w2043;
w2533 <= w2531 and not w2532;
w2534 <= a(5) and not w2533;
w2535 <= a(5) and not w2534;
w2536 <= not w2533 and not w2534;
w2537 <= not w2535 and not w2536;
w2538 <= w2526 and not w2537;
w2539 <= w2526 and not w2538;
w2540 <= not w2537 and not w2538;
w2541 <= not w2539 and not w2540;
w2542 <= not w2397 and w2541;
w2543 <= w2397 and not w2541;
w2544 <= not w2542 and not w2543;
w2545 <= b(26) and w9;
w2546 <= b(24) and w27;
w2547 <= b(25) and w4;
w2548 <= not w2546 and not w2547;
w2549 <= not w2545 and w2548;
w2550 <= not w2224 and not w2226;
w2551 <= not b(25) and not b(26);
w2552 <= b(25) and b(26);
w2553 <= not w2551 and not w2552;
w2554 <= not w2550 and w2553;
w2555 <= w2550 and not w2553;
w2556 <= not w2554 and not w2555;
w2557 <= w12 and w2556;
w2558 <= w2549 and not w2557;
w2559 <= a(2) and not w2558;
w2560 <= a(2) and not w2559;
w2561 <= not w2558 and not w2559;
w2562 <= not w2560 and not w2561;
w2563 <= not w2544 and not w2562;
w2564 <= w2544 and w2562;
w2565 <= not w2563 and not w2564;
w2566 <= not w2395 and w2565;
w2567 <= w2395 and not w2565;
w2568 <= not w2566 and not w2567;
w2569 <= not w2563 and not w2566;
w2570 <= b(24) and w105;
w2571 <= b(22) and w146;
w2572 <= b(23) and w100;
w2573 <= not w2571 and not w2572;
w2574 <= not w2570 and w2573;
w2575 <= w108 and w2201;
w2576 <= w2574 and not w2575;
w2577 <= a(5) and not w2576;
w2578 <= a(5) and not w2577;
w2579 <= not w2576 and not w2577;
w2580 <= not w2578 and not w2579;
w2581 <= b(15) and w694;
w2582 <= b(13) and w799;
w2583 <= b(14) and w689;
w2584 <= not w2582 and not w2583;
w2585 <= not w2581 and w2584;
w2586 <= w697 and w874;
w2587 <= w2585 and not w2586;
w2588 <= a(14) and not w2587;
w2589 <= a(14) and not w2588;
w2590 <= not w2587 and not w2588;
w2591 <= not w2589 and not w2590;
w2592 <= not w2479 and not w2481;
w2593 <= b(12) and w1045;
w2594 <= b(10) and w1134;
w2595 <= b(11) and w1040;
w2596 <= not w2594 and not w2595;
w2597 <= not w2593 and w2596;
w2598 <= w585 and w1048;
w2599 <= w2597 and not w2598;
w2600 <= a(17) and not w2599;
w2601 <= a(17) and not w2600;
w2602 <= not w2599 and not w2600;
w2603 <= not w2601 and not w2602;
w2604 <= not w2473 and not w2475;
w2605 <= b(6) and w1791;
w2606 <= b(4) and w1941;
w2607 <= b(5) and w1786;
w2608 <= not w2606 and not w2607;
w2609 <= not w2605 and w2608;
w2610 <= w202 and w1794;
w2611 <= w2609 and not w2610;
w2612 <= a(23) and not w2611;
w2613 <= a(23) and not w2612;
w2614 <= not w2611 and not w2612;
w2615 <= not w2613 and not w2614;
w2616 <= a(26) and not a(27);
w2617 <= not a(26) and a(27);
w2618 <= not w2616 and not w2617;
w2619 <= b(0) and not w2618;
w2620 <= not w2440 and w2619;
w2621 <= w2440 and not w2619;
w2622 <= not w2620 and not w2621;
w2623 <= b(3) and w2282;
w2624 <= b(1) and w2428;
w2625 <= b(2) and w2277;
w2626 <= not w2624 and not w2625;
w2627 <= not w2623 and w2626;
w2628 <= w61 and w2285;
w2629 <= w2627 and not w2628;
w2630 <= a(26) and not w2629;
w2631 <= a(26) and not w2630;
w2632 <= not w2629 and not w2630;
w2633 <= not w2631 and not w2632;
w2634 <= not w2622 and not w2633;
w2635 <= w2622 and w2633;
w2636 <= not w2634 and not w2635;
w2637 <= not w2615 and w2636;
w2638 <= w2636 and not w2637;
w2639 <= not w2615 and not w2637;
w2640 <= not w2638 and not w2639;
w2641 <= not w2458 and w2640;
w2642 <= w2458 and not w2640;
w2643 <= not w2641 and not w2642;
w2644 <= b(9) and w1370;
w2645 <= b(7) and w1506;
w2646 <= b(8) and w1365;
w2647 <= not w2645 and not w2646;
w2648 <= not w2644 and w2647;
w2649 <= w394 and w1373;
w2650 <= w2648 and not w2649;
w2651 <= a(20) and not w2650;
w2652 <= a(20) and not w2651;
w2653 <= not w2650 and not w2651;
w2654 <= not w2652 and not w2653;
w2655 <= not w2643 and not w2654;
w2656 <= w2643 and w2654;
w2657 <= not w2655 and not w2656;
w2658 <= not w2604 and w2657;
w2659 <= w2604 and not w2657;
w2660 <= not w2658 and not w2659;
w2661 <= w2603 and not w2660;
w2662 <= not w2603 and w2660;
w2663 <= not w2661 and not w2662;
w2664 <= not w2592 and w2663;
w2665 <= w2592 and not w2663;
w2666 <= not w2664 and not w2665;
w2667 <= not w2591 and w2666;
w2668 <= w2666 and not w2667;
w2669 <= not w2591 and not w2667;
w2670 <= not w2668 and not w2669;
w2671 <= not w2399 and not w2487;
w2672 <= not w2484 and not w2671;
w2673 <= w2670 and w2672;
w2674 <= not w2670 and not w2672;
w2675 <= not w2673 and not w2674;
w2676 <= b(18) and w443;
w2677 <= b(16) and w510;
w2678 <= b(17) and w438;
w2679 <= not w2677 and not w2678;
w2680 <= not w2676 and w2679;
w2681 <= w446 and w1309;
w2682 <= w2680 and not w2681;
w2683 <= a(11) and not w2682;
w2684 <= a(11) and not w2683;
w2685 <= not w2682 and not w2683;
w2686 <= not w2684 and not w2685;
w2687 <= w2675 and not w2686;
w2688 <= w2675 and not w2687;
w2689 <= not w2686 and not w2687;
w2690 <= not w2688 and not w2689;
w2691 <= not w2502 and not w2506;
w2692 <= w2690 and w2691;
w2693 <= not w2690 and not w2691;
w2694 <= not w2692 and not w2693;
w2695 <= b(21) and w254;
w2696 <= b(19) and w284;
w2697 <= b(20) and w249;
w2698 <= not w2696 and not w2697;
w2699 <= not w2695 and w2698;
w2700 <= w257 and w1727;
w2701 <= w2699 and not w2700;
w2702 <= a(8) and not w2701;
w2703 <= a(8) and not w2702;
w2704 <= not w2701 and not w2702;
w2705 <= not w2703 and not w2704;
w2706 <= not w2694 and w2705;
w2707 <= w2694 and not w2705;
w2708 <= not w2706 and not w2707;
w2709 <= not w2519 and not w2525;
w2710 <= w2708 and not w2709;
w2711 <= not w2708 and w2709;
w2712 <= not w2710 and not w2711;
w2713 <= not w2580 and w2712;
w2714 <= w2712 and not w2713;
w2715 <= not w2580 and not w2713;
w2716 <= not w2714 and not w2715;
w2717 <= not w2397 and not w2541;
w2718 <= not w2538 and not w2717;
w2719 <= w2716 and w2718;
w2720 <= not w2716 and not w2718;
w2721 <= not w2719 and not w2720;
w2722 <= b(27) and w9;
w2723 <= b(25) and w27;
w2724 <= b(26) and w4;
w2725 <= not w2723 and not w2724;
w2726 <= not w2722 and w2725;
w2727 <= not w2552 and not w2554;
w2728 <= not b(26) and not b(27);
w2729 <= b(26) and b(27);
w2730 <= not w2728 and not w2729;
w2731 <= not w2727 and w2730;
w2732 <= w2727 and not w2730;
w2733 <= not w2731 and not w2732;
w2734 <= w12 and w2733;
w2735 <= w2726 and not w2734;
w2736 <= a(2) and not w2735;
w2737 <= a(2) and not w2736;
w2738 <= not w2735 and not w2736;
w2739 <= not w2737 and not w2738;
w2740 <= not w2721 and w2739;
w2741 <= w2721 and not w2739;
w2742 <= not w2740 and not w2741;
w2743 <= not w2569 and w2742;
w2744 <= w2569 and not w2742;
w2745 <= not w2743 and not w2744;
w2746 <= not w2741 and not w2743;
w2747 <= b(25) and w105;
w2748 <= b(23) and w146;
w2749 <= b(24) and w100;
w2750 <= not w2748 and not w2749;
w2751 <= not w2747 and w2750;
w2752 <= w108 and w2228;
w2753 <= w2751 and not w2752;
w2754 <= a(5) and not w2753;
w2755 <= a(5) and not w2754;
w2756 <= not w2753 and not w2754;
w2757 <= not w2755 and not w2756;
w2758 <= not w2458 and not w2640;
w2759 <= not w2637 and not w2758;
w2760 <= b(7) and w1791;
w2761 <= b(5) and w1941;
w2762 <= b(6) and w1786;
w2763 <= not w2761 and not w2762;
w2764 <= not w2760 and w2763;
w2765 <= w227 and w1794;
w2766 <= w2764 and not w2765;
w2767 <= a(23) and not w2766;
w2768 <= a(23) and not w2767;
w2769 <= not w2766 and not w2767;
w2770 <= not w2768 and not w2769;
w2771 <= w2440 and w2619;
w2772 <= not w2634 and not w2771;
w2773 <= b(4) and w2282;
w2774 <= b(2) and w2428;
w2775 <= b(3) and w2277;
w2776 <= not w2774 and not w2775;
w2777 <= not w2773 and w2776;
w2778 <= w89 and w2285;
w2779 <= w2777 and not w2778;
w2780 <= a(26) and not w2779;
w2781 <= a(26) and not w2780;
w2782 <= not w2779 and not w2780;
w2783 <= not w2781 and not w2782;
w2784 <= a(29) and not w2619;
w2785 <= not a(27) and a(28);
w2786 <= a(27) and not a(28);
w2787 <= not w2785 and not w2786;
w2788 <= w2618 and not w2787;
w2789 <= b(0) and w2788;
w2790 <= not a(28) and a(29);
w2791 <= a(28) and not a(29);
w2792 <= not w2790 and not w2791;
w2793 <= not w2618 and w2792;
w2794 <= b(1) and w2793;
w2795 <= not w2789 and not w2794;
w2796 <= not w2618 and not w2792;
w2797 <= not w15 and w2796;
w2798 <= w2795 and not w2797;
w2799 <= a(29) and not w2798;
w2800 <= a(29) and not w2799;
w2801 <= not w2798 and not w2799;
w2802 <= not w2800 and not w2801;
w2803 <= w2784 and not w2802;
w2804 <= not w2784 and w2802;
w2805 <= not w2803 and not w2804;
w2806 <= w2783 and w2805;
w2807 <= not w2783 and not w2805;
w2808 <= not w2806 and not w2807;
w2809 <= not w2772 and not w2808;
w2810 <= w2772 and w2808;
w2811 <= not w2809 and not w2810;
w2812 <= not w2770 and w2811;
w2813 <= w2770 and not w2811;
w2814 <= not w2812 and not w2813;
w2815 <= not w2759 and w2814;
w2816 <= w2759 and not w2814;
w2817 <= not w2815 and not w2816;
w2818 <= b(10) and w1370;
w2819 <= b(8) and w1506;
w2820 <= b(9) and w1365;
w2821 <= not w2819 and not w2820;
w2822 <= not w2818 and w2821;
w2823 <= w481 and w1373;
w2824 <= w2822 and not w2823;
w2825 <= a(20) and not w2824;
w2826 <= a(20) and not w2825;
w2827 <= not w2824 and not w2825;
w2828 <= not w2826 and not w2827;
w2829 <= w2817 and not w2828;
w2830 <= w2817 and not w2829;
w2831 <= not w2828 and not w2829;
w2832 <= not w2830 and not w2831;
w2833 <= not w2655 and not w2658;
w2834 <= w2832 and w2833;
w2835 <= not w2832 and not w2833;
w2836 <= not w2834 and not w2835;
w2837 <= b(13) and w1045;
w2838 <= b(11) and w1134;
w2839 <= b(12) and w1040;
w2840 <= not w2838 and not w2839;
w2841 <= not w2837 and w2840;
w2842 <= w751 and w1048;
w2843 <= w2841 and not w2842;
w2844 <= a(17) and not w2843;
w2845 <= a(17) and not w2844;
w2846 <= not w2843 and not w2844;
w2847 <= not w2845 and not w2846;
w2848 <= w2836 and not w2847;
w2849 <= w2836 and not w2848;
w2850 <= not w2847 and not w2848;
w2851 <= not w2849 and not w2850;
w2852 <= not w2662 and not w2664;
w2853 <= not w2851 and not w2852;
w2854 <= not w2851 and not w2853;
w2855 <= not w2852 and not w2853;
w2856 <= not w2854 and not w2855;
w2857 <= b(16) and w694;
w2858 <= b(14) and w799;
w2859 <= b(15) and w689;
w2860 <= not w2858 and not w2859;
w2861 <= not w2857 and w2860;
w2862 <= w697 and w980;
w2863 <= w2861 and not w2862;
w2864 <= a(14) and not w2863;
w2865 <= a(14) and not w2864;
w2866 <= not w2863 and not w2864;
w2867 <= not w2865 and not w2866;
w2868 <= not w2856 and not w2867;
w2869 <= not w2856 and not w2868;
w2870 <= not w2867 and not w2868;
w2871 <= not w2869 and not w2870;
w2872 <= not w2667 and not w2674;
w2873 <= w2871 and w2872;
w2874 <= not w2871 and not w2872;
w2875 <= not w2873 and not w2874;
w2876 <= b(19) and w443;
w2877 <= b(17) and w510;
w2878 <= b(18) and w438;
w2879 <= not w2877 and not w2878;
w2880 <= not w2876 and w2879;
w2881 <= w446 and w1451;
w2882 <= w2880 and not w2881;
w2883 <= a(11) and not w2882;
w2884 <= a(11) and not w2883;
w2885 <= not w2882 and not w2883;
w2886 <= not w2884 and not w2885;
w2887 <= w2875 and not w2886;
w2888 <= w2875 and not w2887;
w2889 <= not w2886 and not w2887;
w2890 <= not w2888 and not w2889;
w2891 <= not w2687 and not w2693;
w2892 <= w2890 and w2891;
w2893 <= not w2890 and not w2891;
w2894 <= not w2892 and not w2893;
w2895 <= b(22) and w254;
w2896 <= b(20) and w284;
w2897 <= b(21) and w249;
w2898 <= not w2896 and not w2897;
w2899 <= not w2895 and w2898;
w2900 <= w257 and w1888;
w2901 <= w2899 and not w2900;
w2902 <= a(8) and not w2901;
w2903 <= a(8) and not w2902;
w2904 <= not w2901 and not w2902;
w2905 <= not w2903 and not w2904;
w2906 <= not w2894 and w2905;
w2907 <= w2894 and not w2905;
w2908 <= not w2906 and not w2907;
w2909 <= not w2707 and not w2710;
w2910 <= w2908 and not w2909;
w2911 <= not w2908 and w2909;
w2912 <= not w2910 and not w2911;
w2913 <= not w2757 and w2912;
w2914 <= w2912 and not w2913;
w2915 <= not w2757 and not w2913;
w2916 <= not w2914 and not w2915;
w2917 <= not w2713 and not w2720;
w2918 <= w2916 and w2917;
w2919 <= not w2916 and not w2917;
w2920 <= not w2918 and not w2919;
w2921 <= b(28) and w9;
w2922 <= b(26) and w27;
w2923 <= b(27) and w4;
w2924 <= not w2922 and not w2923;
w2925 <= not w2921 and w2924;
w2926 <= not w2729 and not w2731;
w2927 <= not b(27) and not b(28);
w2928 <= b(27) and b(28);
w2929 <= not w2927 and not w2928;
w2930 <= not w2926 and w2929;
w2931 <= w2926 and not w2929;
w2932 <= not w2930 and not w2931;
w2933 <= w12 and w2932;
w2934 <= w2925 and not w2933;
w2935 <= a(2) and not w2934;
w2936 <= a(2) and not w2935;
w2937 <= not w2934 and not w2935;
w2938 <= not w2936 and not w2937;
w2939 <= not w2920 and w2938;
w2940 <= w2920 and not w2938;
w2941 <= not w2939 and not w2940;
w2942 <= not w2746 and w2941;
w2943 <= w2746 and not w2941;
w2944 <= not w2942 and not w2943;
w2945 <= not w2913 and not w2919;
w2946 <= b(26) and w105;
w2947 <= b(24) and w146;
w2948 <= b(25) and w100;
w2949 <= not w2947 and not w2948;
w2950 <= not w2946 and w2949;
w2951 <= w108 and w2556;
w2952 <= w2950 and not w2951;
w2953 <= a(5) and not w2952;
w2954 <= a(5) and not w2953;
w2955 <= not w2952 and not w2953;
w2956 <= not w2954 and not w2955;
w2957 <= not w2887 and not w2893;
w2958 <= b(14) and w1045;
w2959 <= b(12) and w1134;
w2960 <= b(13) and w1040;
w2961 <= not w2959 and not w2960;
w2962 <= not w2958 and w2961;
w2963 <= w777 and w1048;
w2964 <= w2962 and not w2963;
w2965 <= a(17) and not w2964;
w2966 <= a(17) and not w2965;
w2967 <= not w2964 and not w2965;
w2968 <= not w2966 and not w2967;
w2969 <= not w2829 and not w2835;
w2970 <= b(11) and w1370;
w2971 <= b(9) and w1506;
w2972 <= b(10) and w1365;
w2973 <= not w2971 and not w2972;
w2974 <= not w2970 and w2973;
w2975 <= w561 and w1373;
w2976 <= w2974 and not w2975;
w2977 <= a(20) and not w2976;
w2978 <= a(20) and not w2977;
w2979 <= not w2976 and not w2977;
w2980 <= not w2978 and not w2979;
w2981 <= not w2812 and not w2815;
w2982 <= not w2783 and w2805;
w2983 <= not w2809 and not w2982;
w2984 <= b(2) and w2793;
w2985 <= w2618 and not w2792;
w2986 <= w2787 and w2985;
w2987 <= b(0) and w2986;
w2988 <= b(1) and w2788;
w2989 <= not w2987 and not w2988;
w2990 <= not w2984 and w2989;
w2991 <= w39 and w2796;
w2992 <= w2990 and not w2991;
w2993 <= a(29) and not w2992;
w2994 <= a(29) and not w2993;
w2995 <= not w2992 and not w2993;
w2996 <= not w2994 and not w2995;
w2997 <= not w2803 and w2996;
w2998 <= w2803 and not w2996;
w2999 <= not w2997 and not w2998;
w3000 <= b(5) and w2282;
w3001 <= b(3) and w2428;
w3002 <= b(4) and w2277;
w3003 <= not w3001 and not w3002;
w3004 <= not w3000 and w3003;
w3005 <= w137 and w2285;
w3006 <= w3004 and not w3005;
w3007 <= a(26) and not w3006;
w3008 <= a(26) and not w3007;
w3009 <= not w3006 and not w3007;
w3010 <= not w3008 and not w3009;
w3011 <= w2999 and not w3010;
w3012 <= not w2999 and w3010;
w3013 <= not w2983 and not w3012;
w3014 <= not w3011 and w3013;
w3015 <= not w2983 and not w3014;
w3016 <= not w3011 and not w3014;
w3017 <= not w3012 and w3016;
w3018 <= not w3015 and not w3017;
w3019 <= b(8) and w1791;
w3020 <= b(6) and w1941;
w3021 <= b(7) and w1786;
w3022 <= not w3020 and not w3021;
w3023 <= not w3019 and w3022;
w3024 <= w328 and w1794;
w3025 <= w3023 and not w3024;
w3026 <= a(23) and not w3025;
w3027 <= a(23) and not w3026;
w3028 <= not w3025 and not w3026;
w3029 <= not w3027 and not w3028;
w3030 <= w3018 and w3029;
w3031 <= not w3018 and not w3029;
w3032 <= not w3030 and not w3031;
w3033 <= not w2981 and w3032;
w3034 <= w2981 and not w3032;
w3035 <= not w3033 and not w3034;
w3036 <= w2980 and not w3035;
w3037 <= not w2980 and w3035;
w3038 <= not w3036 and not w3037;
w3039 <= not w2969 and w3038;
w3040 <= w2969 and not w3038;
w3041 <= not w3039 and not w3040;
w3042 <= not w2968 and w3041;
w3043 <= w3041 and not w3042;
w3044 <= not w2968 and not w3042;
w3045 <= not w3043 and not w3044;
w3046 <= not w2848 and not w2853;
w3047 <= w3045 and w3046;
w3048 <= not w3045 and not w3046;
w3049 <= not w3047 and not w3048;
w3050 <= b(17) and w694;
w3051 <= b(15) and w799;
w3052 <= b(16) and w689;
w3053 <= not w3051 and not w3052;
w3054 <= not w3050 and w3053;
w3055 <= w697 and w1099;
w3056 <= w3054 and not w3055;
w3057 <= a(14) and not w3056;
w3058 <= a(14) and not w3057;
w3059 <= not w3056 and not w3057;
w3060 <= not w3058 and not w3059;
w3061 <= w3049 and not w3060;
w3062 <= w3049 and not w3061;
w3063 <= not w3060 and not w3061;
w3064 <= not w3062 and not w3063;
w3065 <= not w2868 and not w2874;
w3066 <= w3064 and w3065;
w3067 <= not w3064 and not w3065;
w3068 <= not w3066 and not w3067;
w3069 <= b(20) and w443;
w3070 <= b(18) and w510;
w3071 <= b(19) and w438;
w3072 <= not w3070 and not w3071;
w3073 <= not w3069 and w3072;
w3074 <= w446 and w1589;
w3075 <= w3073 and not w3074;
w3076 <= a(11) and not w3075;
w3077 <= a(11) and not w3076;
w3078 <= not w3075 and not w3076;
w3079 <= not w3077 and not w3078;
w3080 <= w3068 and not w3079;
w3081 <= not w3068 and w3079;
w3082 <= not w2957 and not w3081;
w3083 <= not w3080 and w3082;
w3084 <= not w2957 and not w3083;
w3085 <= not w3080 and not w3083;
w3086 <= not w3081 and w3085;
w3087 <= not w3084 and not w3086;
w3088 <= b(23) and w254;
w3089 <= b(21) and w284;
w3090 <= b(22) and w249;
w3091 <= not w3089 and not w3090;
w3092 <= not w3088 and w3091;
w3093 <= w257 and w2043;
w3094 <= w3092 and not w3093;
w3095 <= a(8) and not w3094;
w3096 <= a(8) and not w3095;
w3097 <= not w3094 and not w3095;
w3098 <= not w3096 and not w3097;
w3099 <= not w3087 and not w3098;
w3100 <= not w3087 and not w3099;
w3101 <= not w3098 and not w3099;
w3102 <= not w3100 and not w3101;
w3103 <= not w2907 and not w2910;
w3104 <= not w3102 and not w3103;
w3105 <= w3102 and w3103;
w3106 <= not w3104 and not w3105;
w3107 <= not w2956 and w3106;
w3108 <= not w2956 and not w3107;
w3109 <= w3106 and not w3107;
w3110 <= not w3108 and not w3109;
w3111 <= not w2945 and not w3110;
w3112 <= not w2945 and not w3111;
w3113 <= not w3110 and not w3111;
w3114 <= not w3112 and not w3113;
w3115 <= b(29) and w9;
w3116 <= b(27) and w27;
w3117 <= b(28) and w4;
w3118 <= not w3116 and not w3117;
w3119 <= not w3115 and w3118;
w3120 <= not w2928 and not w2930;
w3121 <= not b(28) and not b(29);
w3122 <= b(28) and b(29);
w3123 <= not w3121 and not w3122;
w3124 <= not w3120 and w3123;
w3125 <= w3120 and not w3123;
w3126 <= not w3124 and not w3125;
w3127 <= w12 and w3126;
w3128 <= w3119 and not w3127;
w3129 <= a(2) and not w3128;
w3130 <= a(2) and not w3129;
w3131 <= not w3128 and not w3129;
w3132 <= not w3130 and not w3131;
w3133 <= not w3114 and not w3132;
w3134 <= not w3114 and not w3133;
w3135 <= not w3132 and not w3133;
w3136 <= not w3134 and not w3135;
w3137 <= not w2940 and not w2942;
w3138 <= not w3136 and not w3137;
w3139 <= w3136 and w3137;
w3140 <= not w3138 and not w3139;
w3141 <= not w3099 and not w3104;
w3142 <= b(15) and w1045;
w3143 <= b(13) and w1134;
w3144 <= b(14) and w1040;
w3145 <= not w3143 and not w3144;
w3146 <= not w3142 and w3145;
w3147 <= w874 and w1048;
w3148 <= w3146 and not w3147;
w3149 <= a(17) and not w3148;
w3150 <= a(17) and not w3149;
w3151 <= not w3148 and not w3149;
w3152 <= not w3150 and not w3151;
w3153 <= not w3037 and not w3039;
w3154 <= b(12) and w1370;
w3155 <= b(10) and w1506;
w3156 <= b(11) and w1365;
w3157 <= not w3155 and not w3156;
w3158 <= not w3154 and w3157;
w3159 <= w585 and w1373;
w3160 <= w3158 and not w3159;
w3161 <= a(20) and not w3160;
w3162 <= a(20) and not w3161;
w3163 <= not w3160 and not w3161;
w3164 <= not w3162 and not w3163;
w3165 <= not w3031 and not w3033;
w3166 <= b(6) and w2282;
w3167 <= b(4) and w2428;
w3168 <= b(5) and w2277;
w3169 <= not w3167 and not w3168;
w3170 <= not w3166 and w3169;
w3171 <= w202 and w2285;
w3172 <= w3170 and not w3171;
w3173 <= a(26) and not w3172;
w3174 <= a(26) and not w3173;
w3175 <= not w3172 and not w3173;
w3176 <= not w3174 and not w3175;
w3177 <= a(29) and not a(30);
w3178 <= not a(29) and a(30);
w3179 <= not w3177 and not w3178;
w3180 <= b(0) and not w3179;
w3181 <= not w2998 and w3180;
w3182 <= w2998 and not w3180;
w3183 <= not w3181 and not w3182;
w3184 <= b(3) and w2793;
w3185 <= b(1) and w2986;
w3186 <= b(2) and w2788;
w3187 <= not w3185 and not w3186;
w3188 <= not w3184 and w3187;
w3189 <= w61 and w2796;
w3190 <= w3188 and not w3189;
w3191 <= a(29) and not w3190;
w3192 <= a(29) and not w3191;
w3193 <= not w3190 and not w3191;
w3194 <= not w3192 and not w3193;
w3195 <= not w3183 and not w3194;
w3196 <= w3183 and w3194;
w3197 <= not w3195 and not w3196;
w3198 <= not w3176 and w3197;
w3199 <= w3197 and not w3198;
w3200 <= not w3176 and not w3198;
w3201 <= not w3199 and not w3200;
w3202 <= not w3016 and w3201;
w3203 <= w3016 and not w3201;
w3204 <= not w3202 and not w3203;
w3205 <= b(9) and w1791;
w3206 <= b(7) and w1941;
w3207 <= b(8) and w1786;
w3208 <= not w3206 and not w3207;
w3209 <= not w3205 and w3208;
w3210 <= w394 and w1794;
w3211 <= w3209 and not w3210;
w3212 <= a(23) and not w3211;
w3213 <= a(23) and not w3212;
w3214 <= not w3211 and not w3212;
w3215 <= not w3213 and not w3214;
w3216 <= not w3204 and not w3215;
w3217 <= w3204 and w3215;
w3218 <= not w3216 and not w3217;
w3219 <= not w3165 and w3218;
w3220 <= w3165 and not w3218;
w3221 <= not w3219 and not w3220;
w3222 <= w3164 and not w3221;
w3223 <= not w3164 and w3221;
w3224 <= not w3222 and not w3223;
w3225 <= not w3153 and w3224;
w3226 <= w3153 and not w3224;
w3227 <= not w3225 and not w3226;
w3228 <= not w3152 and w3227;
w3229 <= w3227 and not w3228;
w3230 <= not w3152 and not w3228;
w3231 <= not w3229 and not w3230;
w3232 <= not w3042 and not w3048;
w3233 <= w3231 and w3232;
w3234 <= not w3231 and not w3232;
w3235 <= not w3233 and not w3234;
w3236 <= b(18) and w694;
w3237 <= b(16) and w799;
w3238 <= b(17) and w689;
w3239 <= not w3237 and not w3238;
w3240 <= not w3236 and w3239;
w3241 <= w697 and w1309;
w3242 <= w3240 and not w3241;
w3243 <= a(14) and not w3242;
w3244 <= a(14) and not w3243;
w3245 <= not w3242 and not w3243;
w3246 <= not w3244 and not w3245;
w3247 <= w3235 and not w3246;
w3248 <= w3235 and not w3247;
w3249 <= not w3246 and not w3247;
w3250 <= not w3248 and not w3249;
w3251 <= not w3061 and not w3067;
w3252 <= w3250 and w3251;
w3253 <= not w3250 and not w3251;
w3254 <= not w3252 and not w3253;
w3255 <= b(21) and w443;
w3256 <= b(19) and w510;
w3257 <= b(20) and w438;
w3258 <= not w3256 and not w3257;
w3259 <= not w3255 and w3258;
w3260 <= w446 and w1727;
w3261 <= w3259 and not w3260;
w3262 <= a(11) and not w3261;
w3263 <= a(11) and not w3262;
w3264 <= not w3261 and not w3262;
w3265 <= not w3263 and not w3264;
w3266 <= w3254 and not w3265;
w3267 <= w3254 and not w3266;
w3268 <= not w3265 and not w3266;
w3269 <= not w3267 and not w3268;
w3270 <= not w3085 and w3269;
w3271 <= w3085 and not w3269;
w3272 <= not w3270 and not w3271;
w3273 <= b(24) and w254;
w3274 <= b(22) and w284;
w3275 <= b(23) and w249;
w3276 <= not w3274 and not w3275;
w3277 <= not w3273 and w3276;
w3278 <= w257 and w2201;
w3279 <= w3277 and not w3278;
w3280 <= a(8) and not w3279;
w3281 <= a(8) and not w3280;
w3282 <= not w3279 and not w3280;
w3283 <= not w3281 and not w3282;
w3284 <= not w3272 and not w3283;
w3285 <= w3272 and w3283;
w3286 <= not w3284 and not w3285;
w3287 <= w3141 and not w3286;
w3288 <= not w3141 and w3286;
w3289 <= not w3287 and not w3288;
w3290 <= b(27) and w105;
w3291 <= b(25) and w146;
w3292 <= b(26) and w100;
w3293 <= not w3291 and not w3292;
w3294 <= not w3290 and w3293;
w3295 <= w108 and w2733;
w3296 <= w3294 and not w3295;
w3297 <= a(5) and not w3296;
w3298 <= a(5) and not w3297;
w3299 <= not w3296 and not w3297;
w3300 <= not w3298 and not w3299;
w3301 <= w3289 and not w3300;
w3302 <= w3289 and not w3301;
w3303 <= not w3300 and not w3301;
w3304 <= not w3302 and not w3303;
w3305 <= not w3107 and not w3111;
w3306 <= w3304 and w3305;
w3307 <= not w3304 and not w3305;
w3308 <= not w3306 and not w3307;
w3309 <= b(30) and w9;
w3310 <= b(28) and w27;
w3311 <= b(29) and w4;
w3312 <= not w3310 and not w3311;
w3313 <= not w3309 and w3312;
w3314 <= not w3122 and not w3124;
w3315 <= not b(29) and not b(30);
w3316 <= b(29) and b(30);
w3317 <= not w3315 and not w3316;
w3318 <= not w3314 and w3317;
w3319 <= w3314 and not w3317;
w3320 <= not w3318 and not w3319;
w3321 <= w12 and w3320;
w3322 <= w3313 and not w3321;
w3323 <= a(2) and not w3322;
w3324 <= a(2) and not w3323;
w3325 <= not w3322 and not w3323;
w3326 <= not w3324 and not w3325;
w3327 <= w3308 and not w3326;
w3328 <= w3308 and not w3327;
w3329 <= not w3326 and not w3327;
w3330 <= not w3328 and not w3329;
w3331 <= not w3133 and not w3138;
w3332 <= not w3330 and not w3331;
w3333 <= w3330 and w3331;
w3334 <= not w3332 and not w3333;
w3335 <= b(16) and w1045;
w3336 <= b(14) and w1134;
w3337 <= b(15) and w1040;
w3338 <= not w3336 and not w3337;
w3339 <= not w3335 and w3338;
w3340 <= w980 and w1048;
w3341 <= w3339 and not w3340;
w3342 <= a(17) and not w3341;
w3343 <= a(17) and not w3342;
w3344 <= not w3341 and not w3342;
w3345 <= not w3343 and not w3344;
w3346 <= not w3016 and not w3201;
w3347 <= not w3198 and not w3346;
w3348 <= b(7) and w2282;
w3349 <= b(5) and w2428;
w3350 <= b(6) and w2277;
w3351 <= not w3349 and not w3350;
w3352 <= not w3348 and w3351;
w3353 <= w227 and w2285;
w3354 <= w3352 and not w3353;
w3355 <= a(26) and not w3354;
w3356 <= a(26) and not w3355;
w3357 <= not w3354 and not w3355;
w3358 <= not w3356 and not w3357;
w3359 <= w2998 and w3180;
w3360 <= not w3195 and not w3359;
w3361 <= b(4) and w2793;
w3362 <= b(2) and w2986;
w3363 <= b(3) and w2788;
w3364 <= not w3362 and not w3363;
w3365 <= not w3361 and w3364;
w3366 <= w89 and w2796;
w3367 <= w3365 and not w3366;
w3368 <= a(29) and not w3367;
w3369 <= a(29) and not w3368;
w3370 <= not w3367 and not w3368;
w3371 <= not w3369 and not w3370;
w3372 <= a(32) and not w3180;
w3373 <= not a(30) and a(31);
w3374 <= a(30) and not a(31);
w3375 <= not w3373 and not w3374;
w3376 <= w3179 and not w3375;
w3377 <= b(0) and w3376;
w3378 <= not a(31) and a(32);
w3379 <= a(31) and not a(32);
w3380 <= not w3378 and not w3379;
w3381 <= not w3179 and w3380;
w3382 <= b(1) and w3381;
w3383 <= not w3377 and not w3382;
w3384 <= not w3179 and not w3380;
w3385 <= not w15 and w3384;
w3386 <= w3383 and not w3385;
w3387 <= a(32) and not w3386;
w3388 <= a(32) and not w3387;
w3389 <= not w3386 and not w3387;
w3390 <= not w3388 and not w3389;
w3391 <= w3372 and not w3390;
w3392 <= not w3372 and w3390;
w3393 <= not w3391 and not w3392;
w3394 <= w3371 and w3393;
w3395 <= not w3371 and not w3393;
w3396 <= not w3394 and not w3395;
w3397 <= not w3360 and not w3396;
w3398 <= w3360 and w3396;
w3399 <= not w3397 and not w3398;
w3400 <= not w3358 and w3399;
w3401 <= w3358 and not w3399;
w3402 <= not w3400 and not w3401;
w3403 <= not w3347 and w3402;
w3404 <= w3347 and not w3402;
w3405 <= not w3403 and not w3404;
w3406 <= b(10) and w1791;
w3407 <= b(8) and w1941;
w3408 <= b(9) and w1786;
w3409 <= not w3407 and not w3408;
w3410 <= not w3406 and w3409;
w3411 <= w481 and w1794;
w3412 <= w3410 and not w3411;
w3413 <= a(23) and not w3412;
w3414 <= a(23) and not w3413;
w3415 <= not w3412 and not w3413;
w3416 <= not w3414 and not w3415;
w3417 <= w3405 and not w3416;
w3418 <= w3405 and not w3417;
w3419 <= not w3416 and not w3417;
w3420 <= not w3418 and not w3419;
w3421 <= not w3216 and not w3219;
w3422 <= w3420 and w3421;
w3423 <= not w3420 and not w3421;
w3424 <= not w3422 and not w3423;
w3425 <= b(13) and w1370;
w3426 <= b(11) and w1506;
w3427 <= b(12) and w1365;
w3428 <= not w3426 and not w3427;
w3429 <= not w3425 and w3428;
w3430 <= w751 and w1373;
w3431 <= w3429 and not w3430;
w3432 <= a(20) and not w3431;
w3433 <= a(20) and not w3432;
w3434 <= not w3431 and not w3432;
w3435 <= not w3433 and not w3434;
w3436 <= not w3424 and w3435;
w3437 <= w3424 and not w3435;
w3438 <= not w3436 and not w3437;
w3439 <= not w3223 and not w3225;
w3440 <= w3438 and not w3439;
w3441 <= not w3438 and w3439;
w3442 <= not w3440 and not w3441;
w3443 <= not w3345 and w3442;
w3444 <= w3442 and not w3443;
w3445 <= not w3345 and not w3443;
w3446 <= not w3444 and not w3445;
w3447 <= not w3228 and not w3234;
w3448 <= w3446 and w3447;
w3449 <= not w3446 and not w3447;
w3450 <= not w3448 and not w3449;
w3451 <= b(19) and w694;
w3452 <= b(17) and w799;
w3453 <= b(18) and w689;
w3454 <= not w3452 and not w3453;
w3455 <= not w3451 and w3454;
w3456 <= w697 and w1451;
w3457 <= w3455 and not w3456;
w3458 <= a(14) and not w3457;
w3459 <= a(14) and not w3458;
w3460 <= not w3457 and not w3458;
w3461 <= not w3459 and not w3460;
w3462 <= w3450 and not w3461;
w3463 <= w3450 and not w3462;
w3464 <= not w3461 and not w3462;
w3465 <= not w3463 and not w3464;
w3466 <= not w3247 and not w3253;
w3467 <= w3465 and w3466;
w3468 <= not w3465 and not w3466;
w3469 <= not w3467 and not w3468;
w3470 <= b(22) and w443;
w3471 <= b(20) and w510;
w3472 <= b(21) and w438;
w3473 <= not w3471 and not w3472;
w3474 <= not w3470 and w3473;
w3475 <= w446 and w1888;
w3476 <= w3474 and not w3475;
w3477 <= a(11) and not w3476;
w3478 <= a(11) and not w3477;
w3479 <= not w3476 and not w3477;
w3480 <= not w3478 and not w3479;
w3481 <= w3469 and not w3480;
w3482 <= w3469 and not w3481;
w3483 <= not w3480 and not w3481;
w3484 <= not w3482 and not w3483;
w3485 <= not w3085 and not w3269;
w3486 <= not w3266 and not w3485;
w3487 <= w3484 and w3486;
w3488 <= not w3484 and not w3486;
w3489 <= not w3487 and not w3488;
w3490 <= b(25) and w254;
w3491 <= b(23) and w284;
w3492 <= b(24) and w249;
w3493 <= not w3491 and not w3492;
w3494 <= not w3490 and w3493;
w3495 <= w257 and w2228;
w3496 <= w3494 and not w3495;
w3497 <= a(8) and not w3496;
w3498 <= a(8) and not w3497;
w3499 <= not w3496 and not w3497;
w3500 <= not w3498 and not w3499;
w3501 <= w3489 and not w3500;
w3502 <= w3489 and not w3501;
w3503 <= not w3500 and not w3501;
w3504 <= not w3502 and not w3503;
w3505 <= not w3284 and not w3288;
w3506 <= w3504 and w3505;
w3507 <= not w3504 and not w3505;
w3508 <= not w3506 and not w3507;
w3509 <= b(28) and w105;
w3510 <= b(26) and w146;
w3511 <= b(27) and w100;
w3512 <= not w3510 and not w3511;
w3513 <= not w3509 and w3512;
w3514 <= w108 and w2932;
w3515 <= w3513 and not w3514;
w3516 <= a(5) and not w3515;
w3517 <= a(5) and not w3516;
w3518 <= not w3515 and not w3516;
w3519 <= not w3517 and not w3518;
w3520 <= w3508 and not w3519;
w3521 <= w3508 and not w3520;
w3522 <= not w3519 and not w3520;
w3523 <= not w3521 and not w3522;
w3524 <= not w3301 and not w3307;
w3525 <= w3523 and w3524;
w3526 <= not w3523 and not w3524;
w3527 <= not w3525 and not w3526;
w3528 <= b(31) and w9;
w3529 <= b(29) and w27;
w3530 <= b(30) and w4;
w3531 <= not w3529 and not w3530;
w3532 <= not w3528 and w3531;
w3533 <= not w3316 and not w3318;
w3534 <= not b(30) and not b(31);
w3535 <= b(30) and b(31);
w3536 <= not w3534 and not w3535;
w3537 <= not w3533 and w3536;
w3538 <= w3533 and not w3536;
w3539 <= not w3537 and not w3538;
w3540 <= w12 and w3539;
w3541 <= w3532 and not w3540;
w3542 <= a(2) and not w3541;
w3543 <= a(2) and not w3542;
w3544 <= not w3541 and not w3542;
w3545 <= not w3543 and not w3544;
w3546 <= w3527 and not w3545;
w3547 <= w3527 and not w3546;
w3548 <= not w3545 and not w3546;
w3549 <= not w3547 and not w3548;
w3550 <= not w3327 and not w3332;
w3551 <= not w3549 and not w3550;
w3552 <= w3549 and w3550;
w3553 <= not w3551 and not w3552;
w3554 <= not w3546 and not w3551;
w3555 <= not w3520 and not w3526;
w3556 <= b(26) and w254;
w3557 <= b(24) and w284;
w3558 <= b(25) and w249;
w3559 <= not w3557 and not w3558;
w3560 <= not w3556 and w3559;
w3561 <= w257 and w2556;
w3562 <= w3560 and not w3561;
w3563 <= a(8) and not w3562;
w3564 <= a(8) and not w3563;
w3565 <= not w3562 and not w3563;
w3566 <= not w3564 and not w3565;
w3567 <= not w3481 and not w3488;
w3568 <= not w3462 and not w3468;
w3569 <= b(17) and w1045;
w3570 <= b(15) and w1134;
w3571 <= b(16) and w1040;
w3572 <= not w3570 and not w3571;
w3573 <= not w3569 and w3572;
w3574 <= w1048 and w1099;
w3575 <= w3573 and not w3574;
w3576 <= a(17) and not w3575;
w3577 <= a(17) and not w3576;
w3578 <= not w3575 and not w3576;
w3579 <= not w3577 and not w3578;
w3580 <= not w3437 and not w3440;
w3581 <= not w3417 and not w3423;
w3582 <= not w3371 and w3393;
w3583 <= not w3397 and not w3582;
w3584 <= b(2) and w3381;
w3585 <= w3179 and not w3380;
w3586 <= w3375 and w3585;
w3587 <= b(0) and w3586;
w3588 <= b(1) and w3376;
w3589 <= not w3587 and not w3588;
w3590 <= not w3584 and w3589;
w3591 <= w39 and w3384;
w3592 <= w3590 and not w3591;
w3593 <= a(32) and not w3592;
w3594 <= a(32) and not w3593;
w3595 <= not w3592 and not w3593;
w3596 <= not w3594 and not w3595;
w3597 <= not w3391 and w3596;
w3598 <= w3391 and not w3596;
w3599 <= not w3597 and not w3598;
w3600 <= b(5) and w2793;
w3601 <= b(3) and w2986;
w3602 <= b(4) and w2788;
w3603 <= not w3601 and not w3602;
w3604 <= not w3600 and w3603;
w3605 <= w137 and w2796;
w3606 <= w3604 and not w3605;
w3607 <= a(29) and not w3606;
w3608 <= a(29) and not w3607;
w3609 <= not w3606 and not w3607;
w3610 <= not w3608 and not w3609;
w3611 <= w3599 and not w3610;
w3612 <= not w3599 and w3610;
w3613 <= not w3583 and not w3612;
w3614 <= not w3611 and w3613;
w3615 <= not w3583 and not w3614;
w3616 <= not w3611 and not w3614;
w3617 <= not w3612 and w3616;
w3618 <= not w3615 and not w3617;
w3619 <= b(8) and w2282;
w3620 <= b(6) and w2428;
w3621 <= b(7) and w2277;
w3622 <= not w3620 and not w3621;
w3623 <= not w3619 and w3622;
w3624 <= w328 and w2285;
w3625 <= w3623 and not w3624;
w3626 <= a(26) and not w3625;
w3627 <= a(26) and not w3626;
w3628 <= not w3625 and not w3626;
w3629 <= not w3627 and not w3628;
w3630 <= not w3618 and not w3629;
w3631 <= not w3618 and not w3630;
w3632 <= not w3629 and not w3630;
w3633 <= not w3631 and not w3632;
w3634 <= not w3400 and not w3403;
w3635 <= w3633 and w3634;
w3636 <= not w3633 and not w3634;
w3637 <= not w3635 and not w3636;
w3638 <= b(11) and w1791;
w3639 <= b(9) and w1941;
w3640 <= b(10) and w1786;
w3641 <= not w3639 and not w3640;
w3642 <= not w3638 and w3641;
w3643 <= w561 and w1794;
w3644 <= w3642 and not w3643;
w3645 <= a(23) and not w3644;
w3646 <= a(23) and not w3645;
w3647 <= not w3644 and not w3645;
w3648 <= not w3646 and not w3647;
w3649 <= w3637 and not w3648;
w3650 <= not w3637 and w3648;
w3651 <= not w3581 and not w3650;
w3652 <= not w3649 and w3651;
w3653 <= not w3581 and not w3652;
w3654 <= not w3649 and not w3652;
w3655 <= not w3650 and w3654;
w3656 <= not w3653 and not w3655;
w3657 <= b(14) and w1370;
w3658 <= b(12) and w1506;
w3659 <= b(13) and w1365;
w3660 <= not w3658 and not w3659;
w3661 <= not w3657 and w3660;
w3662 <= w777 and w1373;
w3663 <= w3661 and not w3662;
w3664 <= a(20) and not w3663;
w3665 <= a(20) and not w3664;
w3666 <= not w3663 and not w3664;
w3667 <= not w3665 and not w3666;
w3668 <= w3656 and w3667;
w3669 <= not w3656 and not w3667;
w3670 <= not w3668 and not w3669;
w3671 <= not w3580 and w3670;
w3672 <= w3580 and not w3670;
w3673 <= not w3671 and not w3672;
w3674 <= not w3579 and w3673;
w3675 <= w3673 and not w3674;
w3676 <= not w3579 and not w3674;
w3677 <= not w3675 and not w3676;
w3678 <= not w3443 and not w3449;
w3679 <= w3677 and w3678;
w3680 <= not w3677 and not w3678;
w3681 <= not w3679 and not w3680;
w3682 <= b(20) and w694;
w3683 <= b(18) and w799;
w3684 <= b(19) and w689;
w3685 <= not w3683 and not w3684;
w3686 <= not w3682 and w3685;
w3687 <= w697 and w1589;
w3688 <= w3686 and not w3687;
w3689 <= a(14) and not w3688;
w3690 <= a(14) and not w3689;
w3691 <= not w3688 and not w3689;
w3692 <= not w3690 and not w3691;
w3693 <= w3681 and not w3692;
w3694 <= not w3681 and w3692;
w3695 <= not w3568 and not w3694;
w3696 <= not w3693 and w3695;
w3697 <= not w3568 and not w3696;
w3698 <= not w3693 and not w3696;
w3699 <= not w3694 and w3698;
w3700 <= not w3697 and not w3699;
w3701 <= b(23) and w443;
w3702 <= b(21) and w510;
w3703 <= b(22) and w438;
w3704 <= not w3702 and not w3703;
w3705 <= not w3701 and w3704;
w3706 <= w446 and w2043;
w3707 <= w3705 and not w3706;
w3708 <= a(11) and not w3707;
w3709 <= a(11) and not w3708;
w3710 <= not w3707 and not w3708;
w3711 <= not w3709 and not w3710;
w3712 <= w3700 and w3711;
w3713 <= not w3700 and not w3711;
w3714 <= not w3712 and not w3713;
w3715 <= not w3567 and w3714;
w3716 <= w3567 and not w3714;
w3717 <= not w3715 and not w3716;
w3718 <= not w3566 and w3717;
w3719 <= w3717 and not w3718;
w3720 <= not w3566 and not w3718;
w3721 <= not w3719 and not w3720;
w3722 <= not w3501 and not w3507;
w3723 <= w3721 and w3722;
w3724 <= not w3721 and not w3722;
w3725 <= not w3723 and not w3724;
w3726 <= b(29) and w105;
w3727 <= b(27) and w146;
w3728 <= b(28) and w100;
w3729 <= not w3727 and not w3728;
w3730 <= not w3726 and w3729;
w3731 <= w108 and w3126;
w3732 <= w3730 and not w3731;
w3733 <= a(5) and not w3732;
w3734 <= a(5) and not w3733;
w3735 <= not w3732 and not w3733;
w3736 <= not w3734 and not w3735;
w3737 <= w3725 and not w3736;
w3738 <= not w3725 and w3736;
w3739 <= not w3555 and not w3738;
w3740 <= not w3737 and w3739;
w3741 <= not w3555 and not w3740;
w3742 <= not w3737 and not w3740;
w3743 <= not w3738 and w3742;
w3744 <= not w3741 and not w3743;
w3745 <= b(32) and w9;
w3746 <= b(30) and w27;
w3747 <= b(31) and w4;
w3748 <= not w3746 and not w3747;
w3749 <= not w3745 and w3748;
w3750 <= not w3535 and not w3537;
w3751 <= not b(31) and not b(32);
w3752 <= b(31) and b(32);
w3753 <= not w3751 and not w3752;
w3754 <= not w3750 and w3753;
w3755 <= w3750 and not w3753;
w3756 <= not w3754 and not w3755;
w3757 <= w12 and w3756;
w3758 <= w3749 and not w3757;
w3759 <= a(2) and not w3758;
w3760 <= a(2) and not w3759;
w3761 <= not w3758 and not w3759;
w3762 <= not w3760 and not w3761;
w3763 <= not w3744 and w3762;
w3764 <= w3744 and not w3762;
w3765 <= not w3763 and not w3764;
w3766 <= not w3554 and not w3765;
w3767 <= w3554 and w3765;
w3768 <= not w3766 and not w3767;
w3769 <= not w3744 and not w3762;
w3770 <= not w3766 and not w3769;
w3771 <= b(27) and w254;
w3772 <= b(25) and w284;
w3773 <= b(26) and w249;
w3774 <= not w3772 and not w3773;
w3775 <= not w3771 and w3774;
w3776 <= w257 and w2733;
w3777 <= w3775 and not w3776;
w3778 <= a(8) and not w3777;
w3779 <= a(8) and not w3778;
w3780 <= not w3777 and not w3778;
w3781 <= not w3779 and not w3780;
w3782 <= not w3713 and not w3715;
w3783 <= not w3674 and not w3680;
w3784 <= not w3669 and not w3671;
w3785 <= b(15) and w1370;
w3786 <= b(13) and w1506;
w3787 <= b(14) and w1365;
w3788 <= not w3786 and not w3787;
w3789 <= not w3785 and w3788;
w3790 <= w874 and w1373;
w3791 <= w3789 and not w3790;
w3792 <= a(20) and not w3791;
w3793 <= a(20) and not w3792;
w3794 <= not w3791 and not w3792;
w3795 <= not w3793 and not w3794;
w3796 <= not w3630 and not w3636;
w3797 <= b(6) and w2793;
w3798 <= b(4) and w2986;
w3799 <= b(5) and w2788;
w3800 <= not w3798 and not w3799;
w3801 <= not w3797 and w3800;
w3802 <= w202 and w2796;
w3803 <= w3801 and not w3802;
w3804 <= a(29) and not w3803;
w3805 <= a(29) and not w3804;
w3806 <= not w3803 and not w3804;
w3807 <= not w3805 and not w3806;
w3808 <= a(32) and not a(33);
w3809 <= not a(32) and a(33);
w3810 <= not w3808 and not w3809;
w3811 <= b(0) and not w3810;
w3812 <= not w3598 and w3811;
w3813 <= w3598 and not w3811;
w3814 <= not w3812 and not w3813;
w3815 <= b(3) and w3381;
w3816 <= b(1) and w3586;
w3817 <= b(2) and w3376;
w3818 <= not w3816 and not w3817;
w3819 <= not w3815 and w3818;
w3820 <= w61 and w3384;
w3821 <= w3819 and not w3820;
w3822 <= a(32) and not w3821;
w3823 <= a(32) and not w3822;
w3824 <= not w3821 and not w3822;
w3825 <= not w3823 and not w3824;
w3826 <= not w3814 and not w3825;
w3827 <= w3814 and w3825;
w3828 <= not w3826 and not w3827;
w3829 <= not w3807 and w3828;
w3830 <= w3828 and not w3829;
w3831 <= not w3807 and not w3829;
w3832 <= not w3830 and not w3831;
w3833 <= not w3616 and w3832;
w3834 <= w3616 and not w3832;
w3835 <= not w3833 and not w3834;
w3836 <= b(9) and w2282;
w3837 <= b(7) and w2428;
w3838 <= b(8) and w2277;
w3839 <= not w3837 and not w3838;
w3840 <= not w3836 and w3839;
w3841 <= w394 and w2285;
w3842 <= w3840 and not w3841;
w3843 <= a(26) and not w3842;
w3844 <= a(26) and not w3843;
w3845 <= not w3842 and not w3843;
w3846 <= not w3844 and not w3845;
w3847 <= not w3835 and not w3846;
w3848 <= w3835 and w3846;
w3849 <= not w3847 and not w3848;
w3850 <= w3796 and not w3849;
w3851 <= not w3796 and w3849;
w3852 <= not w3850 and not w3851;
w3853 <= b(12) and w1791;
w3854 <= b(10) and w1941;
w3855 <= b(11) and w1786;
w3856 <= not w3854 and not w3855;
w3857 <= not w3853 and w3856;
w3858 <= w585 and w1794;
w3859 <= w3857 and not w3858;
w3860 <= a(23) and not w3859;
w3861 <= a(23) and not w3860;
w3862 <= not w3859 and not w3860;
w3863 <= not w3861 and not w3862;
w3864 <= not w3852 and w3863;
w3865 <= w3852 and not w3863;
w3866 <= not w3864 and not w3865;
w3867 <= not w3654 and w3866;
w3868 <= w3654 and not w3866;
w3869 <= not w3867 and not w3868;
w3870 <= not w3795 and w3869;
w3871 <= w3869 and not w3870;
w3872 <= not w3795 and not w3870;
w3873 <= not w3871 and not w3872;
w3874 <= not w3784 and w3873;
w3875 <= w3784 and not w3873;
w3876 <= not w3874 and not w3875;
w3877 <= b(18) and w1045;
w3878 <= b(16) and w1134;
w3879 <= b(17) and w1040;
w3880 <= not w3878 and not w3879;
w3881 <= not w3877 and w3880;
w3882 <= w1048 and w1309;
w3883 <= w3881 and not w3882;
w3884 <= a(17) and not w3883;
w3885 <= a(17) and not w3884;
w3886 <= not w3883 and not w3884;
w3887 <= not w3885 and not w3886;
w3888 <= not w3876 and not w3887;
w3889 <= w3876 and w3887;
w3890 <= not w3888 and not w3889;
w3891 <= w3783 and not w3890;
w3892 <= not w3783 and w3890;
w3893 <= not w3891 and not w3892;
w3894 <= b(21) and w694;
w3895 <= b(19) and w799;
w3896 <= b(20) and w689;
w3897 <= not w3895 and not w3896;
w3898 <= not w3894 and w3897;
w3899 <= w697 and w1727;
w3900 <= w3898 and not w3899;
w3901 <= a(14) and not w3900;
w3902 <= a(14) and not w3901;
w3903 <= not w3900 and not w3901;
w3904 <= not w3902 and not w3903;
w3905 <= w3893 and not w3904;
w3906 <= w3893 and not w3905;
w3907 <= not w3904 and not w3905;
w3908 <= not w3906 and not w3907;
w3909 <= not w3698 and w3908;
w3910 <= w3698 and not w3908;
w3911 <= not w3909 and not w3910;
w3912 <= b(24) and w443;
w3913 <= b(22) and w510;
w3914 <= b(23) and w438;
w3915 <= not w3913 and not w3914;
w3916 <= not w3912 and w3915;
w3917 <= w446 and w2201;
w3918 <= w3916 and not w3917;
w3919 <= a(11) and not w3918;
w3920 <= a(11) and not w3919;
w3921 <= not w3918 and not w3919;
w3922 <= not w3920 and not w3921;
w3923 <= w3911 and w3922;
w3924 <= not w3911 and not w3922;
w3925 <= not w3923 and not w3924;
w3926 <= not w3782 and w3925;
w3927 <= w3782 and not w3925;
w3928 <= not w3926 and not w3927;
w3929 <= not w3781 and w3928;
w3930 <= w3928 and not w3929;
w3931 <= not w3781 and not w3929;
w3932 <= not w3930 and not w3931;
w3933 <= not w3718 and not w3724;
w3934 <= w3932 and w3933;
w3935 <= not w3932 and not w3933;
w3936 <= not w3934 and not w3935;
w3937 <= b(30) and w105;
w3938 <= b(28) and w146;
w3939 <= b(29) and w100;
w3940 <= not w3938 and not w3939;
w3941 <= not w3937 and w3940;
w3942 <= w108 and w3320;
w3943 <= w3941 and not w3942;
w3944 <= a(5) and not w3943;
w3945 <= a(5) and not w3944;
w3946 <= not w3943 and not w3944;
w3947 <= not w3945 and not w3946;
w3948 <= w3936 and not w3947;
w3949 <= w3936 and not w3948;
w3950 <= not w3947 and not w3948;
w3951 <= not w3949 and not w3950;
w3952 <= not w3742 and w3951;
w3953 <= w3742 and not w3951;
w3954 <= not w3952 and not w3953;
w3955 <= b(33) and w9;
w3956 <= b(31) and w27;
w3957 <= b(32) and w4;
w3958 <= not w3956 and not w3957;
w3959 <= not w3955 and w3958;
w3960 <= not w3752 and not w3754;
w3961 <= not b(32) and not b(33);
w3962 <= b(32) and b(33);
w3963 <= not w3961 and not w3962;
w3964 <= not w3960 and w3963;
w3965 <= w3960 and not w3963;
w3966 <= not w3964 and not w3965;
w3967 <= w12 and w3966;
w3968 <= w3959 and not w3967;
w3969 <= a(2) and not w3968;
w3970 <= a(2) and not w3969;
w3971 <= not w3968 and not w3969;
w3972 <= not w3970 and not w3971;
w3973 <= not w3954 and not w3972;
w3974 <= w3954 and w3972;
w3975 <= not w3973 and not w3974;
w3976 <= not w3770 and w3975;
w3977 <= w3770 and not w3975;
w3978 <= not w3976 and not w3977;
w3979 <= not w3973 and not w3976;
w3980 <= not w3742 and not w3951;
w3981 <= not w3948 and not w3980;
w3982 <= not w3924 and not w3926;
w3983 <= not w3865 and not w3867;
w3984 <= b(10) and w2282;
w3985 <= b(8) and w2428;
w3986 <= b(9) and w2277;
w3987 <= not w3985 and not w3986;
w3988 <= not w3984 and w3987;
w3989 <= w481 and w2285;
w3990 <= w3988 and not w3989;
w3991 <= a(26) and not w3990;
w3992 <= a(26) and not w3991;
w3993 <= not w3990 and not w3991;
w3994 <= not w3992 and not w3993;
w3995 <= not w3616 and not w3832;
w3996 <= not w3829 and not w3995;
w3997 <= b(7) and w2793;
w3998 <= b(5) and w2986;
w3999 <= b(6) and w2788;
w4000 <= not w3998 and not w3999;
w4001 <= not w3997 and w4000;
w4002 <= w227 and w2796;
w4003 <= w4001 and not w4002;
w4004 <= a(29) and not w4003;
w4005 <= a(29) and not w4004;
w4006 <= not w4003 and not w4004;
w4007 <= not w4005 and not w4006;
w4008 <= w3598 and w3811;
w4009 <= not w3826 and not w4008;
w4010 <= b(4) and w3381;
w4011 <= b(2) and w3586;
w4012 <= b(3) and w3376;
w4013 <= not w4011 and not w4012;
w4014 <= not w4010 and w4013;
w4015 <= w89 and w3384;
w4016 <= w4014 and not w4015;
w4017 <= a(32) and not w4016;
w4018 <= a(32) and not w4017;
w4019 <= not w4016 and not w4017;
w4020 <= not w4018 and not w4019;
w4021 <= a(35) and not w3811;
w4022 <= not a(33) and a(34);
w4023 <= a(33) and not a(34);
w4024 <= not w4022 and not w4023;
w4025 <= w3810 and not w4024;
w4026 <= b(0) and w4025;
w4027 <= not a(34) and a(35);
w4028 <= a(34) and not a(35);
w4029 <= not w4027 and not w4028;
w4030 <= not w3810 and w4029;
w4031 <= b(1) and w4030;
w4032 <= not w4026 and not w4031;
w4033 <= not w3810 and not w4029;
w4034 <= not w15 and w4033;
w4035 <= w4032 and not w4034;
w4036 <= a(35) and not w4035;
w4037 <= a(35) and not w4036;
w4038 <= not w4035 and not w4036;
w4039 <= not w4037 and not w4038;
w4040 <= w4021 and not w4039;
w4041 <= not w4021 and w4039;
w4042 <= not w4040 and not w4041;
w4043 <= w4020 and not w4042;
w4044 <= not w4020 and w4042;
w4045 <= not w4043 and not w4044;
w4046 <= not w4009 and w4045;
w4047 <= w4009 and not w4045;
w4048 <= not w4046 and not w4047;
w4049 <= w4007 and not w4048;
w4050 <= not w4007 and w4048;
w4051 <= not w4049 and not w4050;
w4052 <= not w3996 and w4051;
w4053 <= w3996 and not w4051;
w4054 <= not w4052 and not w4053;
w4055 <= not w3994 and w4054;
w4056 <= w4054 and not w4055;
w4057 <= not w3994 and not w4055;
w4058 <= not w4056 and not w4057;
w4059 <= not w3847 and not w3851;
w4060 <= w4058 and w4059;
w4061 <= not w4058 and not w4059;
w4062 <= not w4060 and not w4061;
w4063 <= b(13) and w1791;
w4064 <= b(11) and w1941;
w4065 <= b(12) and w1786;
w4066 <= not w4064 and not w4065;
w4067 <= not w4063 and w4066;
w4068 <= w751 and w1794;
w4069 <= w4067 and not w4068;
w4070 <= a(23) and not w4069;
w4071 <= a(23) and not w4070;
w4072 <= not w4069 and not w4070;
w4073 <= not w4071 and not w4072;
w4074 <= w4062 and not w4073;
w4075 <= not w4062 and w4073;
w4076 <= not w3983 and not w4075;
w4077 <= not w4074 and w4076;
w4078 <= not w3983 and not w4077;
w4079 <= not w4074 and not w4077;
w4080 <= not w4075 and w4079;
w4081 <= not w4078 and not w4080;
w4082 <= b(16) and w1370;
w4083 <= b(14) and w1506;
w4084 <= b(15) and w1365;
w4085 <= not w4083 and not w4084;
w4086 <= not w4082 and w4085;
w4087 <= w980 and w1373;
w4088 <= w4086 and not w4087;
w4089 <= a(20) and not w4088;
w4090 <= a(20) and not w4089;
w4091 <= not w4088 and not w4089;
w4092 <= not w4090 and not w4091;
w4093 <= not w4081 and not w4092;
w4094 <= not w4081 and not w4093;
w4095 <= not w4092 and not w4093;
w4096 <= not w4094 and not w4095;
w4097 <= not w3784 and not w3873;
w4098 <= not w3870 and not w4097;
w4099 <= w4096 and w4098;
w4100 <= not w4096 and not w4098;
w4101 <= not w4099 and not w4100;
w4102 <= b(19) and w1045;
w4103 <= b(17) and w1134;
w4104 <= b(18) and w1040;
w4105 <= not w4103 and not w4104;
w4106 <= not w4102 and w4105;
w4107 <= w1048 and w1451;
w4108 <= w4106 and not w4107;
w4109 <= a(17) and not w4108;
w4110 <= a(17) and not w4109;
w4111 <= not w4108 and not w4109;
w4112 <= not w4110 and not w4111;
w4113 <= w4101 and not w4112;
w4114 <= w4101 and not w4113;
w4115 <= not w4112 and not w4113;
w4116 <= not w4114 and not w4115;
w4117 <= not w3888 and not w3892;
w4118 <= w4116 and w4117;
w4119 <= not w4116 and not w4117;
w4120 <= not w4118 and not w4119;
w4121 <= b(22) and w694;
w4122 <= b(20) and w799;
w4123 <= b(21) and w689;
w4124 <= not w4122 and not w4123;
w4125 <= not w4121 and w4124;
w4126 <= w697 and w1888;
w4127 <= w4125 and not w4126;
w4128 <= a(14) and not w4127;
w4129 <= a(14) and not w4128;
w4130 <= not w4127 and not w4128;
w4131 <= not w4129 and not w4130;
w4132 <= w4120 and not w4131;
w4133 <= w4120 and not w4132;
w4134 <= not w4131 and not w4132;
w4135 <= not w4133 and not w4134;
w4136 <= not w3698 and not w3908;
w4137 <= not w3905 and not w4136;
w4138 <= w4135 and w4137;
w4139 <= not w4135 and not w4137;
w4140 <= not w4138 and not w4139;
w4141 <= b(25) and w443;
w4142 <= b(23) and w510;
w4143 <= b(24) and w438;
w4144 <= not w4142 and not w4143;
w4145 <= not w4141 and w4144;
w4146 <= w446 and w2228;
w4147 <= w4145 and not w4146;
w4148 <= a(11) and not w4147;
w4149 <= a(11) and not w4148;
w4150 <= not w4147 and not w4148;
w4151 <= not w4149 and not w4150;
w4152 <= w4140 and not w4151;
w4153 <= not w4140 and w4151;
w4154 <= not w3982 and not w4153;
w4155 <= not w4152 and w4154;
w4156 <= not w3982 and not w4155;
w4157 <= not w4152 and not w4155;
w4158 <= not w4153 and w4157;
w4159 <= not w4156 and not w4158;
w4160 <= b(28) and w254;
w4161 <= b(26) and w284;
w4162 <= b(27) and w249;
w4163 <= not w4161 and not w4162;
w4164 <= not w4160 and w4163;
w4165 <= w257 and w2932;
w4166 <= w4164 and not w4165;
w4167 <= a(8) and not w4166;
w4168 <= a(8) and not w4167;
w4169 <= not w4166 and not w4167;
w4170 <= not w4168 and not w4169;
w4171 <= not w4159 and not w4170;
w4172 <= not w4159 and not w4171;
w4173 <= not w4170 and not w4171;
w4174 <= not w4172 and not w4173;
w4175 <= not w3929 and not w3935;
w4176 <= w4174 and w4175;
w4177 <= not w4174 and not w4175;
w4178 <= not w4176 and not w4177;
w4179 <= b(31) and w105;
w4180 <= b(29) and w146;
w4181 <= b(30) and w100;
w4182 <= not w4180 and not w4181;
w4183 <= not w4179 and w4182;
w4184 <= w108 and w3539;
w4185 <= w4183 and not w4184;
w4186 <= a(5) and not w4185;
w4187 <= a(5) and not w4186;
w4188 <= not w4185 and not w4186;
w4189 <= not w4187 and not w4188;
w4190 <= w4178 and not w4189;
w4191 <= not w4178 and w4189;
w4192 <= not w3981 and not w4191;
w4193 <= not w4190 and w4192;
w4194 <= not w3981 and not w4193;
w4195 <= not w4190 and not w4193;
w4196 <= not w4191 and w4195;
w4197 <= not w4194 and not w4196;
w4198 <= b(34) and w9;
w4199 <= b(32) and w27;
w4200 <= b(33) and w4;
w4201 <= not w4199 and not w4200;
w4202 <= not w4198 and w4201;
w4203 <= not w3962 and not w3964;
w4204 <= not b(33) and not b(34);
w4205 <= b(33) and b(34);
w4206 <= not w4204 and not w4205;
w4207 <= not w4203 and w4206;
w4208 <= w4203 and not w4206;
w4209 <= not w4207 and not w4208;
w4210 <= w12 and w4209;
w4211 <= w4202 and not w4210;
w4212 <= a(2) and not w4211;
w4213 <= a(2) and not w4212;
w4214 <= not w4211 and not w4212;
w4215 <= not w4213 and not w4214;
w4216 <= not w4197 and w4215;
w4217 <= w4197 and not w4215;
w4218 <= not w4216 and not w4217;
w4219 <= not w3979 and not w4218;
w4220 <= w3979 and w4218;
w4221 <= not w4219 and not w4220;
w4222 <= not w4197 and not w4215;
w4223 <= not w4219 and not w4222;
w4224 <= b(29) and w254;
w4225 <= b(27) and w284;
w4226 <= b(28) and w249;
w4227 <= not w4225 and not w4226;
w4228 <= not w4224 and w4227;
w4229 <= w257 and w3126;
w4230 <= w4228 and not w4229;
w4231 <= a(8) and not w4230;
w4232 <= a(8) and not w4231;
w4233 <= not w4230 and not w4231;
w4234 <= not w4232 and not w4233;
w4235 <= b(26) and w443;
w4236 <= b(24) and w510;
w4237 <= b(25) and w438;
w4238 <= not w4236 and not w4237;
w4239 <= not w4235 and w4238;
w4240 <= w446 and w2556;
w4241 <= w4239 and not w4240;
w4242 <= a(11) and not w4241;
w4243 <= a(11) and not w4242;
w4244 <= not w4241 and not w4242;
w4245 <= not w4243 and not w4244;
w4246 <= not w4132 and not w4139;
w4247 <= not w4113 and not w4119;
w4248 <= b(17) and w1370;
w4249 <= b(15) and w1506;
w4250 <= b(16) and w1365;
w4251 <= not w4249 and not w4250;
w4252 <= not w4248 and w4251;
w4253 <= w1099 and w1373;
w4254 <= w4252 and not w4253;
w4255 <= a(20) and not w4254;
w4256 <= a(20) and not w4255;
w4257 <= not w4254 and not w4255;
w4258 <= not w4256 and not w4257;
w4259 <= not w4055 and not w4061;
w4260 <= b(11) and w2282;
w4261 <= b(9) and w2428;
w4262 <= b(10) and w2277;
w4263 <= not w4261 and not w4262;
w4264 <= not w4260 and w4263;
w4265 <= w561 and w2285;
w4266 <= w4264 and not w4265;
w4267 <= a(26) and not w4266;
w4268 <= a(26) and not w4267;
w4269 <= not w4266 and not w4267;
w4270 <= not w4268 and not w4269;
w4271 <= not w4050 and not w4052;
w4272 <= not w4044 and not w4046;
w4273 <= b(2) and w4030;
w4274 <= w3810 and not w4029;
w4275 <= w4024 and w4274;
w4276 <= b(0) and w4275;
w4277 <= b(1) and w4025;
w4278 <= not w4276 and not w4277;
w4279 <= not w4273 and w4278;
w4280 <= w39 and w4033;
w4281 <= w4279 and not w4280;
w4282 <= a(35) and not w4281;
w4283 <= a(35) and not w4282;
w4284 <= not w4281 and not w4282;
w4285 <= not w4283 and not w4284;
w4286 <= not w4040 and w4285;
w4287 <= w4040 and not w4285;
w4288 <= not w4286 and not w4287;
w4289 <= b(5) and w3381;
w4290 <= b(3) and w3586;
w4291 <= b(4) and w3376;
w4292 <= not w4290 and not w4291;
w4293 <= not w4289 and w4292;
w4294 <= w137 and w3384;
w4295 <= w4293 and not w4294;
w4296 <= a(32) and not w4295;
w4297 <= a(32) and not w4296;
w4298 <= not w4295 and not w4296;
w4299 <= not w4297 and not w4298;
w4300 <= w4288 and not w4299;
w4301 <= not w4288 and w4299;
w4302 <= not w4272 and not w4301;
w4303 <= not w4300 and w4302;
w4304 <= not w4272 and not w4303;
w4305 <= not w4300 and not w4303;
w4306 <= not w4301 and w4305;
w4307 <= not w4304 and not w4306;
w4308 <= b(8) and w2793;
w4309 <= b(6) and w2986;
w4310 <= b(7) and w2788;
w4311 <= not w4309 and not w4310;
w4312 <= not w4308 and w4311;
w4313 <= w328 and w2796;
w4314 <= w4312 and not w4313;
w4315 <= a(29) and not w4314;
w4316 <= a(29) and not w4315;
w4317 <= not w4314 and not w4315;
w4318 <= not w4316 and not w4317;
w4319 <= not w4307 and not w4318;
w4320 <= not w4307 and not w4319;
w4321 <= not w4318 and not w4319;
w4322 <= not w4320 and not w4321;
w4323 <= not w4271 and not w4322;
w4324 <= w4271 and w4322;
w4325 <= not w4323 and not w4324;
w4326 <= not w4270 and w4325;
w4327 <= not w4270 and not w4326;
w4328 <= w4325 and not w4326;
w4329 <= not w4327 and not w4328;
w4330 <= not w4259 and not w4329;
w4331 <= not w4259 and not w4330;
w4332 <= not w4329 and not w4330;
w4333 <= not w4331 and not w4332;
w4334 <= b(14) and w1791;
w4335 <= b(12) and w1941;
w4336 <= b(13) and w1786;
w4337 <= not w4335 and not w4336;
w4338 <= not w4334 and w4337;
w4339 <= w777 and w1794;
w4340 <= w4338 and not w4339;
w4341 <= a(23) and not w4340;
w4342 <= a(23) and not w4341;
w4343 <= not w4340 and not w4341;
w4344 <= not w4342 and not w4343;
w4345 <= w4333 and w4344;
w4346 <= not w4333 and not w4344;
w4347 <= not w4345 and not w4346;
w4348 <= not w4079 and w4347;
w4349 <= w4079 and not w4347;
w4350 <= not w4348 and not w4349;
w4351 <= not w4258 and w4350;
w4352 <= w4350 and not w4351;
w4353 <= not w4258 and not w4351;
w4354 <= not w4352 and not w4353;
w4355 <= not w4093 and not w4100;
w4356 <= w4354 and w4355;
w4357 <= not w4354 and not w4355;
w4358 <= not w4356 and not w4357;
w4359 <= b(20) and w1045;
w4360 <= b(18) and w1134;
w4361 <= b(19) and w1040;
w4362 <= not w4360 and not w4361;
w4363 <= not w4359 and w4362;
w4364 <= w1048 and w1589;
w4365 <= w4363 and not w4364;
w4366 <= a(17) and not w4365;
w4367 <= a(17) and not w4366;
w4368 <= not w4365 and not w4366;
w4369 <= not w4367 and not w4368;
w4370 <= w4358 and not w4369;
w4371 <= not w4358 and w4369;
w4372 <= not w4247 and not w4371;
w4373 <= not w4370 and w4372;
w4374 <= not w4247 and not w4373;
w4375 <= not w4370 and not w4373;
w4376 <= not w4371 and w4375;
w4377 <= not w4374 and not w4376;
w4378 <= b(23) and w694;
w4379 <= b(21) and w799;
w4380 <= b(22) and w689;
w4381 <= not w4379 and not w4380;
w4382 <= not w4378 and w4381;
w4383 <= w697 and w2043;
w4384 <= w4382 and not w4383;
w4385 <= a(14) and not w4384;
w4386 <= a(14) and not w4385;
w4387 <= not w4384 and not w4385;
w4388 <= not w4386 and not w4387;
w4389 <= w4377 and w4388;
w4390 <= not w4377 and not w4388;
w4391 <= not w4389 and not w4390;
w4392 <= not w4246 and w4391;
w4393 <= w4246 and not w4391;
w4394 <= not w4392 and not w4393;
w4395 <= w4245 and not w4394;
w4396 <= not w4245 and w4394;
w4397 <= not w4395 and not w4396;
w4398 <= not w4157 and w4397;
w4399 <= w4157 and not w4397;
w4400 <= not w4398 and not w4399;
w4401 <= not w4234 and w4400;
w4402 <= w4400 and not w4401;
w4403 <= not w4234 and not w4401;
w4404 <= not w4402 and not w4403;
w4405 <= not w4171 and not w4177;
w4406 <= w4404 and w4405;
w4407 <= not w4404 and not w4405;
w4408 <= not w4406 and not w4407;
w4409 <= b(32) and w105;
w4410 <= b(30) and w146;
w4411 <= b(31) and w100;
w4412 <= not w4410 and not w4411;
w4413 <= not w4409 and w4412;
w4414 <= w108 and w3756;
w4415 <= w4413 and not w4414;
w4416 <= a(5) and not w4415;
w4417 <= a(5) and not w4416;
w4418 <= not w4415 and not w4416;
w4419 <= not w4417 and not w4418;
w4420 <= w4408 and not w4419;
w4421 <= not w4408 and w4419;
w4422 <= not w4195 and not w4421;
w4423 <= not w4420 and w4422;
w4424 <= not w4195 and not w4423;
w4425 <= not w4420 and not w4423;
w4426 <= not w4421 and w4425;
w4427 <= not w4424 and not w4426;
w4428 <= b(35) and w9;
w4429 <= b(33) and w27;
w4430 <= b(34) and w4;
w4431 <= not w4429 and not w4430;
w4432 <= not w4428 and w4431;
w4433 <= not w4205 and not w4207;
w4434 <= not b(34) and not b(35);
w4435 <= b(34) and b(35);
w4436 <= not w4434 and not w4435;
w4437 <= not w4433 and w4436;
w4438 <= w4433 and not w4436;
w4439 <= not w4437 and not w4438;
w4440 <= w12 and w4439;
w4441 <= w4432 and not w4440;
w4442 <= a(2) and not w4441;
w4443 <= a(2) and not w4442;
w4444 <= not w4441 and not w4442;
w4445 <= not w4443 and not w4444;
w4446 <= not w4427 and w4445;
w4447 <= w4427 and not w4445;
w4448 <= not w4446 and not w4447;
w4449 <= not w4223 and not w4448;
w4450 <= w4223 and w4448;
w4451 <= not w4449 and not w4450;
w4452 <= b(33) and w105;
w4453 <= b(31) and w146;
w4454 <= b(32) and w100;
w4455 <= not w4453 and not w4454;
w4456 <= not w4452 and w4455;
w4457 <= w108 and w3966;
w4458 <= w4456 and not w4457;
w4459 <= a(5) and not w4458;
w4460 <= a(5) and not w4459;
w4461 <= not w4458 and not w4459;
w4462 <= not w4460 and not w4461;
w4463 <= not w4401 and not w4407;
w4464 <= not w4396 and not w4398;
w4465 <= b(27) and w443;
w4466 <= b(25) and w510;
w4467 <= b(26) and w438;
w4468 <= not w4466 and not w4467;
w4469 <= not w4465 and w4468;
w4470 <= w446 and w2733;
w4471 <= w4469 and not w4470;
w4472 <= a(11) and not w4471;
w4473 <= a(11) and not w4472;
w4474 <= not w4471 and not w4472;
w4475 <= not w4473 and not w4474;
w4476 <= not w4390 and not w4392;
w4477 <= not w4351 and not w4357;
w4478 <= not w4346 and not w4348;
w4479 <= b(15) and w1791;
w4480 <= b(13) and w1941;
w4481 <= b(14) and w1786;
w4482 <= not w4480 and not w4481;
w4483 <= not w4479 and w4482;
w4484 <= w874 and w1794;
w4485 <= w4483 and not w4484;
w4486 <= a(23) and not w4485;
w4487 <= a(23) and not w4486;
w4488 <= not w4485 and not w4486;
w4489 <= not w4487 and not w4488;
w4490 <= not w4319 and not w4323;
w4491 <= b(6) and w3381;
w4492 <= b(4) and w3586;
w4493 <= b(5) and w3376;
w4494 <= not w4492 and not w4493;
w4495 <= not w4491 and w4494;
w4496 <= w202 and w3384;
w4497 <= w4495 and not w4496;
w4498 <= a(32) and not w4497;
w4499 <= a(32) and not w4498;
w4500 <= not w4497 and not w4498;
w4501 <= not w4499 and not w4500;
w4502 <= a(35) and not a(36);
w4503 <= not a(35) and a(36);
w4504 <= not w4502 and not w4503;
w4505 <= b(0) and not w4504;
w4506 <= not w4287 and w4505;
w4507 <= w4287 and not w4505;
w4508 <= not w4506 and not w4507;
w4509 <= b(3) and w4030;
w4510 <= b(1) and w4275;
w4511 <= b(2) and w4025;
w4512 <= not w4510 and not w4511;
w4513 <= not w4509 and w4512;
w4514 <= w61 and w4033;
w4515 <= w4513 and not w4514;
w4516 <= a(35) and not w4515;
w4517 <= a(35) and not w4516;
w4518 <= not w4515 and not w4516;
w4519 <= not w4517 and not w4518;
w4520 <= not w4508 and not w4519;
w4521 <= w4508 and w4519;
w4522 <= not w4520 and not w4521;
w4523 <= not w4501 and w4522;
w4524 <= w4522 and not w4523;
w4525 <= not w4501 and not w4523;
w4526 <= not w4524 and not w4525;
w4527 <= not w4305 and w4526;
w4528 <= w4305 and not w4526;
w4529 <= not w4527 and not w4528;
w4530 <= b(9) and w2793;
w4531 <= b(7) and w2986;
w4532 <= b(8) and w2788;
w4533 <= not w4531 and not w4532;
w4534 <= not w4530 and w4533;
w4535 <= w394 and w2796;
w4536 <= w4534 and not w4535;
w4537 <= a(29) and not w4536;
w4538 <= a(29) and not w4537;
w4539 <= not w4536 and not w4537;
w4540 <= not w4538 and not w4539;
w4541 <= not w4529 and not w4540;
w4542 <= w4529 and w4540;
w4543 <= not w4541 and not w4542;
w4544 <= w4490 and not w4543;
w4545 <= not w4490 and w4543;
w4546 <= not w4544 and not w4545;
w4547 <= b(12) and w2282;
w4548 <= b(10) and w2428;
w4549 <= b(11) and w2277;
w4550 <= not w4548 and not w4549;
w4551 <= not w4547 and w4550;
w4552 <= w585 and w2285;
w4553 <= w4551 and not w4552;
w4554 <= a(26) and not w4553;
w4555 <= a(26) and not w4554;
w4556 <= not w4553 and not w4554;
w4557 <= not w4555 and not w4556;
w4558 <= not w4546 and w4557;
w4559 <= w4546 and not w4557;
w4560 <= not w4558 and not w4559;
w4561 <= not w4326 and not w4330;
w4562 <= w4560 and not w4561;
w4563 <= not w4560 and w4561;
w4564 <= not w4562 and not w4563;
w4565 <= not w4489 and w4564;
w4566 <= w4564 and not w4565;
w4567 <= not w4489 and not w4565;
w4568 <= not w4566 and not w4567;
w4569 <= not w4478 and w4568;
w4570 <= w4478 and not w4568;
w4571 <= not w4569 and not w4570;
w4572 <= b(18) and w1370;
w4573 <= b(16) and w1506;
w4574 <= b(17) and w1365;
w4575 <= not w4573 and not w4574;
w4576 <= not w4572 and w4575;
w4577 <= w1309 and w1373;
w4578 <= w4576 and not w4577;
w4579 <= a(20) and not w4578;
w4580 <= a(20) and not w4579;
w4581 <= not w4578 and not w4579;
w4582 <= not w4580 and not w4581;
w4583 <= not w4571 and not w4582;
w4584 <= w4571 and w4582;
w4585 <= not w4583 and not w4584;
w4586 <= w4477 and not w4585;
w4587 <= not w4477 and w4585;
w4588 <= not w4586 and not w4587;
w4589 <= b(21) and w1045;
w4590 <= b(19) and w1134;
w4591 <= b(20) and w1040;
w4592 <= not w4590 and not w4591;
w4593 <= not w4589 and w4592;
w4594 <= w1048 and w1727;
w4595 <= w4593 and not w4594;
w4596 <= a(17) and not w4595;
w4597 <= a(17) and not w4596;
w4598 <= not w4595 and not w4596;
w4599 <= not w4597 and not w4598;
w4600 <= w4588 and not w4599;
w4601 <= w4588 and not w4600;
w4602 <= not w4599 and not w4600;
w4603 <= not w4601 and not w4602;
w4604 <= not w4375 and w4603;
w4605 <= w4375 and not w4603;
w4606 <= not w4604 and not w4605;
w4607 <= b(24) and w694;
w4608 <= b(22) and w799;
w4609 <= b(23) and w689;
w4610 <= not w4608 and not w4609;
w4611 <= not w4607 and w4610;
w4612 <= w697 and w2201;
w4613 <= w4611 and not w4612;
w4614 <= a(14) and not w4613;
w4615 <= a(14) and not w4614;
w4616 <= not w4613 and not w4614;
w4617 <= not w4615 and not w4616;
w4618 <= w4606 and w4617;
w4619 <= not w4606 and not w4617;
w4620 <= not w4618 and not w4619;
w4621 <= not w4476 and w4620;
w4622 <= w4476 and not w4620;
w4623 <= not w4621 and not w4622;
w4624 <= not w4475 and w4623;
w4625 <= w4623 and not w4624;
w4626 <= not w4475 and not w4624;
w4627 <= not w4625 and not w4626;
w4628 <= not w4464 and w4627;
w4629 <= w4464 and not w4627;
w4630 <= not w4628 and not w4629;
w4631 <= b(30) and w254;
w4632 <= b(28) and w284;
w4633 <= b(29) and w249;
w4634 <= not w4632 and not w4633;
w4635 <= not w4631 and w4634;
w4636 <= w257 and w3320;
w4637 <= w4635 and not w4636;
w4638 <= a(8) and not w4637;
w4639 <= a(8) and not w4638;
w4640 <= not w4637 and not w4638;
w4641 <= not w4639 and not w4640;
w4642 <= w4630 and w4641;
w4643 <= not w4630 and not w4641;
w4644 <= not w4642 and not w4643;
w4645 <= not w4463 and w4644;
w4646 <= w4463 and not w4644;
w4647 <= not w4645 and not w4646;
w4648 <= not w4462 and w4647;
w4649 <= w4462 and not w4647;
w4650 <= not w4648 and not w4649;
w4651 <= not w4425 and w4650;
w4652 <= w4425 and not w4650;
w4653 <= not w4651 and not w4652;
w4654 <= b(36) and w9;
w4655 <= b(34) and w27;
w4656 <= b(35) and w4;
w4657 <= not w4655 and not w4656;
w4658 <= not w4654 and w4657;
w4659 <= not w4435 and not w4437;
w4660 <= not b(35) and not b(36);
w4661 <= b(35) and b(36);
w4662 <= not w4660 and not w4661;
w4663 <= not w4659 and w4662;
w4664 <= w4659 and not w4662;
w4665 <= not w4663 and not w4664;
w4666 <= w12 and w4665;
w4667 <= w4658 and not w4666;
w4668 <= a(2) and not w4667;
w4669 <= a(2) and not w4668;
w4670 <= not w4667 and not w4668;
w4671 <= not w4669 and not w4670;
w4672 <= w4653 and not w4671;
w4673 <= w4653 and not w4672;
w4674 <= not w4671 and not w4672;
w4675 <= not w4673 and not w4674;
w4676 <= not w4427 and not w4445;
w4677 <= not w4449 and not w4676;
w4678 <= not w4675 and not w4677;
w4679 <= w4675 and w4677;
w4680 <= not w4678 and not w4679;
w4681 <= not w4672 and not w4678;
w4682 <= b(34) and w105;
w4683 <= b(32) and w146;
w4684 <= b(33) and w100;
w4685 <= not w4683 and not w4684;
w4686 <= not w4682 and w4685;
w4687 <= w108 and w4209;
w4688 <= w4686 and not w4687;
w4689 <= a(5) and not w4688;
w4690 <= a(5) and not w4689;
w4691 <= not w4688 and not w4689;
w4692 <= not w4690 and not w4691;
w4693 <= not w4643 and not w4645;
w4694 <= b(31) and w254;
w4695 <= b(29) and w284;
w4696 <= b(30) and w249;
w4697 <= not w4695 and not w4696;
w4698 <= not w4694 and w4697;
w4699 <= w257 and w3539;
w4700 <= w4698 and not w4699;
w4701 <= a(8) and not w4700;
w4702 <= a(8) and not w4701;
w4703 <= not w4700 and not w4701;
w4704 <= not w4702 and not w4703;
w4705 <= not w4464 and not w4627;
w4706 <= not w4624 and not w4705;
w4707 <= not w4619 and not w4621;
w4708 <= b(16) and w1791;
w4709 <= b(14) and w1941;
w4710 <= b(15) and w1786;
w4711 <= not w4709 and not w4710;
w4712 <= not w4708 and w4711;
w4713 <= w980 and w1794;
w4714 <= w4712 and not w4713;
w4715 <= a(23) and not w4714;
w4716 <= a(23) and not w4715;
w4717 <= not w4714 and not w4715;
w4718 <= not w4716 and not w4717;
w4719 <= not w4559 and not w4562;
w4720 <= b(13) and w2282;
w4721 <= b(11) and w2428;
w4722 <= b(12) and w2277;
w4723 <= not w4721 and not w4722;
w4724 <= not w4720 and w4723;
w4725 <= w751 and w2285;
w4726 <= w4724 and not w4725;
w4727 <= a(26) and not w4726;
w4728 <= a(26) and not w4727;
w4729 <= not w4726 and not w4727;
w4730 <= not w4728 and not w4729;
w4731 <= not w4541 and not w4545;
w4732 <= b(10) and w2793;
w4733 <= b(8) and w2986;
w4734 <= b(9) and w2788;
w4735 <= not w4733 and not w4734;
w4736 <= not w4732 and w4735;
w4737 <= w481 and w2796;
w4738 <= w4736 and not w4737;
w4739 <= a(29) and not w4738;
w4740 <= a(29) and not w4739;
w4741 <= not w4738 and not w4739;
w4742 <= not w4740 and not w4741;
w4743 <= not w4305 and not w4526;
w4744 <= not w4523 and not w4743;
w4745 <= b(7) and w3381;
w4746 <= b(5) and w3586;
w4747 <= b(6) and w3376;
w4748 <= not w4746 and not w4747;
w4749 <= not w4745 and w4748;
w4750 <= w227 and w3384;
w4751 <= w4749 and not w4750;
w4752 <= a(32) and not w4751;
w4753 <= a(32) and not w4752;
w4754 <= not w4751 and not w4752;
w4755 <= not w4753 and not w4754;
w4756 <= w4287 and w4505;
w4757 <= not w4520 and not w4756;
w4758 <= b(4) and w4030;
w4759 <= b(2) and w4275;
w4760 <= b(3) and w4025;
w4761 <= not w4759 and not w4760;
w4762 <= not w4758 and w4761;
w4763 <= w89 and w4033;
w4764 <= w4762 and not w4763;
w4765 <= a(35) and not w4764;
w4766 <= a(35) and not w4765;
w4767 <= not w4764 and not w4765;
w4768 <= not w4766 and not w4767;
w4769 <= a(38) and not w4505;
w4770 <= not a(36) and a(37);
w4771 <= a(36) and not a(37);
w4772 <= not w4770 and not w4771;
w4773 <= w4504 and not w4772;
w4774 <= b(0) and w4773;
w4775 <= not a(37) and a(38);
w4776 <= a(37) and not a(38);
w4777 <= not w4775 and not w4776;
w4778 <= not w4504 and w4777;
w4779 <= b(1) and w4778;
w4780 <= not w4774 and not w4779;
w4781 <= not w4504 and not w4777;
w4782 <= not w15 and w4781;
w4783 <= w4780 and not w4782;
w4784 <= a(38) and not w4783;
w4785 <= a(38) and not w4784;
w4786 <= not w4783 and not w4784;
w4787 <= not w4785 and not w4786;
w4788 <= w4769 and not w4787;
w4789 <= not w4769 and w4787;
w4790 <= not w4788 and not w4789;
w4791 <= w4768 and not w4790;
w4792 <= not w4768 and w4790;
w4793 <= not w4791 and not w4792;
w4794 <= not w4757 and w4793;
w4795 <= w4757 and not w4793;
w4796 <= not w4794 and not w4795;
w4797 <= w4755 and not w4796;
w4798 <= not w4755 and w4796;
w4799 <= not w4797 and not w4798;
w4800 <= not w4744 and w4799;
w4801 <= w4744 and not w4799;
w4802 <= not w4800 and not w4801;
w4803 <= w4742 and not w4802;
w4804 <= not w4742 and w4802;
w4805 <= not w4803 and not w4804;
w4806 <= not w4731 and w4805;
w4807 <= w4731 and not w4805;
w4808 <= not w4806 and not w4807;
w4809 <= w4730 and not w4808;
w4810 <= not w4730 and w4808;
w4811 <= not w4809 and not w4810;
w4812 <= not w4719 and w4811;
w4813 <= w4719 and not w4811;
w4814 <= not w4812 and not w4813;
w4815 <= not w4718 and w4814;
w4816 <= w4814 and not w4815;
w4817 <= not w4718 and not w4815;
w4818 <= not w4816 and not w4817;
w4819 <= not w4478 and not w4568;
w4820 <= not w4565 and not w4819;
w4821 <= w4818 and w4820;
w4822 <= not w4818 and not w4820;
w4823 <= not w4821 and not w4822;
w4824 <= b(19) and w1370;
w4825 <= b(17) and w1506;
w4826 <= b(18) and w1365;
w4827 <= not w4825 and not w4826;
w4828 <= not w4824 and w4827;
w4829 <= w1373 and w1451;
w4830 <= w4828 and not w4829;
w4831 <= a(20) and not w4830;
w4832 <= a(20) and not w4831;
w4833 <= not w4830 and not w4831;
w4834 <= not w4832 and not w4833;
w4835 <= w4823 and not w4834;
w4836 <= w4823 and not w4835;
w4837 <= not w4834 and not w4835;
w4838 <= not w4836 and not w4837;
w4839 <= not w4583 and not w4587;
w4840 <= w4838 and w4839;
w4841 <= not w4838 and not w4839;
w4842 <= not w4840 and not w4841;
w4843 <= b(22) and w1045;
w4844 <= b(20) and w1134;
w4845 <= b(21) and w1040;
w4846 <= not w4844 and not w4845;
w4847 <= not w4843 and w4846;
w4848 <= w1048 and w1888;
w4849 <= w4847 and not w4848;
w4850 <= a(17) and not w4849;
w4851 <= a(17) and not w4850;
w4852 <= not w4849 and not w4850;
w4853 <= not w4851 and not w4852;
w4854 <= w4842 and not w4853;
w4855 <= w4842 and not w4854;
w4856 <= not w4853 and not w4854;
w4857 <= not w4855 and not w4856;
w4858 <= not w4375 and not w4603;
w4859 <= not w4600 and not w4858;
w4860 <= w4857 and w4859;
w4861 <= not w4857 and not w4859;
w4862 <= not w4860 and not w4861;
w4863 <= b(25) and w694;
w4864 <= b(23) and w799;
w4865 <= b(24) and w689;
w4866 <= not w4864 and not w4865;
w4867 <= not w4863 and w4866;
w4868 <= w697 and w2228;
w4869 <= w4867 and not w4868;
w4870 <= a(14) and not w4869;
w4871 <= a(14) and not w4870;
w4872 <= not w4869 and not w4870;
w4873 <= not w4871 and not w4872;
w4874 <= w4862 and not w4873;
w4875 <= not w4862 and w4873;
w4876 <= not w4707 and not w4875;
w4877 <= not w4874 and w4876;
w4878 <= not w4707 and not w4877;
w4879 <= not w4874 and not w4877;
w4880 <= not w4875 and w4879;
w4881 <= not w4878 and not w4880;
w4882 <= b(28) and w443;
w4883 <= b(26) and w510;
w4884 <= b(27) and w438;
w4885 <= not w4883 and not w4884;
w4886 <= not w4882 and w4885;
w4887 <= w446 and w2932;
w4888 <= w4886 and not w4887;
w4889 <= a(11) and not w4888;
w4890 <= a(11) and not w4889;
w4891 <= not w4888 and not w4889;
w4892 <= not w4890 and not w4891;
w4893 <= w4881 and w4892;
w4894 <= not w4881 and not w4892;
w4895 <= not w4893 and not w4894;
w4896 <= not w4706 and w4895;
w4897 <= w4706 and not w4895;
w4898 <= not w4896 and not w4897;
w4899 <= w4704 and not w4898;
w4900 <= not w4704 and w4898;
w4901 <= not w4899 and not w4900;
w4902 <= not w4693 and w4901;
w4903 <= w4693 and not w4901;
w4904 <= not w4902 and not w4903;
w4905 <= not w4692 and w4904;
w4906 <= w4904 and not w4905;
w4907 <= not w4692 and not w4905;
w4908 <= not w4906 and not w4907;
w4909 <= not w4648 and not w4651;
w4910 <= w4908 and w4909;
w4911 <= not w4908 and not w4909;
w4912 <= not w4910 and not w4911;
w4913 <= b(37) and w9;
w4914 <= b(35) and w27;
w4915 <= b(36) and w4;
w4916 <= not w4914 and not w4915;
w4917 <= not w4913 and w4916;
w4918 <= not w4661 and not w4663;
w4919 <= not b(36) and not b(37);
w4920 <= b(36) and b(37);
w4921 <= not w4919 and not w4920;
w4922 <= not w4918 and w4921;
w4923 <= w4918 and not w4921;
w4924 <= not w4922 and not w4923;
w4925 <= w12 and w4924;
w4926 <= w4917 and not w4925;
w4927 <= a(2) and not w4926;
w4928 <= a(2) and not w4927;
w4929 <= not w4926 and not w4927;
w4930 <= not w4928 and not w4929;
w4931 <= not w4912 and w4930;
w4932 <= w4912 and not w4930;
w4933 <= not w4931 and not w4932;
w4934 <= not w4681 and w4933;
w4935 <= w4681 and not w4933;
w4936 <= not w4934 and not w4935;
w4937 <= b(38) and w9;
w4938 <= b(36) and w27;
w4939 <= b(37) and w4;
w4940 <= not w4938 and not w4939;
w4941 <= not w4937 and w4940;
w4942 <= not w4920 and not w4922;
w4943 <= not b(37) and not b(38);
w4944 <= b(37) and b(38);
w4945 <= not w4943 and not w4944;
w4946 <= not w4942 and w4945;
w4947 <= w4942 and not w4945;
w4948 <= not w4946 and not w4947;
w4949 <= w12 and w4948;
w4950 <= w4941 and not w4949;
w4951 <= a(2) and not w4950;
w4952 <= a(2) and not w4951;
w4953 <= not w4950 and not w4951;
w4954 <= not w4952 and not w4953;
w4955 <= not w4905 and not w4911;
w4956 <= b(35) and w105;
w4957 <= b(33) and w146;
w4958 <= b(34) and w100;
w4959 <= not w4957 and not w4958;
w4960 <= not w4956 and w4959;
w4961 <= w108 and w4439;
w4962 <= w4960 and not w4961;
w4963 <= a(5) and not w4962;
w4964 <= a(5) and not w4963;
w4965 <= not w4962 and not w4963;
w4966 <= not w4964 and not w4965;
w4967 <= not w4900 and not w4902;
w4968 <= b(32) and w254;
w4969 <= b(30) and w284;
w4970 <= b(31) and w249;
w4971 <= not w4969 and not w4970;
w4972 <= not w4968 and w4971;
w4973 <= w257 and w3756;
w4974 <= w4972 and not w4973;
w4975 <= a(8) and not w4974;
w4976 <= a(8) and not w4975;
w4977 <= not w4974 and not w4975;
w4978 <= not w4976 and not w4977;
w4979 <= not w4894 and not w4896;
w4980 <= b(29) and w443;
w4981 <= b(27) and w510;
w4982 <= b(28) and w438;
w4983 <= not w4981 and not w4982;
w4984 <= not w4980 and w4983;
w4985 <= w446 and w3126;
w4986 <= w4984 and not w4985;
w4987 <= a(11) and not w4986;
w4988 <= a(11) and not w4987;
w4989 <= not w4986 and not w4987;
w4990 <= not w4988 and not w4989;
w4991 <= not w4854 and not w4861;
w4992 <= b(17) and w1791;
w4993 <= b(15) and w1941;
w4994 <= b(16) and w1786;
w4995 <= not w4993 and not w4994;
w4996 <= not w4992 and w4995;
w4997 <= w1099 and w1794;
w4998 <= w4996 and not w4997;
w4999 <= a(23) and not w4998;
w5000 <= a(23) and not w4999;
w5001 <= not w4998 and not w4999;
w5002 <= not w5000 and not w5001;
w5003 <= not w4810 and not w4812;
w5004 <= not w4804 and not w4806;
w5005 <= b(11) and w2793;
w5006 <= b(9) and w2986;
w5007 <= b(10) and w2788;
w5008 <= not w5006 and not w5007;
w5009 <= not w5005 and w5008;
w5010 <= w561 and w2796;
w5011 <= w5009 and not w5010;
w5012 <= a(29) and not w5011;
w5013 <= a(29) and not w5012;
w5014 <= not w5011 and not w5012;
w5015 <= not w5013 and not w5014;
w5016 <= not w4798 and not w4800;
w5017 <= not w4792 and not w4794;
w5018 <= b(2) and w4778;
w5019 <= w4504 and not w4777;
w5020 <= w4772 and w5019;
w5021 <= b(0) and w5020;
w5022 <= b(1) and w4773;
w5023 <= not w5021 and not w5022;
w5024 <= not w5018 and w5023;
w5025 <= w39 and w4781;
w5026 <= w5024 and not w5025;
w5027 <= a(38) and not w5026;
w5028 <= a(38) and not w5027;
w5029 <= not w5026 and not w5027;
w5030 <= not w5028 and not w5029;
w5031 <= not w4788 and w5030;
w5032 <= w4788 and not w5030;
w5033 <= not w5031 and not w5032;
w5034 <= b(5) and w4030;
w5035 <= b(3) and w4275;
w5036 <= b(4) and w4025;
w5037 <= not w5035 and not w5036;
w5038 <= not w5034 and w5037;
w5039 <= w137 and w4033;
w5040 <= w5038 and not w5039;
w5041 <= a(35) and not w5040;
w5042 <= a(35) and not w5041;
w5043 <= not w5040 and not w5041;
w5044 <= not w5042 and not w5043;
w5045 <= w5033 and not w5044;
w5046 <= w5033 and not w5045;
w5047 <= not w5044 and not w5045;
w5048 <= not w5046 and not w5047;
w5049 <= not w5017 and w5048;
w5050 <= w5017 and not w5048;
w5051 <= not w5049 and not w5050;
w5052 <= b(8) and w3381;
w5053 <= b(6) and w3586;
w5054 <= b(7) and w3376;
w5055 <= not w5053 and not w5054;
w5056 <= not w5052 and w5055;
w5057 <= w328 and w3384;
w5058 <= w5056 and not w5057;
w5059 <= a(32) and not w5058;
w5060 <= a(32) and not w5059;
w5061 <= not w5058 and not w5059;
w5062 <= not w5060 and not w5061;
w5063 <= not w5051 and not w5062;
w5064 <= w5051 and w5062;
w5065 <= not w5063 and not w5064;
w5066 <= not w5016 and w5065;
w5067 <= w5016 and not w5065;
w5068 <= not w5066 and not w5067;
w5069 <= not w5015 and w5068;
w5070 <= not w5015 and not w5069;
w5071 <= w5068 and not w5069;
w5072 <= not w5070 and not w5071;
w5073 <= not w5004 and not w5072;
w5074 <= not w5004 and not w5073;
w5075 <= not w5072 and not w5073;
w5076 <= not w5074 and not w5075;
w5077 <= b(14) and w2282;
w5078 <= b(12) and w2428;
w5079 <= b(13) and w2277;
w5080 <= not w5078 and not w5079;
w5081 <= not w5077 and w5080;
w5082 <= w777 and w2285;
w5083 <= w5081 and not w5082;
w5084 <= a(26) and not w5083;
w5085 <= a(26) and not w5084;
w5086 <= not w5083 and not w5084;
w5087 <= not w5085 and not w5086;
w5088 <= w5076 and w5087;
w5089 <= not w5076 and not w5087;
w5090 <= not w5088 and not w5089;
w5091 <= not w5003 and w5090;
w5092 <= w5003 and not w5090;
w5093 <= not w5091 and not w5092;
w5094 <= not w5002 and w5093;
w5095 <= w5093 and not w5094;
w5096 <= not w5002 and not w5094;
w5097 <= not w5095 and not w5096;
w5098 <= not w4815 and not w4822;
w5099 <= w5097 and w5098;
w5100 <= not w5097 and not w5098;
w5101 <= not w5099 and not w5100;
w5102 <= b(20) and w1370;
w5103 <= b(18) and w1506;
w5104 <= b(19) and w1365;
w5105 <= not w5103 and not w5104;
w5106 <= not w5102 and w5105;
w5107 <= w1373 and w1589;
w5108 <= w5106 and not w5107;
w5109 <= a(20) and not w5108;
w5110 <= a(20) and not w5109;
w5111 <= not w5108 and not w5109;
w5112 <= not w5110 and not w5111;
w5113 <= w5101 and not w5112;
w5114 <= w5101 and not w5113;
w5115 <= not w5112 and not w5113;
w5116 <= not w5114 and not w5115;
w5117 <= not w4835 and not w4841;
w5118 <= w5116 and w5117;
w5119 <= not w5116 and not w5117;
w5120 <= not w5118 and not w5119;
w5121 <= b(23) and w1045;
w5122 <= b(21) and w1134;
w5123 <= b(22) and w1040;
w5124 <= not w5122 and not w5123;
w5125 <= not w5121 and w5124;
w5126 <= w1048 and w2043;
w5127 <= w5125 and not w5126;
w5128 <= a(17) and not w5127;
w5129 <= a(17) and not w5128;
w5130 <= not w5127 and not w5128;
w5131 <= not w5129 and not w5130;
w5132 <= w5120 and not w5131;
w5133 <= not w5120 and w5131;
w5134 <= not w4991 and not w5133;
w5135 <= not w5132 and w5134;
w5136 <= not w4991 and not w5135;
w5137 <= not w5132 and not w5135;
w5138 <= not w5133 and w5137;
w5139 <= not w5136 and not w5138;
w5140 <= b(26) and w694;
w5141 <= b(24) and w799;
w5142 <= b(25) and w689;
w5143 <= not w5141 and not w5142;
w5144 <= not w5140 and w5143;
w5145 <= w697 and w2556;
w5146 <= w5144 and not w5145;
w5147 <= a(14) and not w5146;
w5148 <= a(14) and not w5147;
w5149 <= not w5146 and not w5147;
w5150 <= not w5148 and not w5149;
w5151 <= w5139 and w5150;
w5152 <= not w5139 and not w5150;
w5153 <= not w5151 and not w5152;
w5154 <= not w4879 and w5153;
w5155 <= w4879 and not w5153;
w5156 <= not w5154 and not w5155;
w5157 <= w4990 and not w5156;
w5158 <= not w4990 and w5156;
w5159 <= not w5157 and not w5158;
w5160 <= not w4979 and w5159;
w5161 <= w4979 and not w5159;
w5162 <= not w5160 and not w5161;
w5163 <= w4978 and not w5162;
w5164 <= not w4978 and w5162;
w5165 <= not w5163 and not w5164;
w5166 <= not w4967 and w5165;
w5167 <= w4967 and not w5165;
w5168 <= not w5166 and not w5167;
w5169 <= w4966 and not w5168;
w5170 <= not w4966 and w5168;
w5171 <= not w5169 and not w5170;
w5172 <= not w4955 and w5171;
w5173 <= w4955 and not w5171;
w5174 <= not w5172 and not w5173;
w5175 <= not w4954 and w5174;
w5176 <= w5174 and not w5175;
w5177 <= not w4954 and not w5175;
w5178 <= not w5176 and not w5177;
w5179 <= not w4932 and not w4934;
w5180 <= not w5178 and not w5179;
w5181 <= w5178 and w5179;
w5182 <= not w5180 and not w5181;
w5183 <= b(39) and w9;
w5184 <= b(37) and w27;
w5185 <= b(38) and w4;
w5186 <= not w5184 and not w5185;
w5187 <= not w5183 and w5186;
w5188 <= not w4944 and not w4946;
w5189 <= not b(38) and not b(39);
w5190 <= b(38) and b(39);
w5191 <= not w5189 and not w5190;
w5192 <= not w5188 and w5191;
w5193 <= w5188 and not w5191;
w5194 <= not w5192 and not w5193;
w5195 <= w12 and w5194;
w5196 <= w5187 and not w5195;
w5197 <= a(2) and not w5196;
w5198 <= a(2) and not w5197;
w5199 <= not w5196 and not w5197;
w5200 <= not w5198 and not w5199;
w5201 <= not w5170 and not w5172;
w5202 <= not w5164 and not w5166;
w5203 <= b(33) and w254;
w5204 <= b(31) and w284;
w5205 <= b(32) and w249;
w5206 <= not w5204 and not w5205;
w5207 <= not w5203 and w5206;
w5208 <= w257 and w3966;
w5209 <= w5207 and not w5208;
w5210 <= a(8) and not w5209;
w5211 <= a(8) and not w5210;
w5212 <= not w5209 and not w5210;
w5213 <= not w5211 and not w5212;
w5214 <= not w5158 and not w5160;
w5215 <= not w5152 and not w5154;
w5216 <= b(27) and w694;
w5217 <= b(25) and w799;
w5218 <= b(26) and w689;
w5219 <= not w5217 and not w5218;
w5220 <= not w5216 and w5219;
w5221 <= w697 and w2733;
w5222 <= w5220 and not w5221;
w5223 <= a(14) and not w5222;
w5224 <= a(14) and not w5223;
w5225 <= not w5222 and not w5223;
w5226 <= not w5224 and not w5225;
w5227 <= not w5094 and not w5100;
w5228 <= not w5089 and not w5091;
w5229 <= b(15) and w2282;
w5230 <= b(13) and w2428;
w5231 <= b(14) and w2277;
w5232 <= not w5230 and not w5231;
w5233 <= not w5229 and w5232;
w5234 <= w874 and w2285;
w5235 <= w5233 and not w5234;
w5236 <= a(26) and not w5235;
w5237 <= a(26) and not w5236;
w5238 <= not w5235 and not w5236;
w5239 <= not w5237 and not w5238;
w5240 <= b(6) and w4030;
w5241 <= b(4) and w4275;
w5242 <= b(5) and w4025;
w5243 <= not w5241 and not w5242;
w5244 <= not w5240 and w5243;
w5245 <= w202 and w4033;
w5246 <= w5244 and not w5245;
w5247 <= a(35) and not w5246;
w5248 <= a(35) and not w5247;
w5249 <= not w5246 and not w5247;
w5250 <= not w5248 and not w5249;
w5251 <= a(38) and not a(39);
w5252 <= not a(38) and a(39);
w5253 <= not w5251 and not w5252;
w5254 <= b(0) and not w5253;
w5255 <= not w5032 and w5254;
w5256 <= w5032 and not w5254;
w5257 <= not w5255 and not w5256;
w5258 <= b(3) and w4778;
w5259 <= b(1) and w5020;
w5260 <= b(2) and w4773;
w5261 <= not w5259 and not w5260;
w5262 <= not w5258 and w5261;
w5263 <= w61 and w4781;
w5264 <= w5262 and not w5263;
w5265 <= a(38) and not w5264;
w5266 <= a(38) and not w5265;
w5267 <= not w5264 and not w5265;
w5268 <= not w5266 and not w5267;
w5269 <= not w5257 and not w5268;
w5270 <= w5257 and w5268;
w5271 <= not w5269 and not w5270;
w5272 <= not w5250 and w5271;
w5273 <= w5271 and not w5272;
w5274 <= not w5250 and not w5272;
w5275 <= not w5273 and not w5274;
w5276 <= not w5017 and not w5048;
w5277 <= not w5045 and not w5276;
w5278 <= w5275 and w5277;
w5279 <= not w5275 and not w5277;
w5280 <= not w5278 and not w5279;
w5281 <= b(9) and w3381;
w5282 <= b(7) and w3586;
w5283 <= b(8) and w3376;
w5284 <= not w5282 and not w5283;
w5285 <= not w5281 and w5284;
w5286 <= w394 and w3384;
w5287 <= w5285 and not w5286;
w5288 <= a(32) and not w5287;
w5289 <= a(32) and not w5288;
w5290 <= not w5287 and not w5288;
w5291 <= not w5289 and not w5290;
w5292 <= w5280 and not w5291;
w5293 <= w5280 and not w5292;
w5294 <= not w5291 and not w5292;
w5295 <= not w5293 and not w5294;
w5296 <= not w5063 and not w5066;
w5297 <= w5295 and w5296;
w5298 <= not w5295 and not w5296;
w5299 <= not w5297 and not w5298;
w5300 <= b(12) and w2793;
w5301 <= b(10) and w2986;
w5302 <= b(11) and w2788;
w5303 <= not w5301 and not w5302;
w5304 <= not w5300 and w5303;
w5305 <= w585 and w2796;
w5306 <= w5304 and not w5305;
w5307 <= a(29) and not w5306;
w5308 <= a(29) and not w5307;
w5309 <= not w5306 and not w5307;
w5310 <= not w5308 and not w5309;
w5311 <= not w5299 and w5310;
w5312 <= w5299 and not w5310;
w5313 <= not w5311 and not w5312;
w5314 <= not w5069 and not w5073;
w5315 <= w5313 and not w5314;
w5316 <= not w5313 and w5314;
w5317 <= not w5315 and not w5316;
w5318 <= not w5239 and w5317;
w5319 <= w5317 and not w5318;
w5320 <= not w5239 and not w5318;
w5321 <= not w5319 and not w5320;
w5322 <= not w5228 and w5321;
w5323 <= w5228 and not w5321;
w5324 <= not w5322 and not w5323;
w5325 <= b(18) and w1791;
w5326 <= b(16) and w1941;
w5327 <= b(17) and w1786;
w5328 <= not w5326 and not w5327;
w5329 <= not w5325 and w5328;
w5330 <= w1309 and w1794;
w5331 <= w5329 and not w5330;
w5332 <= a(23) and not w5331;
w5333 <= a(23) and not w5332;
w5334 <= not w5331 and not w5332;
w5335 <= not w5333 and not w5334;
w5336 <= not w5324 and not w5335;
w5337 <= w5324 and w5335;
w5338 <= not w5336 and not w5337;
w5339 <= w5227 and not w5338;
w5340 <= not w5227 and w5338;
w5341 <= not w5339 and not w5340;
w5342 <= b(21) and w1370;
w5343 <= b(19) and w1506;
w5344 <= b(20) and w1365;
w5345 <= not w5343 and not w5344;
w5346 <= not w5342 and w5345;
w5347 <= w1373 and w1727;
w5348 <= w5346 and not w5347;
w5349 <= a(20) and not w5348;
w5350 <= a(20) and not w5349;
w5351 <= not w5348 and not w5349;
w5352 <= not w5350 and not w5351;
w5353 <= w5341 and not w5352;
w5354 <= w5341 and not w5353;
w5355 <= not w5352 and not w5353;
w5356 <= not w5354 and not w5355;
w5357 <= not w5113 and not w5119;
w5358 <= w5356 and w5357;
w5359 <= not w5356 and not w5357;
w5360 <= not w5358 and not w5359;
w5361 <= b(24) and w1045;
w5362 <= b(22) and w1134;
w5363 <= b(23) and w1040;
w5364 <= not w5362 and not w5363;
w5365 <= not w5361 and w5364;
w5366 <= w1048 and w2201;
w5367 <= w5365 and not w5366;
w5368 <= a(17) and not w5367;
w5369 <= a(17) and not w5368;
w5370 <= not w5367 and not w5368;
w5371 <= not w5369 and not w5370;
w5372 <= not w5360 and w5371;
w5373 <= w5360 and not w5371;
w5374 <= not w5372 and not w5373;
w5375 <= not w5137 and w5374;
w5376 <= w5137 and not w5374;
w5377 <= not w5375 and not w5376;
w5378 <= not w5226 and w5377;
w5379 <= w5377 and not w5378;
w5380 <= not w5226 and not w5378;
w5381 <= not w5379 and not w5380;
w5382 <= not w5215 and w5381;
w5383 <= w5215 and not w5381;
w5384 <= not w5382 and not w5383;
w5385 <= b(30) and w443;
w5386 <= b(28) and w510;
w5387 <= b(29) and w438;
w5388 <= not w5386 and not w5387;
w5389 <= not w5385 and w5388;
w5390 <= w446 and w3320;
w5391 <= w5389 and not w5390;
w5392 <= a(11) and not w5391;
w5393 <= a(11) and not w5392;
w5394 <= not w5391 and not w5392;
w5395 <= not w5393 and not w5394;
w5396 <= not w5384 and not w5395;
w5397 <= w5384 and w5395;
w5398 <= not w5396 and not w5397;
w5399 <= not w5214 and w5398;
w5400 <= w5214 and not w5398;
w5401 <= not w5399 and not w5400;
w5402 <= not w5213 and w5401;
w5403 <= w5401 and not w5402;
w5404 <= not w5213 and not w5402;
w5405 <= not w5403 and not w5404;
w5406 <= not w5202 and w5405;
w5407 <= w5202 and not w5405;
w5408 <= not w5406 and not w5407;
w5409 <= b(36) and w105;
w5410 <= b(34) and w146;
w5411 <= b(35) and w100;
w5412 <= not w5410 and not w5411;
w5413 <= not w5409 and w5412;
w5414 <= w108 and w4665;
w5415 <= w5413 and not w5414;
w5416 <= a(5) and not w5415;
w5417 <= a(5) and not w5416;
w5418 <= not w5415 and not w5416;
w5419 <= not w5417 and not w5418;
w5420 <= w5408 and w5419;
w5421 <= not w5408 and not w5419;
w5422 <= not w5420 and not w5421;
w5423 <= not w5201 and w5422;
w5424 <= w5201 and not w5422;
w5425 <= not w5423 and not w5424;
w5426 <= not w5200 and w5425;
w5427 <= w5425 and not w5426;
w5428 <= not w5200 and not w5426;
w5429 <= not w5427 and not w5428;
w5430 <= not w5175 and not w5180;
w5431 <= not w5429 and not w5430;
w5432 <= w5429 and w5430;
w5433 <= not w5431 and not w5432;
w5434 <= not w5426 and not w5431;
w5435 <= not w5421 and not w5423;
w5436 <= b(37) and w105;
w5437 <= b(35) and w146;
w5438 <= b(36) and w100;
w5439 <= not w5437 and not w5438;
w5440 <= not w5436 and w5439;
w5441 <= w108 and w4924;
w5442 <= w5440 and not w5441;
w5443 <= a(5) and not w5442;
w5444 <= a(5) and not w5443;
w5445 <= not w5442 and not w5443;
w5446 <= not w5444 and not w5445;
w5447 <= not w5202 and not w5405;
w5448 <= not w5402 and not w5447;
w5449 <= b(34) and w254;
w5450 <= b(32) and w284;
w5451 <= b(33) and w249;
w5452 <= not w5450 and not w5451;
w5453 <= not w5449 and w5452;
w5454 <= w257 and w4209;
w5455 <= w5453 and not w5454;
w5456 <= a(8) and not w5455;
w5457 <= a(8) and not w5456;
w5458 <= not w5455 and not w5456;
w5459 <= not w5457 and not w5458;
w5460 <= not w5396 and not w5399;
w5461 <= not w5215 and not w5381;
w5462 <= not w5378 and not w5461;
w5463 <= b(28) and w694;
w5464 <= b(26) and w799;
w5465 <= b(27) and w689;
w5466 <= not w5464 and not w5465;
w5467 <= not w5463 and w5466;
w5468 <= w697 and w2932;
w5469 <= w5467 and not w5468;
w5470 <= a(14) and not w5469;
w5471 <= a(14) and not w5470;
w5472 <= not w5469 and not w5470;
w5473 <= not w5471 and not w5472;
w5474 <= b(16) and w2282;
w5475 <= b(14) and w2428;
w5476 <= b(15) and w2277;
w5477 <= not w5475 and not w5476;
w5478 <= not w5474 and w5477;
w5479 <= w980 and w2285;
w5480 <= w5478 and not w5479;
w5481 <= a(26) and not w5480;
w5482 <= a(26) and not w5481;
w5483 <= not w5480 and not w5481;
w5484 <= not w5482 and not w5483;
w5485 <= not w5312 and not w5315;
w5486 <= not w5292 and not w5298;
w5487 <= b(7) and w4030;
w5488 <= b(5) and w4275;
w5489 <= b(6) and w4025;
w5490 <= not w5488 and not w5489;
w5491 <= not w5487 and w5490;
w5492 <= w227 and w4033;
w5493 <= w5491 and not w5492;
w5494 <= a(35) and not w5493;
w5495 <= a(35) and not w5494;
w5496 <= not w5493 and not w5494;
w5497 <= not w5495 and not w5496;
w5498 <= w5032 and w5254;
w5499 <= not w5269 and not w5498;
w5500 <= b(4) and w4778;
w5501 <= b(2) and w5020;
w5502 <= b(3) and w4773;
w5503 <= not w5501 and not w5502;
w5504 <= not w5500 and w5503;
w5505 <= w89 and w4781;
w5506 <= w5504 and not w5505;
w5507 <= a(38) and not w5506;
w5508 <= a(38) and not w5507;
w5509 <= not w5506 and not w5507;
w5510 <= not w5508 and not w5509;
w5511 <= a(41) and not w5254;
w5512 <= not a(39) and a(40);
w5513 <= a(39) and not a(40);
w5514 <= not w5512 and not w5513;
w5515 <= w5253 and not w5514;
w5516 <= b(0) and w5515;
w5517 <= not a(40) and a(41);
w5518 <= a(40) and not a(41);
w5519 <= not w5517 and not w5518;
w5520 <= not w5253 and w5519;
w5521 <= b(1) and w5520;
w5522 <= not w5516 and not w5521;
w5523 <= not w5253 and not w5519;
w5524 <= not w15 and w5523;
w5525 <= w5522 and not w5524;
w5526 <= a(41) and not w5525;
w5527 <= a(41) and not w5526;
w5528 <= not w5525 and not w5526;
w5529 <= not w5527 and not w5528;
w5530 <= w5511 and not w5529;
w5531 <= not w5511 and w5529;
w5532 <= not w5530 and not w5531;
w5533 <= w5510 and not w5532;
w5534 <= not w5510 and w5532;
w5535 <= not w5533 and not w5534;
w5536 <= not w5499 and w5535;
w5537 <= w5499 and not w5535;
w5538 <= not w5536 and not w5537;
w5539 <= not w5497 and w5538;
w5540 <= w5538 and not w5539;
w5541 <= not w5497 and not w5539;
w5542 <= not w5540 and not w5541;
w5543 <= not w5272 and not w5279;
w5544 <= w5542 and w5543;
w5545 <= not w5542 and not w5543;
w5546 <= not w5544 and not w5545;
w5547 <= b(10) and w3381;
w5548 <= b(8) and w3586;
w5549 <= b(9) and w3376;
w5550 <= not w5548 and not w5549;
w5551 <= not w5547 and w5550;
w5552 <= w481 and w3384;
w5553 <= w5551 and not w5552;
w5554 <= a(32) and not w5553;
w5555 <= a(32) and not w5554;
w5556 <= not w5553 and not w5554;
w5557 <= not w5555 and not w5556;
w5558 <= w5546 and not w5557;
w5559 <= not w5546 and w5557;
w5560 <= not w5486 and not w5559;
w5561 <= not w5558 and w5560;
w5562 <= not w5486 and not w5561;
w5563 <= not w5558 and not w5561;
w5564 <= not w5559 and w5563;
w5565 <= not w5562 and not w5564;
w5566 <= b(13) and w2793;
w5567 <= b(11) and w2986;
w5568 <= b(12) and w2788;
w5569 <= not w5567 and not w5568;
w5570 <= not w5566 and w5569;
w5571 <= w751 and w2796;
w5572 <= w5570 and not w5571;
w5573 <= a(29) and not w5572;
w5574 <= a(29) and not w5573;
w5575 <= not w5572 and not w5573;
w5576 <= not w5574 and not w5575;
w5577 <= w5565 and w5576;
w5578 <= not w5565 and not w5576;
w5579 <= not w5577 and not w5578;
w5580 <= not w5485 and w5579;
w5581 <= w5485 and not w5579;
w5582 <= not w5580 and not w5581;
w5583 <= not w5484 and w5582;
w5584 <= w5582 and not w5583;
w5585 <= not w5484 and not w5583;
w5586 <= not w5584 and not w5585;
w5587 <= not w5228 and not w5321;
w5588 <= not w5318 and not w5587;
w5589 <= w5586 and w5588;
w5590 <= not w5586 and not w5588;
w5591 <= not w5589 and not w5590;
w5592 <= b(19) and w1791;
w5593 <= b(17) and w1941;
w5594 <= b(18) and w1786;
w5595 <= not w5593 and not w5594;
w5596 <= not w5592 and w5595;
w5597 <= w1451 and w1794;
w5598 <= w5596 and not w5597;
w5599 <= a(23) and not w5598;
w5600 <= a(23) and not w5599;
w5601 <= not w5598 and not w5599;
w5602 <= not w5600 and not w5601;
w5603 <= w5591 and not w5602;
w5604 <= w5591 and not w5603;
w5605 <= not w5602 and not w5603;
w5606 <= not w5604 and not w5605;
w5607 <= not w5336 and not w5340;
w5608 <= w5606 and w5607;
w5609 <= not w5606 and not w5607;
w5610 <= not w5608 and not w5609;
w5611 <= b(22) and w1370;
w5612 <= b(20) and w1506;
w5613 <= b(21) and w1365;
w5614 <= not w5612 and not w5613;
w5615 <= not w5611 and w5614;
w5616 <= w1373 and w1888;
w5617 <= w5615 and not w5616;
w5618 <= a(20) and not w5617;
w5619 <= a(20) and not w5618;
w5620 <= not w5617 and not w5618;
w5621 <= not w5619 and not w5620;
w5622 <= w5610 and not w5621;
w5623 <= w5610 and not w5622;
w5624 <= not w5621 and not w5622;
w5625 <= not w5623 and not w5624;
w5626 <= not w5353 and not w5359;
w5627 <= w5625 and w5626;
w5628 <= not w5625 and not w5626;
w5629 <= not w5627 and not w5628;
w5630 <= b(25) and w1045;
w5631 <= b(23) and w1134;
w5632 <= b(24) and w1040;
w5633 <= not w5631 and not w5632;
w5634 <= not w5630 and w5633;
w5635 <= w1048 and w2228;
w5636 <= w5634 and not w5635;
w5637 <= a(17) and not w5636;
w5638 <= a(17) and not w5637;
w5639 <= not w5636 and not w5637;
w5640 <= not w5638 and not w5639;
w5641 <= w5629 and not w5640;
w5642 <= w5629 and not w5641;
w5643 <= not w5640 and not w5641;
w5644 <= not w5642 and not w5643;
w5645 <= not w5373 and not w5375;
w5646 <= not w5644 and not w5645;
w5647 <= w5644 and w5645;
w5648 <= not w5646 and not w5647;
w5649 <= not w5473 and w5648;
w5650 <= not w5473 and not w5649;
w5651 <= w5648 and not w5649;
w5652 <= not w5650 and not w5651;
w5653 <= not w5462 and not w5652;
w5654 <= not w5462 and not w5653;
w5655 <= not w5652 and not w5653;
w5656 <= not w5654 and not w5655;
w5657 <= b(31) and w443;
w5658 <= b(29) and w510;
w5659 <= b(30) and w438;
w5660 <= not w5658 and not w5659;
w5661 <= not w5657 and w5660;
w5662 <= w446 and w3539;
w5663 <= w5661 and not w5662;
w5664 <= a(11) and not w5663;
w5665 <= a(11) and not w5664;
w5666 <= not w5663 and not w5664;
w5667 <= not w5665 and not w5666;
w5668 <= w5656 and w5667;
w5669 <= not w5656 and not w5667;
w5670 <= not w5668 and not w5669;
w5671 <= not w5460 and w5670;
w5672 <= w5460 and not w5670;
w5673 <= not w5671 and not w5672;
w5674 <= w5459 and not w5673;
w5675 <= not w5459 and w5673;
w5676 <= not w5674 and not w5675;
w5677 <= not w5448 and w5676;
w5678 <= w5448 and not w5676;
w5679 <= not w5677 and not w5678;
w5680 <= not w5446 and w5679;
w5681 <= w5679 and not w5680;
w5682 <= not w5446 and not w5680;
w5683 <= not w5681 and not w5682;
w5684 <= not w5435 and w5683;
w5685 <= w5435 and not w5683;
w5686 <= not w5684 and not w5685;
w5687 <= b(40) and w9;
w5688 <= b(38) and w27;
w5689 <= b(39) and w4;
w5690 <= not w5688 and not w5689;
w5691 <= not w5687 and w5690;
w5692 <= not w5190 and not w5192;
w5693 <= not b(39) and not b(40);
w5694 <= b(39) and b(40);
w5695 <= not w5693 and not w5694;
w5696 <= not w5692 and w5695;
w5697 <= w5692 and not w5695;
w5698 <= not w5696 and not w5697;
w5699 <= w12 and w5698;
w5700 <= w5691 and not w5699;
w5701 <= a(2) and not w5700;
w5702 <= a(2) and not w5701;
w5703 <= not w5700 and not w5701;
w5704 <= not w5702 and not w5703;
w5705 <= not w5686 and not w5704;
w5706 <= w5686 and w5704;
w5707 <= not w5705 and not w5706;
w5708 <= not w5434 and w5707;
w5709 <= w5434 and not w5707;
w5710 <= not w5708 and not w5709;
w5711 <= not w5705 and not w5708;
w5712 <= not w5435 and not w5683;
w5713 <= not w5680 and not w5712;
w5714 <= not w5675 and not w5677;
w5715 <= b(35) and w254;
w5716 <= b(33) and w284;
w5717 <= b(34) and w249;
w5718 <= not w5716 and not w5717;
w5719 <= not w5715 and w5718;
w5720 <= w257 and w4439;
w5721 <= w5719 and not w5720;
w5722 <= a(8) and not w5721;
w5723 <= a(8) and not w5722;
w5724 <= not w5721 and not w5722;
w5725 <= not w5723 and not w5724;
w5726 <= not w5669 and not w5671;
w5727 <= b(32) and w443;
w5728 <= b(30) and w510;
w5729 <= b(31) and w438;
w5730 <= not w5728 and not w5729;
w5731 <= not w5727 and w5730;
w5732 <= w446 and w3756;
w5733 <= w5731 and not w5732;
w5734 <= a(11) and not w5733;
w5735 <= a(11) and not w5734;
w5736 <= not w5733 and not w5734;
w5737 <= not w5735 and not w5736;
w5738 <= not w5649 and not w5653;
w5739 <= b(29) and w694;
w5740 <= b(27) and w799;
w5741 <= b(28) and w689;
w5742 <= not w5740 and not w5741;
w5743 <= not w5739 and w5742;
w5744 <= w697 and w3126;
w5745 <= w5743 and not w5744;
w5746 <= a(14) and not w5745;
w5747 <= a(14) and not w5746;
w5748 <= not w5745 and not w5746;
w5749 <= not w5747 and not w5748;
w5750 <= not w5641 and not w5646;
w5751 <= not w5622 and not w5628;
w5752 <= b(20) and w1791;
w5753 <= b(18) and w1941;
w5754 <= b(19) and w1786;
w5755 <= not w5753 and not w5754;
w5756 <= not w5752 and w5755;
w5757 <= w1589 and w1794;
w5758 <= w5756 and not w5757;
w5759 <= a(23) and not w5758;
w5760 <= a(23) and not w5759;
w5761 <= not w5758 and not w5759;
w5762 <= not w5760 and not w5761;
w5763 <= not w5583 and not w5590;
w5764 <= b(17) and w2282;
w5765 <= b(15) and w2428;
w5766 <= b(16) and w2277;
w5767 <= not w5765 and not w5766;
w5768 <= not w5764 and w5767;
w5769 <= w1099 and w2285;
w5770 <= w5768 and not w5769;
w5771 <= a(26) and not w5770;
w5772 <= a(26) and not w5771;
w5773 <= not w5770 and not w5771;
w5774 <= not w5772 and not w5773;
w5775 <= not w5578 and not w5580;
w5776 <= b(14) and w2793;
w5777 <= b(12) and w2986;
w5778 <= b(13) and w2788;
w5779 <= not w5777 and not w5778;
w5780 <= not w5776 and w5779;
w5781 <= w777 and w2796;
w5782 <= w5780 and not w5781;
w5783 <= a(29) and not w5782;
w5784 <= a(29) and not w5783;
w5785 <= not w5782 and not w5783;
w5786 <= not w5784 and not w5785;
w5787 <= not w5539 and not w5545;
w5788 <= b(8) and w4030;
w5789 <= b(6) and w4275;
w5790 <= b(7) and w4025;
w5791 <= not w5789 and not w5790;
w5792 <= not w5788 and w5791;
w5793 <= w328 and w4033;
w5794 <= w5792 and not w5793;
w5795 <= a(35) and not w5794;
w5796 <= a(35) and not w5795;
w5797 <= not w5794 and not w5795;
w5798 <= not w5796 and not w5797;
w5799 <= not w5534 and not w5536;
w5800 <= b(2) and w5520;
w5801 <= w5253 and not w5519;
w5802 <= w5514 and w5801;
w5803 <= b(0) and w5802;
w5804 <= b(1) and w5515;
w5805 <= not w5803 and not w5804;
w5806 <= not w5800 and w5805;
w5807 <= w39 and w5523;
w5808 <= w5806 and not w5807;
w5809 <= a(41) and not w5808;
w5810 <= a(41) and not w5809;
w5811 <= not w5808 and not w5809;
w5812 <= not w5810 and not w5811;
w5813 <= not w5530 and w5812;
w5814 <= w5530 and not w5812;
w5815 <= not w5813 and not w5814;
w5816 <= b(5) and w4778;
w5817 <= b(3) and w5020;
w5818 <= b(4) and w4773;
w5819 <= not w5817 and not w5818;
w5820 <= not w5816 and w5819;
w5821 <= w137 and w4781;
w5822 <= w5820 and not w5821;
w5823 <= a(38) and not w5822;
w5824 <= a(38) and not w5823;
w5825 <= not w5822 and not w5823;
w5826 <= not w5824 and not w5825;
w5827 <= w5815 and not w5826;
w5828 <= w5815 and not w5827;
w5829 <= not w5826 and not w5827;
w5830 <= not w5828 and not w5829;
w5831 <= not w5799 and not w5830;
w5832 <= w5799 and w5830;
w5833 <= not w5831 and not w5832;
w5834 <= not w5798 and w5833;
w5835 <= not w5798 and not w5834;
w5836 <= w5833 and not w5834;
w5837 <= not w5835 and not w5836;
w5838 <= not w5787 and not w5837;
w5839 <= not w5787 and not w5838;
w5840 <= not w5837 and not w5838;
w5841 <= not w5839 and not w5840;
w5842 <= b(11) and w3381;
w5843 <= b(9) and w3586;
w5844 <= b(10) and w3376;
w5845 <= not w5843 and not w5844;
w5846 <= not w5842 and w5845;
w5847 <= w561 and w3384;
w5848 <= w5846 and not w5847;
w5849 <= a(32) and not w5848;
w5850 <= a(32) and not w5849;
w5851 <= not w5848 and not w5849;
w5852 <= not w5850 and not w5851;
w5853 <= w5841 and w5852;
w5854 <= not w5841 and not w5852;
w5855 <= not w5853 and not w5854;
w5856 <= not w5563 and w5855;
w5857 <= w5563 and not w5855;
w5858 <= not w5856 and not w5857;
w5859 <= w5786 and not w5858;
w5860 <= not w5786 and w5858;
w5861 <= not w5859 and not w5860;
w5862 <= not w5775 and w5861;
w5863 <= w5775 and not w5861;
w5864 <= not w5862 and not w5863;
w5865 <= w5774 and not w5864;
w5866 <= not w5774 and w5864;
w5867 <= not w5865 and not w5866;
w5868 <= not w5763 and w5867;
w5869 <= w5763 and not w5867;
w5870 <= not w5868 and not w5869;
w5871 <= not w5762 and w5870;
w5872 <= w5870 and not w5871;
w5873 <= not w5762 and not w5871;
w5874 <= not w5872 and not w5873;
w5875 <= not w5603 and not w5609;
w5876 <= w5874 and w5875;
w5877 <= not w5874 and not w5875;
w5878 <= not w5876 and not w5877;
w5879 <= b(23) and w1370;
w5880 <= b(21) and w1506;
w5881 <= b(22) and w1365;
w5882 <= not w5880 and not w5881;
w5883 <= not w5879 and w5882;
w5884 <= w1373 and w2043;
w5885 <= w5883 and not w5884;
w5886 <= a(20) and not w5885;
w5887 <= a(20) and not w5886;
w5888 <= not w5885 and not w5886;
w5889 <= not w5887 and not w5888;
w5890 <= w5878 and not w5889;
w5891 <= not w5878 and w5889;
w5892 <= not w5751 and not w5891;
w5893 <= not w5890 and w5892;
w5894 <= not w5751 and not w5893;
w5895 <= not w5890 and not w5893;
w5896 <= not w5891 and w5895;
w5897 <= not w5894 and not w5896;
w5898 <= b(26) and w1045;
w5899 <= b(24) and w1134;
w5900 <= b(25) and w1040;
w5901 <= not w5899 and not w5900;
w5902 <= not w5898 and w5901;
w5903 <= w1048 and w2556;
w5904 <= w5902 and not w5903;
w5905 <= a(17) and not w5904;
w5906 <= a(17) and not w5905;
w5907 <= not w5904 and not w5905;
w5908 <= not w5906 and not w5907;
w5909 <= w5897 and w5908;
w5910 <= not w5897 and not w5908;
w5911 <= not w5909 and not w5910;
w5912 <= not w5750 and w5911;
w5913 <= w5750 and not w5911;
w5914 <= not w5912 and not w5913;
w5915 <= w5749 and not w5914;
w5916 <= not w5749 and w5914;
w5917 <= not w5915 and not w5916;
w5918 <= not w5738 and w5917;
w5919 <= w5738 and not w5917;
w5920 <= not w5918 and not w5919;
w5921 <= w5737 and not w5920;
w5922 <= not w5737 and w5920;
w5923 <= not w5921 and not w5922;
w5924 <= not w5726 and w5923;
w5925 <= w5726 and not w5923;
w5926 <= not w5924 and not w5925;
w5927 <= not w5725 and w5926;
w5928 <= w5926 and not w5927;
w5929 <= not w5725 and not w5927;
w5930 <= not w5928 and not w5929;
w5931 <= not w5714 and w5930;
w5932 <= w5714 and not w5930;
w5933 <= not w5931 and not w5932;
w5934 <= b(38) and w105;
w5935 <= b(36) and w146;
w5936 <= b(37) and w100;
w5937 <= not w5935 and not w5936;
w5938 <= not w5934 and w5937;
w5939 <= w108 and w4948;
w5940 <= w5938 and not w5939;
w5941 <= a(5) and not w5940;
w5942 <= a(5) and not w5941;
w5943 <= not w5940 and not w5941;
w5944 <= not w5942 and not w5943;
w5945 <= not w5933 and not w5944;
w5946 <= w5933 and w5944;
w5947 <= not w5945 and not w5946;
w5948 <= w5713 and not w5947;
w5949 <= not w5713 and w5947;
w5950 <= not w5948 and not w5949;
w5951 <= b(41) and w9;
w5952 <= b(39) and w27;
w5953 <= b(40) and w4;
w5954 <= not w5952 and not w5953;
w5955 <= not w5951 and w5954;
w5956 <= not w5694 and not w5696;
w5957 <= not b(40) and not b(41);
w5958 <= b(40) and b(41);
w5959 <= not w5957 and not w5958;
w5960 <= not w5956 and w5959;
w5961 <= w5956 and not w5959;
w5962 <= not w5960 and not w5961;
w5963 <= w12 and w5962;
w5964 <= w5955 and not w5963;
w5965 <= a(2) and not w5964;
w5966 <= a(2) and not w5965;
w5967 <= not w5964 and not w5965;
w5968 <= not w5966 and not w5967;
w5969 <= not w5950 and w5968;
w5970 <= w5950 and not w5968;
w5971 <= not w5969 and not w5970;
w5972 <= not w5711 and w5971;
w5973 <= w5711 and not w5971;
w5974 <= not w5972 and not w5973;
w5975 <= not w5945 and not w5949;
w5976 <= b(39) and w105;
w5977 <= b(37) and w146;
w5978 <= b(38) and w100;
w5979 <= not w5977 and not w5978;
w5980 <= not w5976 and w5979;
w5981 <= w108 and w5194;
w5982 <= w5980 and not w5981;
w5983 <= a(5) and not w5982;
w5984 <= a(5) and not w5983;
w5985 <= not w5982 and not w5983;
w5986 <= not w5984 and not w5985;
w5987 <= not w5714 and not w5930;
w5988 <= not w5927 and not w5987;
w5989 <= not w5922 and not w5924;
w5990 <= b(33) and w443;
w5991 <= b(31) and w510;
w5992 <= b(32) and w438;
w5993 <= not w5991 and not w5992;
w5994 <= not w5990 and w5993;
w5995 <= w446 and w3966;
w5996 <= w5994 and not w5995;
w5997 <= a(11) and not w5996;
w5998 <= a(11) and not w5997;
w5999 <= not w5996 and not w5997;
w6000 <= not w5998 and not w5999;
w6001 <= not w5916 and not w5918;
w6002 <= not w5910 and not w5912;
w6003 <= b(27) and w1045;
w6004 <= b(25) and w1134;
w6005 <= b(26) and w1040;
w6006 <= not w6004 and not w6005;
w6007 <= not w6003 and w6006;
w6008 <= w1048 and w2733;
w6009 <= w6007 and not w6008;
w6010 <= a(17) and not w6009;
w6011 <= a(17) and not w6010;
w6012 <= not w6009 and not w6010;
w6013 <= not w6011 and not w6012;
w6014 <= b(21) and w1791;
w6015 <= b(19) and w1941;
w6016 <= b(20) and w1786;
w6017 <= not w6015 and not w6016;
w6018 <= not w6014 and w6017;
w6019 <= w1727 and w1794;
w6020 <= w6018 and not w6019;
w6021 <= a(23) and not w6020;
w6022 <= a(23) and not w6021;
w6023 <= not w6020 and not w6021;
w6024 <= not w6022 and not w6023;
w6025 <= not w5866 and not w5868;
w6026 <= not w5860 and not w5862;
w6027 <= not w5854 and not w5856;
w6028 <= b(12) and w3381;
w6029 <= b(10) and w3586;
w6030 <= b(11) and w3376;
w6031 <= not w6029 and not w6030;
w6032 <= not w6028 and w6031;
w6033 <= w585 and w3384;
w6034 <= w6032 and not w6033;
w6035 <= a(32) and not w6034;
w6036 <= a(32) and not w6035;
w6037 <= not w6034 and not w6035;
w6038 <= not w6036 and not w6037;
w6039 <= not w5834 and not w5838;
w6040 <= b(6) and w4778;
w6041 <= b(4) and w5020;
w6042 <= b(5) and w4773;
w6043 <= not w6041 and not w6042;
w6044 <= not w6040 and w6043;
w6045 <= w202 and w4781;
w6046 <= w6044 and not w6045;
w6047 <= a(38) and not w6046;
w6048 <= a(38) and not w6047;
w6049 <= not w6046 and not w6047;
w6050 <= not w6048 and not w6049;
w6051 <= a(41) and not a(42);
w6052 <= not a(41) and a(42);
w6053 <= not w6051 and not w6052;
w6054 <= b(0) and not w6053;
w6055 <= not w5814 and w6054;
w6056 <= w5814 and not w6054;
w6057 <= not w6055 and not w6056;
w6058 <= b(3) and w5520;
w6059 <= b(1) and w5802;
w6060 <= b(2) and w5515;
w6061 <= not w6059 and not w6060;
w6062 <= not w6058 and w6061;
w6063 <= w61 and w5523;
w6064 <= w6062 and not w6063;
w6065 <= a(41) and not w6064;
w6066 <= a(41) and not w6065;
w6067 <= not w6064 and not w6065;
w6068 <= not w6066 and not w6067;
w6069 <= not w6057 and not w6068;
w6070 <= w6057 and w6068;
w6071 <= not w6069 and not w6070;
w6072 <= not w6050 and w6071;
w6073 <= w6071 and not w6072;
w6074 <= not w6050 and not w6072;
w6075 <= not w6073 and not w6074;
w6076 <= not w5827 and not w5831;
w6077 <= w6075 and w6076;
w6078 <= not w6075 and not w6076;
w6079 <= not w6077 and not w6078;
w6080 <= b(9) and w4030;
w6081 <= b(7) and w4275;
w6082 <= b(8) and w4025;
w6083 <= not w6081 and not w6082;
w6084 <= not w6080 and w6083;
w6085 <= w394 and w4033;
w6086 <= w6084 and not w6085;
w6087 <= a(35) and not w6086;
w6088 <= a(35) and not w6087;
w6089 <= not w6086 and not w6087;
w6090 <= not w6088 and not w6089;
w6091 <= not w6079 and w6090;
w6092 <= w6079 and not w6090;
w6093 <= not w6091 and not w6092;
w6094 <= not w6039 and w6093;
w6095 <= w6039 and not w6093;
w6096 <= not w6094 and not w6095;
w6097 <= not w6038 and w6096;
w6098 <= not w6038 and not w6097;
w6099 <= w6096 and not w6097;
w6100 <= not w6098 and not w6099;
w6101 <= not w6027 and not w6100;
w6102 <= not w6027 and not w6101;
w6103 <= not w6100 and not w6101;
w6104 <= not w6102 and not w6103;
w6105 <= b(15) and w2793;
w6106 <= b(13) and w2986;
w6107 <= b(14) and w2788;
w6108 <= not w6106 and not w6107;
w6109 <= not w6105 and w6108;
w6110 <= w874 and w2796;
w6111 <= w6109 and not w6110;
w6112 <= a(29) and not w6111;
w6113 <= a(29) and not w6112;
w6114 <= not w6111 and not w6112;
w6115 <= not w6113 and not w6114;
w6116 <= not w6104 and not w6115;
w6117 <= not w6104 and not w6116;
w6118 <= not w6115 and not w6116;
w6119 <= not w6117 and not w6118;
w6120 <= not w6026 and w6119;
w6121 <= w6026 and not w6119;
w6122 <= not w6120 and not w6121;
w6123 <= b(18) and w2282;
w6124 <= b(16) and w2428;
w6125 <= b(17) and w2277;
w6126 <= not w6124 and not w6125;
w6127 <= not w6123 and w6126;
w6128 <= w1309 and w2285;
w6129 <= w6127 and not w6128;
w6130 <= a(26) and not w6129;
w6131 <= a(26) and not w6130;
w6132 <= not w6129 and not w6130;
w6133 <= not w6131 and not w6132;
w6134 <= not w6122 and not w6133;
w6135 <= w6122 and w6133;
w6136 <= not w6134 and not w6135;
w6137 <= not w6025 and w6136;
w6138 <= w6025 and not w6136;
w6139 <= not w6137 and not w6138;
w6140 <= not w6024 and w6139;
w6141 <= w6139 and not w6140;
w6142 <= not w6024 and not w6140;
w6143 <= not w6141 and not w6142;
w6144 <= not w5871 and not w5877;
w6145 <= w6143 and w6144;
w6146 <= not w6143 and not w6144;
w6147 <= not w6145 and not w6146;
w6148 <= b(24) and w1370;
w6149 <= b(22) and w1506;
w6150 <= b(23) and w1365;
w6151 <= not w6149 and not w6150;
w6152 <= not w6148 and w6151;
w6153 <= w1373 and w2201;
w6154 <= w6152 and not w6153;
w6155 <= a(20) and not w6154;
w6156 <= a(20) and not w6155;
w6157 <= not w6154 and not w6155;
w6158 <= not w6156 and not w6157;
w6159 <= not w6147 and w6158;
w6160 <= w6147 and not w6158;
w6161 <= not w6159 and not w6160;
w6162 <= not w5895 and w6161;
w6163 <= w5895 and not w6161;
w6164 <= not w6162 and not w6163;
w6165 <= not w6013 and w6164;
w6166 <= w6164 and not w6165;
w6167 <= not w6013 and not w6165;
w6168 <= not w6166 and not w6167;
w6169 <= not w6002 and w6168;
w6170 <= w6002 and not w6168;
w6171 <= not w6169 and not w6170;
w6172 <= b(30) and w694;
w6173 <= b(28) and w799;
w6174 <= b(29) and w689;
w6175 <= not w6173 and not w6174;
w6176 <= not w6172 and w6175;
w6177 <= w697 and w3320;
w6178 <= w6176 and not w6177;
w6179 <= a(14) and not w6178;
w6180 <= a(14) and not w6179;
w6181 <= not w6178 and not w6179;
w6182 <= not w6180 and not w6181;
w6183 <= not w6171 and not w6182;
w6184 <= w6171 and w6182;
w6185 <= not w6183 and not w6184;
w6186 <= not w6001 and w6185;
w6187 <= w6001 and not w6185;
w6188 <= not w6186 and not w6187;
w6189 <= not w6000 and w6188;
w6190 <= w6188 and not w6189;
w6191 <= not w6000 and not w6189;
w6192 <= not w6190 and not w6191;
w6193 <= not w5989 and w6192;
w6194 <= w5989 and not w6192;
w6195 <= not w6193 and not w6194;
w6196 <= b(36) and w254;
w6197 <= b(34) and w284;
w6198 <= b(35) and w249;
w6199 <= not w6197 and not w6198;
w6200 <= not w6196 and w6199;
w6201 <= w257 and w4665;
w6202 <= w6200 and not w6201;
w6203 <= a(8) and not w6202;
w6204 <= a(8) and not w6203;
w6205 <= not w6202 and not w6203;
w6206 <= not w6204 and not w6205;
w6207 <= w6195 and w6206;
w6208 <= not w6195 and not w6206;
w6209 <= not w6207 and not w6208;
w6210 <= not w5988 and w6209;
w6211 <= w5988 and not w6209;
w6212 <= not w6210 and not w6211;
w6213 <= not w5986 and w6212;
w6214 <= not w5986 and not w6213;
w6215 <= w6212 and not w6213;
w6216 <= not w6214 and not w6215;
w6217 <= not w5975 and not w6216;
w6218 <= not w5975 and not w6217;
w6219 <= not w6216 and not w6217;
w6220 <= not w6218 and not w6219;
w6221 <= b(42) and w9;
w6222 <= b(40) and w27;
w6223 <= b(41) and w4;
w6224 <= not w6222 and not w6223;
w6225 <= not w6221 and w6224;
w6226 <= not w5958 and not w5960;
w6227 <= not b(41) and not b(42);
w6228 <= b(41) and b(42);
w6229 <= not w6227 and not w6228;
w6230 <= not w6226 and w6229;
w6231 <= w6226 and not w6229;
w6232 <= not w6230 and not w6231;
w6233 <= w12 and w6232;
w6234 <= w6225 and not w6233;
w6235 <= a(2) and not w6234;
w6236 <= a(2) and not w6235;
w6237 <= not w6234 and not w6235;
w6238 <= not w6236 and not w6237;
w6239 <= not w6220 and not w6238;
w6240 <= not w6220 and not w6239;
w6241 <= not w6238 and not w6239;
w6242 <= not w6240 and not w6241;
w6243 <= not w5970 and not w5972;
w6244 <= not w6242 and not w6243;
w6245 <= w6242 and w6243;
w6246 <= not w6244 and not w6245;
w6247 <= b(43) and w9;
w6248 <= b(41) and w27;
w6249 <= b(42) and w4;
w6250 <= not w6248 and not w6249;
w6251 <= not w6247 and w6250;
w6252 <= not w6228 and not w6230;
w6253 <= not b(42) and not b(43);
w6254 <= b(42) and b(43);
w6255 <= not w6253 and not w6254;
w6256 <= not w6252 and w6255;
w6257 <= w6252 and not w6255;
w6258 <= not w6256 and not w6257;
w6259 <= w12 and w6258;
w6260 <= w6251 and not w6259;
w6261 <= a(2) and not w6260;
w6262 <= a(2) and not w6261;
w6263 <= not w6260 and not w6261;
w6264 <= not w6262 and not w6263;
w6265 <= not w6213 and not w6217;
w6266 <= not w6208 and not w6210;
w6267 <= b(34) and w443;
w6268 <= b(32) and w510;
w6269 <= b(33) and w438;
w6270 <= not w6268 and not w6269;
w6271 <= not w6267 and w6270;
w6272 <= w446 and w4209;
w6273 <= w6271 and not w6272;
w6274 <= a(11) and not w6273;
w6275 <= a(11) and not w6274;
w6276 <= not w6273 and not w6274;
w6277 <= not w6275 and not w6276;
w6278 <= not w6183 and not w6186;
w6279 <= not w6002 and not w6168;
w6280 <= not w6165 and not w6279;
w6281 <= b(28) and w1045;
w6282 <= b(26) and w1134;
w6283 <= b(27) and w1040;
w6284 <= not w6282 and not w6283;
w6285 <= not w6281 and w6284;
w6286 <= w1048 and w2932;
w6287 <= w6285 and not w6286;
w6288 <= a(17) and not w6287;
w6289 <= a(17) and not w6288;
w6290 <= not w6287 and not w6288;
w6291 <= not w6289 and not w6290;
w6292 <= b(16) and w2793;
w6293 <= b(14) and w2986;
w6294 <= b(15) and w2788;
w6295 <= not w6293 and not w6294;
w6296 <= not w6292 and w6295;
w6297 <= w980 and w2796;
w6298 <= w6296 and not w6297;
w6299 <= a(29) and not w6298;
w6300 <= a(29) and not w6299;
w6301 <= not w6298 and not w6299;
w6302 <= not w6300 and not w6301;
w6303 <= not w6097 and not w6101;
w6304 <= not w6092 and not w6094;
w6305 <= b(7) and w4778;
w6306 <= b(5) and w5020;
w6307 <= b(6) and w4773;
w6308 <= not w6306 and not w6307;
w6309 <= not w6305 and w6308;
w6310 <= w227 and w4781;
w6311 <= w6309 and not w6310;
w6312 <= a(38) and not w6311;
w6313 <= a(38) and not w6312;
w6314 <= not w6311 and not w6312;
w6315 <= not w6313 and not w6314;
w6316 <= w5814 and w6054;
w6317 <= not w6069 and not w6316;
w6318 <= b(4) and w5520;
w6319 <= b(2) and w5802;
w6320 <= b(3) and w5515;
w6321 <= not w6319 and not w6320;
w6322 <= not w6318 and w6321;
w6323 <= w89 and w5523;
w6324 <= w6322 and not w6323;
w6325 <= a(41) and not w6324;
w6326 <= a(41) and not w6325;
w6327 <= not w6324 and not w6325;
w6328 <= not w6326 and not w6327;
w6329 <= a(44) and not w6054;
w6330 <= not a(42) and a(43);
w6331 <= a(42) and not a(43);
w6332 <= not w6330 and not w6331;
w6333 <= w6053 and not w6332;
w6334 <= b(0) and w6333;
w6335 <= not a(43) and a(44);
w6336 <= a(43) and not a(44);
w6337 <= not w6335 and not w6336;
w6338 <= not w6053 and w6337;
w6339 <= b(1) and w6338;
w6340 <= not w6334 and not w6339;
w6341 <= not w6053 and not w6337;
w6342 <= not w15 and w6341;
w6343 <= w6340 and not w6342;
w6344 <= a(44) and not w6343;
w6345 <= a(44) and not w6344;
w6346 <= not w6343 and not w6344;
w6347 <= not w6345 and not w6346;
w6348 <= w6329 and not w6347;
w6349 <= not w6329 and w6347;
w6350 <= not w6348 and not w6349;
w6351 <= w6328 and not w6350;
w6352 <= not w6328 and w6350;
w6353 <= not w6351 and not w6352;
w6354 <= not w6317 and w6353;
w6355 <= w6317 and not w6353;
w6356 <= not w6354 and not w6355;
w6357 <= not w6315 and w6356;
w6358 <= w6356 and not w6357;
w6359 <= not w6315 and not w6357;
w6360 <= not w6358 and not w6359;
w6361 <= not w6072 and not w6078;
w6362 <= w6360 and w6361;
w6363 <= not w6360 and not w6361;
w6364 <= not w6362 and not w6363;
w6365 <= b(10) and w4030;
w6366 <= b(8) and w4275;
w6367 <= b(9) and w4025;
w6368 <= not w6366 and not w6367;
w6369 <= not w6365 and w6368;
w6370 <= w481 and w4033;
w6371 <= w6369 and not w6370;
w6372 <= a(35) and not w6371;
w6373 <= a(35) and not w6372;
w6374 <= not w6371 and not w6372;
w6375 <= not w6373 and not w6374;
w6376 <= w6364 and not w6375;
w6377 <= not w6364 and w6375;
w6378 <= not w6304 and not w6377;
w6379 <= not w6376 and w6378;
w6380 <= not w6304 and not w6379;
w6381 <= not w6376 and not w6379;
w6382 <= not w6377 and w6381;
w6383 <= not w6380 and not w6382;
w6384 <= b(13) and w3381;
w6385 <= b(11) and w3586;
w6386 <= b(12) and w3376;
w6387 <= not w6385 and not w6386;
w6388 <= not w6384 and w6387;
w6389 <= w751 and w3384;
w6390 <= w6388 and not w6389;
w6391 <= a(32) and not w6390;
w6392 <= a(32) and not w6391;
w6393 <= not w6390 and not w6391;
w6394 <= not w6392 and not w6393;
w6395 <= w6383 and w6394;
w6396 <= not w6383 and not w6394;
w6397 <= not w6395 and not w6396;
w6398 <= not w6303 and w6397;
w6399 <= w6303 and not w6397;
w6400 <= not w6398 and not w6399;
w6401 <= not w6302 and w6400;
w6402 <= w6400 and not w6401;
w6403 <= not w6302 and not w6401;
w6404 <= not w6402 and not w6403;
w6405 <= not w6026 and not w6119;
w6406 <= not w6116 and not w6405;
w6407 <= w6404 and w6406;
w6408 <= not w6404 and not w6406;
w6409 <= not w6407 and not w6408;
w6410 <= b(19) and w2282;
w6411 <= b(17) and w2428;
w6412 <= b(18) and w2277;
w6413 <= not w6411 and not w6412;
w6414 <= not w6410 and w6413;
w6415 <= w1451 and w2285;
w6416 <= w6414 and not w6415;
w6417 <= a(26) and not w6416;
w6418 <= a(26) and not w6417;
w6419 <= not w6416 and not w6417;
w6420 <= not w6418 and not w6419;
w6421 <= w6409 and not w6420;
w6422 <= w6409 and not w6421;
w6423 <= not w6420 and not w6421;
w6424 <= not w6422 and not w6423;
w6425 <= not w6134 and not w6137;
w6426 <= w6424 and w6425;
w6427 <= not w6424 and not w6425;
w6428 <= not w6426 and not w6427;
w6429 <= b(22) and w1791;
w6430 <= b(20) and w1941;
w6431 <= b(21) and w1786;
w6432 <= not w6430 and not w6431;
w6433 <= not w6429 and w6432;
w6434 <= w1794 and w1888;
w6435 <= w6433 and not w6434;
w6436 <= a(23) and not w6435;
w6437 <= a(23) and not w6436;
w6438 <= not w6435 and not w6436;
w6439 <= not w6437 and not w6438;
w6440 <= w6428 and not w6439;
w6441 <= w6428 and not w6440;
w6442 <= not w6439 and not w6440;
w6443 <= not w6441 and not w6442;
w6444 <= not w6140 and not w6146;
w6445 <= w6443 and w6444;
w6446 <= not w6443 and not w6444;
w6447 <= not w6445 and not w6446;
w6448 <= b(25) and w1370;
w6449 <= b(23) and w1506;
w6450 <= b(24) and w1365;
w6451 <= not w6449 and not w6450;
w6452 <= not w6448 and w6451;
w6453 <= w1373 and w2228;
w6454 <= w6452 and not w6453;
w6455 <= a(20) and not w6454;
w6456 <= a(20) and not w6455;
w6457 <= not w6454 and not w6455;
w6458 <= not w6456 and not w6457;
w6459 <= w6447 and not w6458;
w6460 <= w6447 and not w6459;
w6461 <= not w6458 and not w6459;
w6462 <= not w6460 and not w6461;
w6463 <= not w6160 and not w6162;
w6464 <= not w6462 and not w6463;
w6465 <= w6462 and w6463;
w6466 <= not w6464 and not w6465;
w6467 <= not w6291 and w6466;
w6468 <= not w6291 and not w6467;
w6469 <= w6466 and not w6467;
w6470 <= not w6468 and not w6469;
w6471 <= not w6280 and not w6470;
w6472 <= not w6280 and not w6471;
w6473 <= not w6470 and not w6471;
w6474 <= not w6472 and not w6473;
w6475 <= b(31) and w694;
w6476 <= b(29) and w799;
w6477 <= b(30) and w689;
w6478 <= not w6476 and not w6477;
w6479 <= not w6475 and w6478;
w6480 <= w697 and w3539;
w6481 <= w6479 and not w6480;
w6482 <= a(14) and not w6481;
w6483 <= a(14) and not w6482;
w6484 <= not w6481 and not w6482;
w6485 <= not w6483 and not w6484;
w6486 <= w6474 and w6485;
w6487 <= not w6474 and not w6485;
w6488 <= not w6486 and not w6487;
w6489 <= not w6278 and w6488;
w6490 <= w6278 and not w6488;
w6491 <= not w6489 and not w6490;
w6492 <= not w6277 and w6491;
w6493 <= w6491 and not w6492;
w6494 <= not w6277 and not w6492;
w6495 <= not w6493 and not w6494;
w6496 <= not w5989 and not w6192;
w6497 <= not w6189 and not w6496;
w6498 <= w6495 and w6497;
w6499 <= not w6495 and not w6497;
w6500 <= not w6498 and not w6499;
w6501 <= b(37) and w254;
w6502 <= b(35) and w284;
w6503 <= b(36) and w249;
w6504 <= not w6502 and not w6503;
w6505 <= not w6501 and w6504;
w6506 <= w257 and w4924;
w6507 <= w6505 and not w6506;
w6508 <= a(8) and not w6507;
w6509 <= a(8) and not w6508;
w6510 <= not w6507 and not w6508;
w6511 <= not w6509 and not w6510;
w6512 <= w6500 and not w6511;
w6513 <= not w6500 and w6511;
w6514 <= not w6266 and not w6513;
w6515 <= not w6512 and w6514;
w6516 <= not w6266 and not w6515;
w6517 <= not w6512 and not w6515;
w6518 <= not w6513 and w6517;
w6519 <= not w6516 and not w6518;
w6520 <= b(40) and w105;
w6521 <= b(38) and w146;
w6522 <= b(39) and w100;
w6523 <= not w6521 and not w6522;
w6524 <= not w6520 and w6523;
w6525 <= w108 and w5698;
w6526 <= w6524 and not w6525;
w6527 <= a(5) and not w6526;
w6528 <= a(5) and not w6527;
w6529 <= not w6526 and not w6527;
w6530 <= not w6528 and not w6529;
w6531 <= w6519 and w6530;
w6532 <= not w6519 and not w6530;
w6533 <= not w6531 and not w6532;
w6534 <= not w6265 and w6533;
w6535 <= w6265 and not w6533;
w6536 <= not w6534 and not w6535;
w6537 <= not w6264 and w6536;
w6538 <= w6536 and not w6537;
w6539 <= not w6264 and not w6537;
w6540 <= not w6538 and not w6539;
w6541 <= not w6239 and not w6244;
w6542 <= not w6540 and not w6541;
w6543 <= w6540 and w6541;
w6544 <= not w6542 and not w6543;
w6545 <= not w6537 and not w6542;
w6546 <= not w6532 and not w6534;
w6547 <= b(41) and w105;
w6548 <= b(39) and w146;
w6549 <= b(40) and w100;
w6550 <= not w6548 and not w6549;
w6551 <= not w6547 and w6550;
w6552 <= w108 and w5962;
w6553 <= w6551 and not w6552;
w6554 <= a(5) and not w6553;
w6555 <= a(5) and not w6554;
w6556 <= not w6553 and not w6554;
w6557 <= not w6555 and not w6556;
w6558 <= b(35) and w443;
w6559 <= b(33) and w510;
w6560 <= b(34) and w438;
w6561 <= not w6559 and not w6560;
w6562 <= not w6558 and w6561;
w6563 <= w446 and w4439;
w6564 <= w6562 and not w6563;
w6565 <= a(11) and not w6564;
w6566 <= a(11) and not w6565;
w6567 <= not w6564 and not w6565;
w6568 <= not w6566 and not w6567;
w6569 <= not w6487 and not w6489;
w6570 <= b(32) and w694;
w6571 <= b(30) and w799;
w6572 <= b(31) and w689;
w6573 <= not w6571 and not w6572;
w6574 <= not w6570 and w6573;
w6575 <= w697 and w3756;
w6576 <= w6574 and not w6575;
w6577 <= a(14) and not w6576;
w6578 <= a(14) and not w6577;
w6579 <= not w6576 and not w6577;
w6580 <= not w6578 and not w6579;
w6581 <= not w6467 and not w6471;
w6582 <= b(29) and w1045;
w6583 <= b(27) and w1134;
w6584 <= b(28) and w1040;
w6585 <= not w6583 and not w6584;
w6586 <= not w6582 and w6585;
w6587 <= w1048 and w3126;
w6588 <= w6586 and not w6587;
w6589 <= a(17) and not w6588;
w6590 <= a(17) and not w6589;
w6591 <= not w6588 and not w6589;
w6592 <= not w6590 and not w6591;
w6593 <= not w6459 and not w6464;
w6594 <= not w6440 and not w6446;
w6595 <= b(20) and w2282;
w6596 <= b(18) and w2428;
w6597 <= b(19) and w2277;
w6598 <= not w6596 and not w6597;
w6599 <= not w6595 and w6598;
w6600 <= w1589 and w2285;
w6601 <= w6599 and not w6600;
w6602 <= a(26) and not w6601;
w6603 <= a(26) and not w6602;
w6604 <= not w6601 and not w6602;
w6605 <= not w6603 and not w6604;
w6606 <= not w6401 and not w6408;
w6607 <= b(17) and w2793;
w6608 <= b(15) and w2986;
w6609 <= b(16) and w2788;
w6610 <= not w6608 and not w6609;
w6611 <= not w6607 and w6610;
w6612 <= w1099 and w2796;
w6613 <= w6611 and not w6612;
w6614 <= a(29) and not w6613;
w6615 <= a(29) and not w6614;
w6616 <= not w6613 and not w6614;
w6617 <= not w6615 and not w6616;
w6618 <= not w6396 and not w6398;
w6619 <= b(14) and w3381;
w6620 <= b(12) and w3586;
w6621 <= b(13) and w3376;
w6622 <= not w6620 and not w6621;
w6623 <= not w6619 and w6622;
w6624 <= w777 and w3384;
w6625 <= w6623 and not w6624;
w6626 <= a(32) and not w6625;
w6627 <= a(32) and not w6626;
w6628 <= not w6625 and not w6626;
w6629 <= not w6627 and not w6628;
w6630 <= not w6357 and not w6363;
w6631 <= b(8) and w4778;
w6632 <= b(6) and w5020;
w6633 <= b(7) and w4773;
w6634 <= not w6632 and not w6633;
w6635 <= not w6631 and w6634;
w6636 <= w328 and w4781;
w6637 <= w6635 and not w6636;
w6638 <= a(38) and not w6637;
w6639 <= a(38) and not w6638;
w6640 <= not w6637 and not w6638;
w6641 <= not w6639 and not w6640;
w6642 <= not w6352 and not w6354;
w6643 <= b(2) and w6338;
w6644 <= w6053 and not w6337;
w6645 <= w6332 and w6644;
w6646 <= b(0) and w6645;
w6647 <= b(1) and w6333;
w6648 <= not w6646 and not w6647;
w6649 <= not w6643 and w6648;
w6650 <= w39 and w6341;
w6651 <= w6649 and not w6650;
w6652 <= a(44) and not w6651;
w6653 <= a(44) and not w6652;
w6654 <= not w6651 and not w6652;
w6655 <= not w6653 and not w6654;
w6656 <= not w6348 and w6655;
w6657 <= w6348 and not w6655;
w6658 <= not w6656 and not w6657;
w6659 <= b(5) and w5520;
w6660 <= b(3) and w5802;
w6661 <= b(4) and w5515;
w6662 <= not w6660 and not w6661;
w6663 <= not w6659 and w6662;
w6664 <= w137 and w5523;
w6665 <= w6663 and not w6664;
w6666 <= a(41) and not w6665;
w6667 <= a(41) and not w6666;
w6668 <= not w6665 and not w6666;
w6669 <= not w6667 and not w6668;
w6670 <= w6658 and not w6669;
w6671 <= w6658 and not w6670;
w6672 <= not w6669 and not w6670;
w6673 <= not w6671 and not w6672;
w6674 <= not w6642 and not w6673;
w6675 <= w6642 and w6673;
w6676 <= not w6674 and not w6675;
w6677 <= not w6641 and w6676;
w6678 <= not w6641 and not w6677;
w6679 <= w6676 and not w6677;
w6680 <= not w6678 and not w6679;
w6681 <= not w6630 and not w6680;
w6682 <= not w6630 and not w6681;
w6683 <= not w6680 and not w6681;
w6684 <= not w6682 and not w6683;
w6685 <= b(11) and w4030;
w6686 <= b(9) and w4275;
w6687 <= b(10) and w4025;
w6688 <= not w6686 and not w6687;
w6689 <= not w6685 and w6688;
w6690 <= w561 and w4033;
w6691 <= w6689 and not w6690;
w6692 <= a(35) and not w6691;
w6693 <= a(35) and not w6692;
w6694 <= not w6691 and not w6692;
w6695 <= not w6693 and not w6694;
w6696 <= w6684 and w6695;
w6697 <= not w6684 and not w6695;
w6698 <= not w6696 and not w6697;
w6699 <= not w6381 and w6698;
w6700 <= w6381 and not w6698;
w6701 <= not w6699 and not w6700;
w6702 <= w6629 and not w6701;
w6703 <= not w6629 and w6701;
w6704 <= not w6702 and not w6703;
w6705 <= not w6618 and w6704;
w6706 <= w6618 and not w6704;
w6707 <= not w6705 and not w6706;
w6708 <= w6617 and not w6707;
w6709 <= not w6617 and w6707;
w6710 <= not w6708 and not w6709;
w6711 <= not w6606 and w6710;
w6712 <= w6606 and not w6710;
w6713 <= not w6711 and not w6712;
w6714 <= not w6605 and w6713;
w6715 <= w6713 and not w6714;
w6716 <= not w6605 and not w6714;
w6717 <= not w6715 and not w6716;
w6718 <= not w6421 and not w6427;
w6719 <= w6717 and w6718;
w6720 <= not w6717 and not w6718;
w6721 <= not w6719 and not w6720;
w6722 <= b(23) and w1791;
w6723 <= b(21) and w1941;
w6724 <= b(22) and w1786;
w6725 <= not w6723 and not w6724;
w6726 <= not w6722 and w6725;
w6727 <= w1794 and w2043;
w6728 <= w6726 and not w6727;
w6729 <= a(23) and not w6728;
w6730 <= a(23) and not w6729;
w6731 <= not w6728 and not w6729;
w6732 <= not w6730 and not w6731;
w6733 <= w6721 and not w6732;
w6734 <= not w6721 and w6732;
w6735 <= not w6594 and not w6734;
w6736 <= not w6733 and w6735;
w6737 <= not w6594 and not w6736;
w6738 <= not w6733 and not w6736;
w6739 <= not w6734 and w6738;
w6740 <= not w6737 and not w6739;
w6741 <= b(26) and w1370;
w6742 <= b(24) and w1506;
w6743 <= b(25) and w1365;
w6744 <= not w6742 and not w6743;
w6745 <= not w6741 and w6744;
w6746 <= w1373 and w2556;
w6747 <= w6745 and not w6746;
w6748 <= a(20) and not w6747;
w6749 <= a(20) and not w6748;
w6750 <= not w6747 and not w6748;
w6751 <= not w6749 and not w6750;
w6752 <= w6740 and w6751;
w6753 <= not w6740 and not w6751;
w6754 <= not w6752 and not w6753;
w6755 <= not w6593 and w6754;
w6756 <= w6593 and not w6754;
w6757 <= not w6755 and not w6756;
w6758 <= w6592 and not w6757;
w6759 <= not w6592 and w6757;
w6760 <= not w6758 and not w6759;
w6761 <= not w6581 and w6760;
w6762 <= w6581 and not w6760;
w6763 <= not w6761 and not w6762;
w6764 <= w6580 and not w6763;
w6765 <= not w6580 and w6763;
w6766 <= not w6764 and not w6765;
w6767 <= not w6569 and w6766;
w6768 <= w6569 and not w6766;
w6769 <= not w6767 and not w6768;
w6770 <= not w6568 and w6769;
w6771 <= w6769 and not w6770;
w6772 <= not w6568 and not w6770;
w6773 <= not w6771 and not w6772;
w6774 <= not w6492 and not w6499;
w6775 <= w6773 and w6774;
w6776 <= not w6773 and not w6774;
w6777 <= not w6775 and not w6776;
w6778 <= b(38) and w254;
w6779 <= b(36) and w284;
w6780 <= b(37) and w249;
w6781 <= not w6779 and not w6780;
w6782 <= not w6778 and w6781;
w6783 <= w257 and w4948;
w6784 <= w6782 and not w6783;
w6785 <= a(8) and not w6784;
w6786 <= a(8) and not w6785;
w6787 <= not w6784 and not w6785;
w6788 <= not w6786 and not w6787;
w6789 <= w6777 and not w6788;
w6790 <= w6777 and not w6789;
w6791 <= not w6788 and not w6789;
w6792 <= not w6790 and not w6791;
w6793 <= not w6517 and not w6792;
w6794 <= w6517 and w6792;
w6795 <= not w6793 and not w6794;
w6796 <= not w6557 and w6795;
w6797 <= not w6557 and not w6796;
w6798 <= w6795 and not w6796;
w6799 <= not w6797 and not w6798;
w6800 <= not w6546 and not w6799;
w6801 <= not w6546 and not w6800;
w6802 <= not w6799 and not w6800;
w6803 <= not w6801 and not w6802;
w6804 <= b(44) and w9;
w6805 <= b(42) and w27;
w6806 <= b(43) and w4;
w6807 <= not w6805 and not w6806;
w6808 <= not w6804 and w6807;
w6809 <= not w6254 and not w6256;
w6810 <= not b(43) and not b(44);
w6811 <= b(43) and b(44);
w6812 <= not w6810 and not w6811;
w6813 <= not w6809 and w6812;
w6814 <= w6809 and not w6812;
w6815 <= not w6813 and not w6814;
w6816 <= w12 and w6815;
w6817 <= w6808 and not w6816;
w6818 <= a(2) and not w6817;
w6819 <= a(2) and not w6818;
w6820 <= not w6817 and not w6818;
w6821 <= not w6819 and not w6820;
w6822 <= not w6803 and w6821;
w6823 <= w6803 and not w6821;
w6824 <= not w6822 and not w6823;
w6825 <= not w6545 and not w6824;
w6826 <= w6545 and w6824;
w6827 <= not w6825 and not w6826;
w6828 <= not w6803 and not w6821;
w6829 <= not w6825 and not w6828;
w6830 <= not w6770 and not w6776;
w6831 <= not w6765 and not w6767;
w6832 <= b(33) and w694;
w6833 <= b(31) and w799;
w6834 <= b(32) and w689;
w6835 <= not w6833 and not w6834;
w6836 <= not w6832 and w6835;
w6837 <= w697 and w3966;
w6838 <= w6836 and not w6837;
w6839 <= a(14) and not w6838;
w6840 <= a(14) and not w6839;
w6841 <= not w6838 and not w6839;
w6842 <= not w6840 and not w6841;
w6843 <= not w6759 and not w6761;
w6844 <= not w6753 and not w6755;
w6845 <= b(27) and w1370;
w6846 <= b(25) and w1506;
w6847 <= b(26) and w1365;
w6848 <= not w6846 and not w6847;
w6849 <= not w6845 and w6848;
w6850 <= w1373 and w2733;
w6851 <= w6849 and not w6850;
w6852 <= a(20) and not w6851;
w6853 <= a(20) and not w6852;
w6854 <= not w6851 and not w6852;
w6855 <= not w6853 and not w6854;
w6856 <= b(21) and w2282;
w6857 <= b(19) and w2428;
w6858 <= b(20) and w2277;
w6859 <= not w6857 and not w6858;
w6860 <= not w6856 and w6859;
w6861 <= w1727 and w2285;
w6862 <= w6860 and not w6861;
w6863 <= a(26) and not w6862;
w6864 <= a(26) and not w6863;
w6865 <= not w6862 and not w6863;
w6866 <= not w6864 and not w6865;
w6867 <= not w6709 and not w6711;
w6868 <= not w6703 and not w6705;
w6869 <= not w6697 and not w6699;
w6870 <= b(12) and w4030;
w6871 <= b(10) and w4275;
w6872 <= b(11) and w4025;
w6873 <= not w6871 and not w6872;
w6874 <= not w6870 and w6873;
w6875 <= w585 and w4033;
w6876 <= w6874 and not w6875;
w6877 <= a(35) and not w6876;
w6878 <= a(35) and not w6877;
w6879 <= not w6876 and not w6877;
w6880 <= not w6878 and not w6879;
w6881 <= not w6677 and not w6681;
w6882 <= b(6) and w5520;
w6883 <= b(4) and w5802;
w6884 <= b(5) and w5515;
w6885 <= not w6883 and not w6884;
w6886 <= not w6882 and w6885;
w6887 <= w202 and w5523;
w6888 <= w6886 and not w6887;
w6889 <= a(41) and not w6888;
w6890 <= a(41) and not w6889;
w6891 <= not w6888 and not w6889;
w6892 <= not w6890 and not w6891;
w6893 <= a(44) and not a(45);
w6894 <= not a(44) and a(45);
w6895 <= not w6893 and not w6894;
w6896 <= b(0) and not w6895;
w6897 <= not w6657 and w6896;
w6898 <= w6657 and not w6896;
w6899 <= not w6897 and not w6898;
w6900 <= b(3) and w6338;
w6901 <= b(1) and w6645;
w6902 <= b(2) and w6333;
w6903 <= not w6901 and not w6902;
w6904 <= not w6900 and w6903;
w6905 <= w61 and w6341;
w6906 <= w6904 and not w6905;
w6907 <= a(44) and not w6906;
w6908 <= a(44) and not w6907;
w6909 <= not w6906 and not w6907;
w6910 <= not w6908 and not w6909;
w6911 <= not w6899 and not w6910;
w6912 <= w6899 and w6910;
w6913 <= not w6911 and not w6912;
w6914 <= not w6892 and w6913;
w6915 <= w6913 and not w6914;
w6916 <= not w6892 and not w6914;
w6917 <= not w6915 and not w6916;
w6918 <= not w6670 and not w6674;
w6919 <= w6917 and w6918;
w6920 <= not w6917 and not w6918;
w6921 <= not w6919 and not w6920;
w6922 <= b(9) and w4778;
w6923 <= b(7) and w5020;
w6924 <= b(8) and w4773;
w6925 <= not w6923 and not w6924;
w6926 <= not w6922 and w6925;
w6927 <= w394 and w4781;
w6928 <= w6926 and not w6927;
w6929 <= a(38) and not w6928;
w6930 <= a(38) and not w6929;
w6931 <= not w6928 and not w6929;
w6932 <= not w6930 and not w6931;
w6933 <= not w6921 and w6932;
w6934 <= w6921 and not w6932;
w6935 <= not w6933 and not w6934;
w6936 <= not w6881 and w6935;
w6937 <= w6881 and not w6935;
w6938 <= not w6936 and not w6937;
w6939 <= not w6880 and w6938;
w6940 <= not w6880 and not w6939;
w6941 <= w6938 and not w6939;
w6942 <= not w6940 and not w6941;
w6943 <= not w6869 and not w6942;
w6944 <= not w6869 and not w6943;
w6945 <= not w6942 and not w6943;
w6946 <= not w6944 and not w6945;
w6947 <= b(15) and w3381;
w6948 <= b(13) and w3586;
w6949 <= b(14) and w3376;
w6950 <= not w6948 and not w6949;
w6951 <= not w6947 and w6950;
w6952 <= w874 and w3384;
w6953 <= w6951 and not w6952;
w6954 <= a(32) and not w6953;
w6955 <= a(32) and not w6954;
w6956 <= not w6953 and not w6954;
w6957 <= not w6955 and not w6956;
w6958 <= not w6946 and not w6957;
w6959 <= not w6946 and not w6958;
w6960 <= not w6957 and not w6958;
w6961 <= not w6959 and not w6960;
w6962 <= not w6868 and w6961;
w6963 <= w6868 and not w6961;
w6964 <= not w6962 and not w6963;
w6965 <= b(18) and w2793;
w6966 <= b(16) and w2986;
w6967 <= b(17) and w2788;
w6968 <= not w6966 and not w6967;
w6969 <= not w6965 and w6968;
w6970 <= w1309 and w2796;
w6971 <= w6969 and not w6970;
w6972 <= a(29) and not w6971;
w6973 <= a(29) and not w6972;
w6974 <= not w6971 and not w6972;
w6975 <= not w6973 and not w6974;
w6976 <= not w6964 and not w6975;
w6977 <= w6964 and w6975;
w6978 <= not w6976 and not w6977;
w6979 <= not w6867 and w6978;
w6980 <= w6867 and not w6978;
w6981 <= not w6979 and not w6980;
w6982 <= not w6866 and w6981;
w6983 <= w6981 and not w6982;
w6984 <= not w6866 and not w6982;
w6985 <= not w6983 and not w6984;
w6986 <= not w6714 and not w6720;
w6987 <= w6985 and w6986;
w6988 <= not w6985 and not w6986;
w6989 <= not w6987 and not w6988;
w6990 <= b(24) and w1791;
w6991 <= b(22) and w1941;
w6992 <= b(23) and w1786;
w6993 <= not w6991 and not w6992;
w6994 <= not w6990 and w6993;
w6995 <= w1794 and w2201;
w6996 <= w6994 and not w6995;
w6997 <= a(23) and not w6996;
w6998 <= a(23) and not w6997;
w6999 <= not w6996 and not w6997;
w7000 <= not w6998 and not w6999;
w7001 <= not w6989 and w7000;
w7002 <= w6989 and not w7000;
w7003 <= not w7001 and not w7002;
w7004 <= not w6738 and w7003;
w7005 <= w6738 and not w7003;
w7006 <= not w7004 and not w7005;
w7007 <= not w6855 and w7006;
w7008 <= w7006 and not w7007;
w7009 <= not w6855 and not w7007;
w7010 <= not w7008 and not w7009;
w7011 <= not w6844 and w7010;
w7012 <= w6844 and not w7010;
w7013 <= not w7011 and not w7012;
w7014 <= b(30) and w1045;
w7015 <= b(28) and w1134;
w7016 <= b(29) and w1040;
w7017 <= not w7015 and not w7016;
w7018 <= not w7014 and w7017;
w7019 <= w1048 and w3320;
w7020 <= w7018 and not w7019;
w7021 <= a(17) and not w7020;
w7022 <= a(17) and not w7021;
w7023 <= not w7020 and not w7021;
w7024 <= not w7022 and not w7023;
w7025 <= not w7013 and not w7024;
w7026 <= w7013 and w7024;
w7027 <= not w7025 and not w7026;
w7028 <= not w6843 and w7027;
w7029 <= w6843 and not w7027;
w7030 <= not w7028 and not w7029;
w7031 <= not w6842 and w7030;
w7032 <= w7030 and not w7031;
w7033 <= not w6842 and not w7031;
w7034 <= not w7032 and not w7033;
w7035 <= not w6831 and w7034;
w7036 <= w6831 and not w7034;
w7037 <= not w7035 and not w7036;
w7038 <= b(36) and w443;
w7039 <= b(34) and w510;
w7040 <= b(35) and w438;
w7041 <= not w7039 and not w7040;
w7042 <= not w7038 and w7041;
w7043 <= w446 and w4665;
w7044 <= w7042 and not w7043;
w7045 <= a(11) and not w7044;
w7046 <= a(11) and not w7045;
w7047 <= not w7044 and not w7045;
w7048 <= not w7046 and not w7047;
w7049 <= not w7037 and not w7048;
w7050 <= w7037 and w7048;
w7051 <= not w7049 and not w7050;
w7052 <= w6830 and not w7051;
w7053 <= not w6830 and w7051;
w7054 <= not w7052 and not w7053;
w7055 <= b(39) and w254;
w7056 <= b(37) and w284;
w7057 <= b(38) and w249;
w7058 <= not w7056 and not w7057;
w7059 <= not w7055 and w7058;
w7060 <= w257 and w5194;
w7061 <= w7059 and not w7060;
w7062 <= a(8) and not w7061;
w7063 <= a(8) and not w7062;
w7064 <= not w7061 and not w7062;
w7065 <= not w7063 and not w7064;
w7066 <= w7054 and not w7065;
w7067 <= w7054 and not w7066;
w7068 <= not w7065 and not w7066;
w7069 <= not w7067 and not w7068;
w7070 <= not w6789 and not w6793;
w7071 <= w7069 and w7070;
w7072 <= not w7069 and not w7070;
w7073 <= not w7071 and not w7072;
w7074 <= b(42) and w105;
w7075 <= b(40) and w146;
w7076 <= b(41) and w100;
w7077 <= not w7075 and not w7076;
w7078 <= not w7074 and w7077;
w7079 <= w108 and w6232;
w7080 <= w7078 and not w7079;
w7081 <= a(5) and not w7080;
w7082 <= a(5) and not w7081;
w7083 <= not w7080 and not w7081;
w7084 <= not w7082 and not w7083;
w7085 <= w7073 and not w7084;
w7086 <= w7073 and not w7085;
w7087 <= not w7084 and not w7085;
w7088 <= not w7086 and not w7087;
w7089 <= not w6796 and not w6800;
w7090 <= w7088 and w7089;
w7091 <= not w7088 and not w7089;
w7092 <= not w7090 and not w7091;
w7093 <= b(45) and w9;
w7094 <= b(43) and w27;
w7095 <= b(44) and w4;
w7096 <= not w7094 and not w7095;
w7097 <= not w7093 and w7096;
w7098 <= not w6811 and not w6813;
w7099 <= not b(44) and not b(45);
w7100 <= b(44) and b(45);
w7101 <= not w7099 and not w7100;
w7102 <= not w7098 and w7101;
w7103 <= w7098 and not w7101;
w7104 <= not w7102 and not w7103;
w7105 <= w12 and w7104;
w7106 <= w7097 and not w7105;
w7107 <= a(2) and not w7106;
w7108 <= a(2) and not w7107;
w7109 <= not w7106 and not w7107;
w7110 <= not w7108 and not w7109;
w7111 <= not w7092 and w7110;
w7112 <= w7092 and not w7110;
w7113 <= not w7111 and not w7112;
w7114 <= not w6829 and w7113;
w7115 <= w6829 and not w7113;
w7116 <= not w7114 and not w7115;
w7117 <= not w7066 and not w7072;
w7118 <= b(34) and w694;
w7119 <= b(32) and w799;
w7120 <= b(33) and w689;
w7121 <= not w7119 and not w7120;
w7122 <= not w7118 and w7121;
w7123 <= w697 and w4209;
w7124 <= w7122 and not w7123;
w7125 <= a(14) and not w7124;
w7126 <= a(14) and not w7125;
w7127 <= not w7124 and not w7125;
w7128 <= not w7126 and not w7127;
w7129 <= not w7025 and not w7028;
w7130 <= not w6844 and not w7010;
w7131 <= not w7007 and not w7130;
w7132 <= b(28) and w1370;
w7133 <= b(26) and w1506;
w7134 <= b(27) and w1365;
w7135 <= not w7133 and not w7134;
w7136 <= not w7132 and w7135;
w7137 <= w1373 and w2932;
w7138 <= w7136 and not w7137;
w7139 <= a(20) and not w7138;
w7140 <= a(20) and not w7139;
w7141 <= not w7138 and not w7139;
w7142 <= not w7140 and not w7141;
w7143 <= b(16) and w3381;
w7144 <= b(14) and w3586;
w7145 <= b(15) and w3376;
w7146 <= not w7144 and not w7145;
w7147 <= not w7143 and w7146;
w7148 <= w980 and w3384;
w7149 <= w7147 and not w7148;
w7150 <= a(32) and not w7149;
w7151 <= a(32) and not w7150;
w7152 <= not w7149 and not w7150;
w7153 <= not w7151 and not w7152;
w7154 <= not w6939 and not w6943;
w7155 <= not w6934 and not w6936;
w7156 <= b(7) and w5520;
w7157 <= b(5) and w5802;
w7158 <= b(6) and w5515;
w7159 <= not w7157 and not w7158;
w7160 <= not w7156 and w7159;
w7161 <= w227 and w5523;
w7162 <= w7160 and not w7161;
w7163 <= a(41) and not w7162;
w7164 <= a(41) and not w7163;
w7165 <= not w7162 and not w7163;
w7166 <= not w7164 and not w7165;
w7167 <= w6657 and w6896;
w7168 <= not w6911 and not w7167;
w7169 <= b(4) and w6338;
w7170 <= b(2) and w6645;
w7171 <= b(3) and w6333;
w7172 <= not w7170 and not w7171;
w7173 <= not w7169 and w7172;
w7174 <= w89 and w6341;
w7175 <= w7173 and not w7174;
w7176 <= a(44) and not w7175;
w7177 <= a(44) and not w7176;
w7178 <= not w7175 and not w7176;
w7179 <= not w7177 and not w7178;
w7180 <= a(47) and not w6896;
w7181 <= not a(45) and a(46);
w7182 <= a(45) and not a(46);
w7183 <= not w7181 and not w7182;
w7184 <= w6895 and not w7183;
w7185 <= b(0) and w7184;
w7186 <= not a(46) and a(47);
w7187 <= a(46) and not a(47);
w7188 <= not w7186 and not w7187;
w7189 <= not w6895 and w7188;
w7190 <= b(1) and w7189;
w7191 <= not w7185 and not w7190;
w7192 <= not w6895 and not w7188;
w7193 <= not w15 and w7192;
w7194 <= w7191 and not w7193;
w7195 <= a(47) and not w7194;
w7196 <= a(47) and not w7195;
w7197 <= not w7194 and not w7195;
w7198 <= not w7196 and not w7197;
w7199 <= w7180 and not w7198;
w7200 <= not w7180 and w7198;
w7201 <= not w7199 and not w7200;
w7202 <= w7179 and not w7201;
w7203 <= not w7179 and w7201;
w7204 <= not w7202 and not w7203;
w7205 <= not w7168 and w7204;
w7206 <= w7168 and not w7204;
w7207 <= not w7205 and not w7206;
w7208 <= not w7166 and w7207;
w7209 <= w7207 and not w7208;
w7210 <= not w7166 and not w7208;
w7211 <= not w7209 and not w7210;
w7212 <= not w6914 and not w6920;
w7213 <= w7211 and w7212;
w7214 <= not w7211 and not w7212;
w7215 <= not w7213 and not w7214;
w7216 <= b(10) and w4778;
w7217 <= b(8) and w5020;
w7218 <= b(9) and w4773;
w7219 <= not w7217 and not w7218;
w7220 <= not w7216 and w7219;
w7221 <= w481 and w4781;
w7222 <= w7220 and not w7221;
w7223 <= a(38) and not w7222;
w7224 <= a(38) and not w7223;
w7225 <= not w7222 and not w7223;
w7226 <= not w7224 and not w7225;
w7227 <= w7215 and not w7226;
w7228 <= not w7215 and w7226;
w7229 <= not w7155 and not w7228;
w7230 <= not w7227 and w7229;
w7231 <= not w7155 and not w7230;
w7232 <= not w7227 and not w7230;
w7233 <= not w7228 and w7232;
w7234 <= not w7231 and not w7233;
w7235 <= b(13) and w4030;
w7236 <= b(11) and w4275;
w7237 <= b(12) and w4025;
w7238 <= not w7236 and not w7237;
w7239 <= not w7235 and w7238;
w7240 <= w751 and w4033;
w7241 <= w7239 and not w7240;
w7242 <= a(35) and not w7241;
w7243 <= a(35) and not w7242;
w7244 <= not w7241 and not w7242;
w7245 <= not w7243 and not w7244;
w7246 <= w7234 and w7245;
w7247 <= not w7234 and not w7245;
w7248 <= not w7246 and not w7247;
w7249 <= not w7154 and w7248;
w7250 <= w7154 and not w7248;
w7251 <= not w7249 and not w7250;
w7252 <= not w7153 and w7251;
w7253 <= w7251 and not w7252;
w7254 <= not w7153 and not w7252;
w7255 <= not w7253 and not w7254;
w7256 <= not w6868 and not w6961;
w7257 <= not w6958 and not w7256;
w7258 <= w7255 and w7257;
w7259 <= not w7255 and not w7257;
w7260 <= not w7258 and not w7259;
w7261 <= b(19) and w2793;
w7262 <= b(17) and w2986;
w7263 <= b(18) and w2788;
w7264 <= not w7262 and not w7263;
w7265 <= not w7261 and w7264;
w7266 <= w1451 and w2796;
w7267 <= w7265 and not w7266;
w7268 <= a(29) and not w7267;
w7269 <= a(29) and not w7268;
w7270 <= not w7267 and not w7268;
w7271 <= not w7269 and not w7270;
w7272 <= w7260 and not w7271;
w7273 <= w7260 and not w7272;
w7274 <= not w7271 and not w7272;
w7275 <= not w7273 and not w7274;
w7276 <= not w6976 and not w6979;
w7277 <= w7275 and w7276;
w7278 <= not w7275 and not w7276;
w7279 <= not w7277 and not w7278;
w7280 <= b(22) and w2282;
w7281 <= b(20) and w2428;
w7282 <= b(21) and w2277;
w7283 <= not w7281 and not w7282;
w7284 <= not w7280 and w7283;
w7285 <= w1888 and w2285;
w7286 <= w7284 and not w7285;
w7287 <= a(26) and not w7286;
w7288 <= a(26) and not w7287;
w7289 <= not w7286 and not w7287;
w7290 <= not w7288 and not w7289;
w7291 <= w7279 and not w7290;
w7292 <= w7279 and not w7291;
w7293 <= not w7290 and not w7291;
w7294 <= not w7292 and not w7293;
w7295 <= not w6982 and not w6988;
w7296 <= w7294 and w7295;
w7297 <= not w7294 and not w7295;
w7298 <= not w7296 and not w7297;
w7299 <= b(25) and w1791;
w7300 <= b(23) and w1941;
w7301 <= b(24) and w1786;
w7302 <= not w7300 and not w7301;
w7303 <= not w7299 and w7302;
w7304 <= w1794 and w2228;
w7305 <= w7303 and not w7304;
w7306 <= a(23) and not w7305;
w7307 <= a(23) and not w7306;
w7308 <= not w7305 and not w7306;
w7309 <= not w7307 and not w7308;
w7310 <= w7298 and not w7309;
w7311 <= w7298 and not w7310;
w7312 <= not w7309 and not w7310;
w7313 <= not w7311 and not w7312;
w7314 <= not w7002 and not w7004;
w7315 <= not w7313 and not w7314;
w7316 <= w7313 and w7314;
w7317 <= not w7315 and not w7316;
w7318 <= not w7142 and w7317;
w7319 <= not w7142 and not w7318;
w7320 <= w7317 and not w7318;
w7321 <= not w7319 and not w7320;
w7322 <= not w7131 and not w7321;
w7323 <= not w7131 and not w7322;
w7324 <= not w7321 and not w7322;
w7325 <= not w7323 and not w7324;
w7326 <= b(31) and w1045;
w7327 <= b(29) and w1134;
w7328 <= b(30) and w1040;
w7329 <= not w7327 and not w7328;
w7330 <= not w7326 and w7329;
w7331 <= w1048 and w3539;
w7332 <= w7330 and not w7331;
w7333 <= a(17) and not w7332;
w7334 <= a(17) and not w7333;
w7335 <= not w7332 and not w7333;
w7336 <= not w7334 and not w7335;
w7337 <= w7325 and w7336;
w7338 <= not w7325 and not w7336;
w7339 <= not w7337 and not w7338;
w7340 <= not w7129 and w7339;
w7341 <= w7129 and not w7339;
w7342 <= not w7340 and not w7341;
w7343 <= not w7128 and w7342;
w7344 <= w7342 and not w7343;
w7345 <= not w7128 and not w7343;
w7346 <= not w7344 and not w7345;
w7347 <= not w6831 and not w7034;
w7348 <= not w7031 and not w7347;
w7349 <= w7346 and w7348;
w7350 <= not w7346 and not w7348;
w7351 <= not w7349 and not w7350;
w7352 <= b(37) and w443;
w7353 <= b(35) and w510;
w7354 <= b(36) and w438;
w7355 <= not w7353 and not w7354;
w7356 <= not w7352 and w7355;
w7357 <= w446 and w4924;
w7358 <= w7356 and not w7357;
w7359 <= a(11) and not w7358;
w7360 <= a(11) and not w7359;
w7361 <= not w7358 and not w7359;
w7362 <= not w7360 and not w7361;
w7363 <= w7351 and not w7362;
w7364 <= w7351 and not w7363;
w7365 <= not w7362 and not w7363;
w7366 <= not w7364 and not w7365;
w7367 <= not w7049 and not w7053;
w7368 <= w7366 and w7367;
w7369 <= not w7366 and not w7367;
w7370 <= not w7368 and not w7369;
w7371 <= b(40) and w254;
w7372 <= b(38) and w284;
w7373 <= b(39) and w249;
w7374 <= not w7372 and not w7373;
w7375 <= not w7371 and w7374;
w7376 <= w257 and w5698;
w7377 <= w7375 and not w7376;
w7378 <= a(8) and not w7377;
w7379 <= a(8) and not w7378;
w7380 <= not w7377 and not w7378;
w7381 <= not w7379 and not w7380;
w7382 <= w7370 and not w7381;
w7383 <= not w7370 and w7381;
w7384 <= not w7117 and not w7383;
w7385 <= not w7382 and w7384;
w7386 <= not w7117 and not w7385;
w7387 <= not w7382 and not w7385;
w7388 <= not w7383 and w7387;
w7389 <= not w7386 and not w7388;
w7390 <= b(43) and w105;
w7391 <= b(41) and w146;
w7392 <= b(42) and w100;
w7393 <= not w7391 and not w7392;
w7394 <= not w7390 and w7393;
w7395 <= w108 and w6258;
w7396 <= w7394 and not w7395;
w7397 <= a(5) and not w7396;
w7398 <= a(5) and not w7397;
w7399 <= not w7396 and not w7397;
w7400 <= not w7398 and not w7399;
w7401 <= not w7389 and not w7400;
w7402 <= not w7389 and not w7401;
w7403 <= not w7400 and not w7401;
w7404 <= not w7402 and not w7403;
w7405 <= not w7085 and not w7091;
w7406 <= w7404 and w7405;
w7407 <= not w7404 and not w7405;
w7408 <= not w7406 and not w7407;
w7409 <= b(46) and w9;
w7410 <= b(44) and w27;
w7411 <= b(45) and w4;
w7412 <= not w7410 and not w7411;
w7413 <= not w7409 and w7412;
w7414 <= not w7100 and not w7102;
w7415 <= not b(45) and not b(46);
w7416 <= b(45) and b(46);
w7417 <= not w7415 and not w7416;
w7418 <= not w7414 and w7417;
w7419 <= w7414 and not w7417;
w7420 <= not w7418 and not w7419;
w7421 <= w12 and w7420;
w7422 <= w7413 and not w7421;
w7423 <= a(2) and not w7422;
w7424 <= a(2) and not w7423;
w7425 <= not w7422 and not w7423;
w7426 <= not w7424 and not w7425;
w7427 <= w7408 and not w7426;
w7428 <= w7408 and not w7427;
w7429 <= not w7426 and not w7427;
w7430 <= not w7428 and not w7429;
w7431 <= not w7112 and not w7114;
w7432 <= not w7430 and not w7431;
w7433 <= w7430 and w7431;
w7434 <= not w7432 and not w7433;
w7435 <= b(47) and w9;
w7436 <= b(45) and w27;
w7437 <= b(46) and w4;
w7438 <= not w7436 and not w7437;
w7439 <= not w7435 and w7438;
w7440 <= not w7416 and not w7418;
w7441 <= not b(46) and not b(47);
w7442 <= b(46) and b(47);
w7443 <= not w7441 and not w7442;
w7444 <= not w7440 and w7443;
w7445 <= w7440 and not w7443;
w7446 <= not w7444 and not w7445;
w7447 <= w12 and w7446;
w7448 <= w7439 and not w7447;
w7449 <= a(2) and not w7448;
w7450 <= a(2) and not w7449;
w7451 <= not w7448 and not w7449;
w7452 <= not w7450 and not w7451;
w7453 <= not w7401 and not w7407;
w7454 <= b(35) and w694;
w7455 <= b(33) and w799;
w7456 <= b(34) and w689;
w7457 <= not w7455 and not w7456;
w7458 <= not w7454 and w7457;
w7459 <= w697 and w4439;
w7460 <= w7458 and not w7459;
w7461 <= a(14) and not w7460;
w7462 <= a(14) and not w7461;
w7463 <= not w7460 and not w7461;
w7464 <= not w7462 and not w7463;
w7465 <= not w7338 and not w7340;
w7466 <= b(32) and w1045;
w7467 <= b(30) and w1134;
w7468 <= b(31) and w1040;
w7469 <= not w7467 and not w7468;
w7470 <= not w7466 and w7469;
w7471 <= w1048 and w3756;
w7472 <= w7470 and not w7471;
w7473 <= a(17) and not w7472;
w7474 <= a(17) and not w7473;
w7475 <= not w7472 and not w7473;
w7476 <= not w7474 and not w7475;
w7477 <= not w7318 and not w7322;
w7478 <= b(29) and w1370;
w7479 <= b(27) and w1506;
w7480 <= b(28) and w1365;
w7481 <= not w7479 and not w7480;
w7482 <= not w7478 and w7481;
w7483 <= w1373 and w3126;
w7484 <= w7482 and not w7483;
w7485 <= a(20) and not w7484;
w7486 <= a(20) and not w7485;
w7487 <= not w7484 and not w7485;
w7488 <= not w7486 and not w7487;
w7489 <= not w7310 and not w7315;
w7490 <= not w7291 and not w7297;
w7491 <= not w7252 and not w7259;
w7492 <= b(17) and w3381;
w7493 <= b(15) and w3586;
w7494 <= b(16) and w3376;
w7495 <= not w7493 and not w7494;
w7496 <= not w7492 and w7495;
w7497 <= w1099 and w3384;
w7498 <= w7496 and not w7497;
w7499 <= a(32) and not w7498;
w7500 <= a(32) and not w7499;
w7501 <= not w7498 and not w7499;
w7502 <= not w7500 and not w7501;
w7503 <= not w7247 and not w7249;
w7504 <= b(14) and w4030;
w7505 <= b(12) and w4275;
w7506 <= b(13) and w4025;
w7507 <= not w7505 and not w7506;
w7508 <= not w7504 and w7507;
w7509 <= w777 and w4033;
w7510 <= w7508 and not w7509;
w7511 <= a(35) and not w7510;
w7512 <= a(35) and not w7511;
w7513 <= not w7510 and not w7511;
w7514 <= not w7512 and not w7513;
w7515 <= not w7208 and not w7214;
w7516 <= b(8) and w5520;
w7517 <= b(6) and w5802;
w7518 <= b(7) and w5515;
w7519 <= not w7517 and not w7518;
w7520 <= not w7516 and w7519;
w7521 <= w328 and w5523;
w7522 <= w7520 and not w7521;
w7523 <= a(41) and not w7522;
w7524 <= a(41) and not w7523;
w7525 <= not w7522 and not w7523;
w7526 <= not w7524 and not w7525;
w7527 <= not w7203 and not w7205;
w7528 <= b(2) and w7189;
w7529 <= w6895 and not w7188;
w7530 <= w7183 and w7529;
w7531 <= b(0) and w7530;
w7532 <= b(1) and w7184;
w7533 <= not w7531 and not w7532;
w7534 <= not w7528 and w7533;
w7535 <= w39 and w7192;
w7536 <= w7534 and not w7535;
w7537 <= a(47) and not w7536;
w7538 <= a(47) and not w7537;
w7539 <= not w7536 and not w7537;
w7540 <= not w7538 and not w7539;
w7541 <= not w7199 and w7540;
w7542 <= w7199 and not w7540;
w7543 <= not w7541 and not w7542;
w7544 <= b(5) and w6338;
w7545 <= b(3) and w6645;
w7546 <= b(4) and w6333;
w7547 <= not w7545 and not w7546;
w7548 <= not w7544 and w7547;
w7549 <= w137 and w6341;
w7550 <= w7548 and not w7549;
w7551 <= a(44) and not w7550;
w7552 <= a(44) and not w7551;
w7553 <= not w7550 and not w7551;
w7554 <= not w7552 and not w7553;
w7555 <= w7543 and not w7554;
w7556 <= w7543 and not w7555;
w7557 <= not w7554 and not w7555;
w7558 <= not w7556 and not w7557;
w7559 <= not w7527 and not w7558;
w7560 <= w7527 and w7558;
w7561 <= not w7559 and not w7560;
w7562 <= not w7526 and w7561;
w7563 <= not w7526 and not w7562;
w7564 <= w7561 and not w7562;
w7565 <= not w7563 and not w7564;
w7566 <= not w7515 and not w7565;
w7567 <= not w7515 and not w7566;
w7568 <= not w7565 and not w7566;
w7569 <= not w7567 and not w7568;
w7570 <= b(11) and w4778;
w7571 <= b(9) and w5020;
w7572 <= b(10) and w4773;
w7573 <= not w7571 and not w7572;
w7574 <= not w7570 and w7573;
w7575 <= w561 and w4781;
w7576 <= w7574 and not w7575;
w7577 <= a(38) and not w7576;
w7578 <= a(38) and not w7577;
w7579 <= not w7576 and not w7577;
w7580 <= not w7578 and not w7579;
w7581 <= w7569 and w7580;
w7582 <= not w7569 and not w7580;
w7583 <= not w7581 and not w7582;
w7584 <= not w7232 and w7583;
w7585 <= w7232 and not w7583;
w7586 <= not w7584 and not w7585;
w7587 <= not w7514 and w7586;
w7588 <= w7586 and not w7587;
w7589 <= not w7514 and not w7587;
w7590 <= not w7588 and not w7589;
w7591 <= not w7503 and not w7590;
w7592 <= w7503 and w7590;
w7593 <= not w7591 and not w7592;
w7594 <= not w7502 and w7593;
w7595 <= not w7502 and not w7594;
w7596 <= w7593 and not w7594;
w7597 <= not w7595 and not w7596;
w7598 <= not w7491 and not w7597;
w7599 <= not w7491 and not w7598;
w7600 <= not w7597 and not w7598;
w7601 <= not w7599 and not w7600;
w7602 <= b(20) and w2793;
w7603 <= b(18) and w2986;
w7604 <= b(19) and w2788;
w7605 <= not w7603 and not w7604;
w7606 <= not w7602 and w7605;
w7607 <= w1589 and w2796;
w7608 <= w7606 and not w7607;
w7609 <= a(29) and not w7608;
w7610 <= a(29) and not w7609;
w7611 <= not w7608 and not w7609;
w7612 <= not w7610 and not w7611;
w7613 <= not w7601 and not w7612;
w7614 <= not w7601 and not w7613;
w7615 <= not w7612 and not w7613;
w7616 <= not w7614 and not w7615;
w7617 <= not w7272 and not w7278;
w7618 <= w7616 and w7617;
w7619 <= not w7616 and not w7617;
w7620 <= not w7618 and not w7619;
w7621 <= b(23) and w2282;
w7622 <= b(21) and w2428;
w7623 <= b(22) and w2277;
w7624 <= not w7622 and not w7623;
w7625 <= not w7621 and w7624;
w7626 <= w2043 and w2285;
w7627 <= w7625 and not w7626;
w7628 <= a(26) and not w7627;
w7629 <= a(26) and not w7628;
w7630 <= not w7627 and not w7628;
w7631 <= not w7629 and not w7630;
w7632 <= w7620 and not w7631;
w7633 <= not w7620 and w7631;
w7634 <= not w7490 and not w7633;
w7635 <= not w7632 and w7634;
w7636 <= not w7490 and not w7635;
w7637 <= not w7632 and not w7635;
w7638 <= not w7633 and w7637;
w7639 <= not w7636 and not w7638;
w7640 <= b(26) and w1791;
w7641 <= b(24) and w1941;
w7642 <= b(25) and w1786;
w7643 <= not w7641 and not w7642;
w7644 <= not w7640 and w7643;
w7645 <= w1794 and w2556;
w7646 <= w7644 and not w7645;
w7647 <= a(23) and not w7646;
w7648 <= a(23) and not w7647;
w7649 <= not w7646 and not w7647;
w7650 <= not w7648 and not w7649;
w7651 <= w7639 and w7650;
w7652 <= not w7639 and not w7650;
w7653 <= not w7651 and not w7652;
w7654 <= not w7489 and w7653;
w7655 <= w7489 and not w7653;
w7656 <= not w7654 and not w7655;
w7657 <= w7488 and not w7656;
w7658 <= not w7488 and w7656;
w7659 <= not w7657 and not w7658;
w7660 <= not w7477 and w7659;
w7661 <= w7477 and not w7659;
w7662 <= not w7660 and not w7661;
w7663 <= w7476 and not w7662;
w7664 <= not w7476 and w7662;
w7665 <= not w7663 and not w7664;
w7666 <= not w7465 and w7665;
w7667 <= w7465 and not w7665;
w7668 <= not w7666 and not w7667;
w7669 <= not w7464 and w7668;
w7670 <= w7668 and not w7669;
w7671 <= not w7464 and not w7669;
w7672 <= not w7670 and not w7671;
w7673 <= not w7343 and not w7350;
w7674 <= w7672 and w7673;
w7675 <= not w7672 and not w7673;
w7676 <= not w7674 and not w7675;
w7677 <= b(38) and w443;
w7678 <= b(36) and w510;
w7679 <= b(37) and w438;
w7680 <= not w7678 and not w7679;
w7681 <= not w7677 and w7680;
w7682 <= w446 and w4948;
w7683 <= w7681 and not w7682;
w7684 <= a(11) and not w7683;
w7685 <= a(11) and not w7684;
w7686 <= not w7683 and not w7684;
w7687 <= not w7685 and not w7686;
w7688 <= w7676 and not w7687;
w7689 <= w7676 and not w7688;
w7690 <= not w7687 and not w7688;
w7691 <= not w7689 and not w7690;
w7692 <= not w7363 and not w7369;
w7693 <= w7691 and w7692;
w7694 <= not w7691 and not w7692;
w7695 <= not w7693 and not w7694;
w7696 <= b(41) and w254;
w7697 <= b(39) and w284;
w7698 <= b(40) and w249;
w7699 <= not w7697 and not w7698;
w7700 <= not w7696 and w7699;
w7701 <= w257 and w5962;
w7702 <= w7700 and not w7701;
w7703 <= a(8) and not w7702;
w7704 <= a(8) and not w7703;
w7705 <= not w7702 and not w7703;
w7706 <= not w7704 and not w7705;
w7707 <= w7695 and not w7706;
w7708 <= not w7695 and w7706;
w7709 <= not w7387 and not w7708;
w7710 <= not w7707 and w7709;
w7711 <= not w7387 and not w7710;
w7712 <= not w7707 and not w7710;
w7713 <= not w7708 and w7712;
w7714 <= not w7711 and not w7713;
w7715 <= b(44) and w105;
w7716 <= b(42) and w146;
w7717 <= b(43) and w100;
w7718 <= not w7716 and not w7717;
w7719 <= not w7715 and w7718;
w7720 <= w108 and w6815;
w7721 <= w7719 and not w7720;
w7722 <= a(5) and not w7721;
w7723 <= a(5) and not w7722;
w7724 <= not w7721 and not w7722;
w7725 <= not w7723 and not w7724;
w7726 <= w7714 and w7725;
w7727 <= not w7714 and not w7725;
w7728 <= not w7726 and not w7727;
w7729 <= not w7453 and w7728;
w7730 <= w7453 and not w7728;
w7731 <= not w7729 and not w7730;
w7732 <= not w7452 and w7731;
w7733 <= w7731 and not w7732;
w7734 <= not w7452 and not w7732;
w7735 <= not w7733 and not w7734;
w7736 <= not w7427 and not w7432;
w7737 <= not w7735 and not w7736;
w7738 <= w7735 and w7736;
w7739 <= not w7737 and not w7738;
w7740 <= not w7732 and not w7737;
w7741 <= b(48) and w9;
w7742 <= b(46) and w27;
w7743 <= b(47) and w4;
w7744 <= not w7742 and not w7743;
w7745 <= not w7741 and w7744;
w7746 <= not w7442 and not w7444;
w7747 <= not b(47) and not b(48);
w7748 <= b(47) and b(48);
w7749 <= not w7747 and not w7748;
w7750 <= not w7746 and w7749;
w7751 <= w7746 and not w7749;
w7752 <= not w7750 and not w7751;
w7753 <= w12 and w7752;
w7754 <= w7745 and not w7753;
w7755 <= a(2) and not w7754;
w7756 <= a(2) and not w7755;
w7757 <= not w7754 and not w7755;
w7758 <= not w7756 and not w7757;
w7759 <= not w7727 and not w7729;
w7760 <= not w7669 and not w7675;
w7761 <= not w7664 and not w7666;
w7762 <= b(33) and w1045;
w7763 <= b(31) and w1134;
w7764 <= b(32) and w1040;
w7765 <= not w7763 and not w7764;
w7766 <= not w7762 and w7765;
w7767 <= w1048 and w3966;
w7768 <= w7766 and not w7767;
w7769 <= a(17) and not w7768;
w7770 <= a(17) and not w7769;
w7771 <= not w7768 and not w7769;
w7772 <= not w7770 and not w7771;
w7773 <= not w7658 and not w7660;
w7774 <= not w7652 and not w7654;
w7775 <= b(27) and w1791;
w7776 <= b(25) and w1941;
w7777 <= b(26) and w1786;
w7778 <= not w7776 and not w7777;
w7779 <= not w7775 and w7778;
w7780 <= w1794 and w2733;
w7781 <= w7779 and not w7780;
w7782 <= a(23) and not w7781;
w7783 <= a(23) and not w7782;
w7784 <= not w7781 and not w7782;
w7785 <= not w7783 and not w7784;
w7786 <= not w7587 and not w7591;
w7787 <= b(15) and w4030;
w7788 <= b(13) and w4275;
w7789 <= b(14) and w4025;
w7790 <= not w7788 and not w7789;
w7791 <= not w7787 and w7790;
w7792 <= w874 and w4033;
w7793 <= w7791 and not w7792;
w7794 <= a(35) and not w7793;
w7795 <= a(35) and not w7794;
w7796 <= not w7793 and not w7794;
w7797 <= not w7795 and not w7796;
w7798 <= not w7582 and not w7584;
w7799 <= b(12) and w4778;
w7800 <= b(10) and w5020;
w7801 <= b(11) and w4773;
w7802 <= not w7800 and not w7801;
w7803 <= not w7799 and w7802;
w7804 <= w585 and w4781;
w7805 <= w7803 and not w7804;
w7806 <= a(38) and not w7805;
w7807 <= a(38) and not w7806;
w7808 <= not w7805 and not w7806;
w7809 <= not w7807 and not w7808;
w7810 <= not w7562 and not w7566;
w7811 <= b(6) and w6338;
w7812 <= b(4) and w6645;
w7813 <= b(5) and w6333;
w7814 <= not w7812 and not w7813;
w7815 <= not w7811 and w7814;
w7816 <= w202 and w6341;
w7817 <= w7815 and not w7816;
w7818 <= a(44) and not w7817;
w7819 <= a(44) and not w7818;
w7820 <= not w7817 and not w7818;
w7821 <= not w7819 and not w7820;
w7822 <= a(47) and not a(48);
w7823 <= not a(47) and a(48);
w7824 <= not w7822 and not w7823;
w7825 <= b(0) and not w7824;
w7826 <= not w7542 and w7825;
w7827 <= w7542 and not w7825;
w7828 <= not w7826 and not w7827;
w7829 <= b(3) and w7189;
w7830 <= b(1) and w7530;
w7831 <= b(2) and w7184;
w7832 <= not w7830 and not w7831;
w7833 <= not w7829 and w7832;
w7834 <= w61 and w7192;
w7835 <= w7833 and not w7834;
w7836 <= a(47) and not w7835;
w7837 <= a(47) and not w7836;
w7838 <= not w7835 and not w7836;
w7839 <= not w7837 and not w7838;
w7840 <= not w7828 and not w7839;
w7841 <= w7828 and w7839;
w7842 <= not w7840 and not w7841;
w7843 <= not w7821 and w7842;
w7844 <= w7842 and not w7843;
w7845 <= not w7821 and not w7843;
w7846 <= not w7844 and not w7845;
w7847 <= not w7555 and not w7559;
w7848 <= w7846 and w7847;
w7849 <= not w7846 and not w7847;
w7850 <= not w7848 and not w7849;
w7851 <= b(9) and w5520;
w7852 <= b(7) and w5802;
w7853 <= b(8) and w5515;
w7854 <= not w7852 and not w7853;
w7855 <= not w7851 and w7854;
w7856 <= w394 and w5523;
w7857 <= w7855 and not w7856;
w7858 <= a(41) and not w7857;
w7859 <= a(41) and not w7858;
w7860 <= not w7857 and not w7858;
w7861 <= not w7859 and not w7860;
w7862 <= not w7850 and w7861;
w7863 <= w7850 and not w7861;
w7864 <= not w7862 and not w7863;
w7865 <= not w7810 and w7864;
w7866 <= w7810 and not w7864;
w7867 <= not w7865 and not w7866;
w7868 <= not w7809 and w7867;
w7869 <= not w7809 and not w7868;
w7870 <= w7867 and not w7868;
w7871 <= not w7869 and not w7870;
w7872 <= not w7798 and not w7871;
w7873 <= w7798 and not w7870;
w7874 <= not w7869 and w7873;
w7875 <= not w7872 and not w7874;
w7876 <= not w7797 and w7875;
w7877 <= w7797 and not w7875;
w7878 <= not w7876 and not w7877;
w7879 <= not w7786 and w7878;
w7880 <= w7786 and not w7878;
w7881 <= not w7879 and not w7880;
w7882 <= b(18) and w3381;
w7883 <= b(16) and w3586;
w7884 <= b(17) and w3376;
w7885 <= not w7883 and not w7884;
w7886 <= not w7882 and w7885;
w7887 <= w1309 and w3384;
w7888 <= w7886 and not w7887;
w7889 <= a(32) and not w7888;
w7890 <= a(32) and not w7889;
w7891 <= not w7888 and not w7889;
w7892 <= not w7890 and not w7891;
w7893 <= w7881 and not w7892;
w7894 <= w7881 and not w7893;
w7895 <= not w7892 and not w7893;
w7896 <= not w7894 and not w7895;
w7897 <= not w7594 and not w7598;
w7898 <= w7896 and w7897;
w7899 <= not w7896 and not w7897;
w7900 <= not w7898 and not w7899;
w7901 <= b(21) and w2793;
w7902 <= b(19) and w2986;
w7903 <= b(20) and w2788;
w7904 <= not w7902 and not w7903;
w7905 <= not w7901 and w7904;
w7906 <= w1727 and w2796;
w7907 <= w7905 and not w7906;
w7908 <= a(29) and not w7907;
w7909 <= a(29) and not w7908;
w7910 <= not w7907 and not w7908;
w7911 <= not w7909 and not w7910;
w7912 <= w7900 and not w7911;
w7913 <= w7900 and not w7912;
w7914 <= not w7911 and not w7912;
w7915 <= not w7913 and not w7914;
w7916 <= not w7613 and not w7619;
w7917 <= w7915 and w7916;
w7918 <= not w7915 and not w7916;
w7919 <= not w7917 and not w7918;
w7920 <= b(24) and w2282;
w7921 <= b(22) and w2428;
w7922 <= b(23) and w2277;
w7923 <= not w7921 and not w7922;
w7924 <= not w7920 and w7923;
w7925 <= w2201 and w2285;
w7926 <= w7924 and not w7925;
w7927 <= a(26) and not w7926;
w7928 <= a(26) and not w7927;
w7929 <= not w7926 and not w7927;
w7930 <= not w7928 and not w7929;
w7931 <= not w7919 and w7930;
w7932 <= w7919 and not w7930;
w7933 <= not w7931 and not w7932;
w7934 <= not w7637 and w7933;
w7935 <= w7637 and not w7933;
w7936 <= not w7934 and not w7935;
w7937 <= not w7785 and w7936;
w7938 <= w7936 and not w7937;
w7939 <= not w7785 and not w7937;
w7940 <= not w7938 and not w7939;
w7941 <= not w7774 and w7940;
w7942 <= w7774 and not w7940;
w7943 <= not w7941 and not w7942;
w7944 <= b(30) and w1370;
w7945 <= b(28) and w1506;
w7946 <= b(29) and w1365;
w7947 <= not w7945 and not w7946;
w7948 <= not w7944 and w7947;
w7949 <= w1373 and w3320;
w7950 <= w7948 and not w7949;
w7951 <= a(20) and not w7950;
w7952 <= a(20) and not w7951;
w7953 <= not w7950 and not w7951;
w7954 <= not w7952 and not w7953;
w7955 <= not w7943 and not w7954;
w7956 <= w7943 and w7954;
w7957 <= not w7955 and not w7956;
w7958 <= not w7773 and w7957;
w7959 <= w7773 and not w7957;
w7960 <= not w7958 and not w7959;
w7961 <= not w7772 and w7960;
w7962 <= w7960 and not w7961;
w7963 <= not w7772 and not w7961;
w7964 <= not w7962 and not w7963;
w7965 <= not w7761 and w7964;
w7966 <= w7761 and not w7964;
w7967 <= not w7965 and not w7966;
w7968 <= b(36) and w694;
w7969 <= b(34) and w799;
w7970 <= b(35) and w689;
w7971 <= not w7969 and not w7970;
w7972 <= not w7968 and w7971;
w7973 <= w697 and w4665;
w7974 <= w7972 and not w7973;
w7975 <= a(14) and not w7974;
w7976 <= a(14) and not w7975;
w7977 <= not w7974 and not w7975;
w7978 <= not w7976 and not w7977;
w7979 <= not w7967 and not w7978;
w7980 <= w7967 and w7978;
w7981 <= not w7979 and not w7980;
w7982 <= w7760 and not w7981;
w7983 <= not w7760 and w7981;
w7984 <= not w7982 and not w7983;
w7985 <= b(39) and w443;
w7986 <= b(37) and w510;
w7987 <= b(38) and w438;
w7988 <= not w7986 and not w7987;
w7989 <= not w7985 and w7988;
w7990 <= w446 and w5194;
w7991 <= w7989 and not w7990;
w7992 <= a(11) and not w7991;
w7993 <= a(11) and not w7992;
w7994 <= not w7991 and not w7992;
w7995 <= not w7993 and not w7994;
w7996 <= w7984 and not w7995;
w7997 <= w7984 and not w7996;
w7998 <= not w7995 and not w7996;
w7999 <= not w7997 and not w7998;
w8000 <= not w7688 and not w7694;
w8001 <= w7999 and w8000;
w8002 <= not w7999 and not w8000;
w8003 <= not w8001 and not w8002;
w8004 <= b(42) and w254;
w8005 <= b(40) and w284;
w8006 <= b(41) and w249;
w8007 <= not w8005 and not w8006;
w8008 <= not w8004 and w8007;
w8009 <= w257 and w6232;
w8010 <= w8008 and not w8009;
w8011 <= a(8) and not w8010;
w8012 <= a(8) and not w8011;
w8013 <= not w8010 and not w8011;
w8014 <= not w8012 and not w8013;
w8015 <= w8003 and not w8014;
w8016 <= w8003 and not w8015;
w8017 <= not w8014 and not w8015;
w8018 <= not w8016 and not w8017;
w8019 <= not w7712 and w8018;
w8020 <= w7712 and not w8018;
w8021 <= not w8019 and not w8020;
w8022 <= b(45) and w105;
w8023 <= b(43) and w146;
w8024 <= b(44) and w100;
w8025 <= not w8023 and not w8024;
w8026 <= not w8022 and w8025;
w8027 <= w108 and w7104;
w8028 <= w8026 and not w8027;
w8029 <= a(5) and not w8028;
w8030 <= a(5) and not w8029;
w8031 <= not w8028 and not w8029;
w8032 <= not w8030 and not w8031;
w8033 <= not w8021 and not w8032;
w8034 <= w8021 and w8032;
w8035 <= not w8033 and not w8034;
w8036 <= not w7759 and w8035;
w8037 <= w7759 and not w8035;
w8038 <= not w8036 and not w8037;
w8039 <= w7758 and not w8038;
w8040 <= not w7758 and w8038;
w8041 <= not w8039 and not w8040;
w8042 <= not w7740 and w8041;
w8043 <= w7740 and not w8041;
w8044 <= not w8042 and not w8043;
w8045 <= not w8040 and not w8042;
w8046 <= not w7774 and not w7940;
w8047 <= not w7937 and not w8046;
w8048 <= b(28) and w1791;
w8049 <= b(26) and w1941;
w8050 <= b(27) and w1786;
w8051 <= not w8049 and not w8050;
w8052 <= not w8048 and w8051;
w8053 <= w1794 and w2932;
w8054 <= w8052 and not w8053;
w8055 <= a(23) and not w8054;
w8056 <= a(23) and not w8055;
w8057 <= not w8054 and not w8055;
w8058 <= not w8056 and not w8057;
w8059 <= b(16) and w4030;
w8060 <= b(14) and w4275;
w8061 <= b(15) and w4025;
w8062 <= not w8060 and not w8061;
w8063 <= not w8059 and w8062;
w8064 <= w980 and w4033;
w8065 <= w8063 and not w8064;
w8066 <= a(35) and not w8065;
w8067 <= a(35) and not w8066;
w8068 <= not w8065 and not w8066;
w8069 <= not w8067 and not w8068;
w8070 <= not w7868 and not w7872;
w8071 <= not w7863 and not w7865;
w8072 <= b(7) and w6338;
w8073 <= b(5) and w6645;
w8074 <= b(6) and w6333;
w8075 <= not w8073 and not w8074;
w8076 <= not w8072 and w8075;
w8077 <= w227 and w6341;
w8078 <= w8076 and not w8077;
w8079 <= a(44) and not w8078;
w8080 <= a(44) and not w8079;
w8081 <= not w8078 and not w8079;
w8082 <= not w8080 and not w8081;
w8083 <= w7542 and w7825;
w8084 <= not w7840 and not w8083;
w8085 <= b(4) and w7189;
w8086 <= b(2) and w7530;
w8087 <= b(3) and w7184;
w8088 <= not w8086 and not w8087;
w8089 <= not w8085 and w8088;
w8090 <= w89 and w7192;
w8091 <= w8089 and not w8090;
w8092 <= a(47) and not w8091;
w8093 <= a(47) and not w8092;
w8094 <= not w8091 and not w8092;
w8095 <= not w8093 and not w8094;
w8096 <= a(50) and not w7825;
w8097 <= not a(48) and a(49);
w8098 <= a(48) and not a(49);
w8099 <= not w8097 and not w8098;
w8100 <= w7824 and not w8099;
w8101 <= b(0) and w8100;
w8102 <= not a(49) and a(50);
w8103 <= a(49) and not a(50);
w8104 <= not w8102 and not w8103;
w8105 <= not w7824 and w8104;
w8106 <= b(1) and w8105;
w8107 <= not w8101 and not w8106;
w8108 <= not w7824 and not w8104;
w8109 <= not w15 and w8108;
w8110 <= w8107 and not w8109;
w8111 <= a(50) and not w8110;
w8112 <= a(50) and not w8111;
w8113 <= not w8110 and not w8111;
w8114 <= not w8112 and not w8113;
w8115 <= w8096 and not w8114;
w8116 <= not w8096 and w8114;
w8117 <= not w8115 and not w8116;
w8118 <= w8095 and not w8117;
w8119 <= not w8095 and w8117;
w8120 <= not w8118 and not w8119;
w8121 <= not w8084 and w8120;
w8122 <= w8084 and not w8120;
w8123 <= not w8121 and not w8122;
w8124 <= not w8082 and w8123;
w8125 <= w8123 and not w8124;
w8126 <= not w8082 and not w8124;
w8127 <= not w8125 and not w8126;
w8128 <= not w7843 and not w7849;
w8129 <= w8127 and w8128;
w8130 <= not w8127 and not w8128;
w8131 <= not w8129 and not w8130;
w8132 <= b(10) and w5520;
w8133 <= b(8) and w5802;
w8134 <= b(9) and w5515;
w8135 <= not w8133 and not w8134;
w8136 <= not w8132 and w8135;
w8137 <= w481 and w5523;
w8138 <= w8136 and not w8137;
w8139 <= a(41) and not w8138;
w8140 <= a(41) and not w8139;
w8141 <= not w8138 and not w8139;
w8142 <= not w8140 and not w8141;
w8143 <= w8131 and not w8142;
w8144 <= not w8131 and w8142;
w8145 <= not w8071 and not w8144;
w8146 <= not w8143 and w8145;
w8147 <= not w8071 and not w8146;
w8148 <= not w8143 and not w8146;
w8149 <= not w8144 and w8148;
w8150 <= not w8147 and not w8149;
w8151 <= b(13) and w4778;
w8152 <= b(11) and w5020;
w8153 <= b(12) and w4773;
w8154 <= not w8152 and not w8153;
w8155 <= not w8151 and w8154;
w8156 <= w751 and w4781;
w8157 <= w8155 and not w8156;
w8158 <= a(38) and not w8157;
w8159 <= a(38) and not w8158;
w8160 <= not w8157 and not w8158;
w8161 <= not w8159 and not w8160;
w8162 <= w8150 and w8161;
w8163 <= not w8150 and not w8161;
w8164 <= not w8162 and not w8163;
w8165 <= not w8070 and w8164;
w8166 <= w8070 and not w8164;
w8167 <= not w8165 and not w8166;
w8168 <= not w8069 and w8167;
w8169 <= w8167 and not w8168;
w8170 <= not w8069 and not w8168;
w8171 <= not w8169 and not w8170;
w8172 <= not w7876 and not w7879;
w8173 <= w8171 and w8172;
w8174 <= not w8171 and not w8172;
w8175 <= not w8173 and not w8174;
w8176 <= b(19) and w3381;
w8177 <= b(17) and w3586;
w8178 <= b(18) and w3376;
w8179 <= not w8177 and not w8178;
w8180 <= not w8176 and w8179;
w8181 <= w1451 and w3384;
w8182 <= w8180 and not w8181;
w8183 <= a(32) and not w8182;
w8184 <= a(32) and not w8183;
w8185 <= not w8182 and not w8183;
w8186 <= not w8184 and not w8185;
w8187 <= w8175 and not w8186;
w8188 <= w8175 and not w8187;
w8189 <= not w8186 and not w8187;
w8190 <= not w8188 and not w8189;
w8191 <= not w7893 and not w7899;
w8192 <= w8190 and w8191;
w8193 <= not w8190 and not w8191;
w8194 <= not w8192 and not w8193;
w8195 <= b(22) and w2793;
w8196 <= b(20) and w2986;
w8197 <= b(21) and w2788;
w8198 <= not w8196 and not w8197;
w8199 <= not w8195 and w8198;
w8200 <= w1888 and w2796;
w8201 <= w8199 and not w8200;
w8202 <= a(29) and not w8201;
w8203 <= a(29) and not w8202;
w8204 <= not w8201 and not w8202;
w8205 <= not w8203 and not w8204;
w8206 <= w8194 and not w8205;
w8207 <= w8194 and not w8206;
w8208 <= not w8205 and not w8206;
w8209 <= not w8207 and not w8208;
w8210 <= not w7912 and not w7918;
w8211 <= w8209 and w8210;
w8212 <= not w8209 and not w8210;
w8213 <= not w8211 and not w8212;
w8214 <= b(25) and w2282;
w8215 <= b(23) and w2428;
w8216 <= b(24) and w2277;
w8217 <= not w8215 and not w8216;
w8218 <= not w8214 and w8217;
w8219 <= w2228 and w2285;
w8220 <= w8218 and not w8219;
w8221 <= a(26) and not w8220;
w8222 <= a(26) and not w8221;
w8223 <= not w8220 and not w8221;
w8224 <= not w8222 and not w8223;
w8225 <= w8213 and not w8224;
w8226 <= w8213 and not w8225;
w8227 <= not w8224 and not w8225;
w8228 <= not w8226 and not w8227;
w8229 <= not w7932 and not w7934;
w8230 <= not w8228 and not w8229;
w8231 <= w8228 and w8229;
w8232 <= not w8230 and not w8231;
w8233 <= not w8058 and w8232;
w8234 <= not w8058 and not w8233;
w8235 <= w8232 and not w8233;
w8236 <= not w8234 and not w8235;
w8237 <= not w8047 and not w8236;
w8238 <= not w8047 and not w8237;
w8239 <= not w8236 and not w8237;
w8240 <= not w8238 and not w8239;
w8241 <= b(31) and w1370;
w8242 <= b(29) and w1506;
w8243 <= b(30) and w1365;
w8244 <= not w8242 and not w8243;
w8245 <= not w8241 and w8244;
w8246 <= w1373 and w3539;
w8247 <= w8245 and not w8246;
w8248 <= a(20) and not w8247;
w8249 <= a(20) and not w8248;
w8250 <= not w8247 and not w8248;
w8251 <= not w8249 and not w8250;
w8252 <= not w8240 and not w8251;
w8253 <= not w8240 and not w8252;
w8254 <= not w8251 and not w8252;
w8255 <= not w8253 and not w8254;
w8256 <= not w7955 and not w7958;
w8257 <= w8255 and w8256;
w8258 <= not w8255 and not w8256;
w8259 <= not w8257 and not w8258;
w8260 <= b(34) and w1045;
w8261 <= b(32) and w1134;
w8262 <= b(33) and w1040;
w8263 <= not w8261 and not w8262;
w8264 <= not w8260 and w8263;
w8265 <= w1048 and w4209;
w8266 <= w8264 and not w8265;
w8267 <= a(17) and not w8266;
w8268 <= a(17) and not w8267;
w8269 <= not w8266 and not w8267;
w8270 <= not w8268 and not w8269;
w8271 <= w8259 and not w8270;
w8272 <= w8259 and not w8271;
w8273 <= not w8270 and not w8271;
w8274 <= not w8272 and not w8273;
w8275 <= not w7761 and not w7964;
w8276 <= not w7961 and not w8275;
w8277 <= w8274 and w8276;
w8278 <= not w8274 and not w8276;
w8279 <= not w8277 and not w8278;
w8280 <= b(37) and w694;
w8281 <= b(35) and w799;
w8282 <= b(36) and w689;
w8283 <= not w8281 and not w8282;
w8284 <= not w8280 and w8283;
w8285 <= w697 and w4924;
w8286 <= w8284 and not w8285;
w8287 <= a(14) and not w8286;
w8288 <= a(14) and not w8287;
w8289 <= not w8286 and not w8287;
w8290 <= not w8288 and not w8289;
w8291 <= w8279 and not w8290;
w8292 <= w8279 and not w8291;
w8293 <= not w8290 and not w8291;
w8294 <= not w8292 and not w8293;
w8295 <= not w7979 and not w7983;
w8296 <= w8294 and w8295;
w8297 <= not w8294 and not w8295;
w8298 <= not w8296 and not w8297;
w8299 <= b(40) and w443;
w8300 <= b(38) and w510;
w8301 <= b(39) and w438;
w8302 <= not w8300 and not w8301;
w8303 <= not w8299 and w8302;
w8304 <= w446 and w5698;
w8305 <= w8303 and not w8304;
w8306 <= a(11) and not w8305;
w8307 <= a(11) and not w8306;
w8308 <= not w8305 and not w8306;
w8309 <= not w8307 and not w8308;
w8310 <= w8298 and not w8309;
w8311 <= w8298 and not w8310;
w8312 <= not w8309 and not w8310;
w8313 <= not w8311 and not w8312;
w8314 <= not w7996 and not w8002;
w8315 <= w8313 and w8314;
w8316 <= not w8313 and not w8314;
w8317 <= not w8315 and not w8316;
w8318 <= b(43) and w254;
w8319 <= b(41) and w284;
w8320 <= b(42) and w249;
w8321 <= not w8319 and not w8320;
w8322 <= not w8318 and w8321;
w8323 <= w257 and w6258;
w8324 <= w8322 and not w8323;
w8325 <= a(8) and not w8324;
w8326 <= a(8) and not w8325;
w8327 <= not w8324 and not w8325;
w8328 <= not w8326 and not w8327;
w8329 <= w8317 and not w8328;
w8330 <= w8317 and not w8329;
w8331 <= not w8328 and not w8329;
w8332 <= not w8330 and not w8331;
w8333 <= not w7712 and not w8018;
w8334 <= not w8015 and not w8333;
w8335 <= w8332 and w8334;
w8336 <= not w8332 and not w8334;
w8337 <= not w8335 and not w8336;
w8338 <= b(46) and w105;
w8339 <= b(44) and w146;
w8340 <= b(45) and w100;
w8341 <= not w8339 and not w8340;
w8342 <= not w8338 and w8341;
w8343 <= w108 and w7420;
w8344 <= w8342 and not w8343;
w8345 <= a(5) and not w8344;
w8346 <= a(5) and not w8345;
w8347 <= not w8344 and not w8345;
w8348 <= not w8346 and not w8347;
w8349 <= w8337 and not w8348;
w8350 <= w8337 and not w8349;
w8351 <= not w8348 and not w8349;
w8352 <= not w8350 and not w8351;
w8353 <= not w8033 and not w8036;
w8354 <= w8352 and w8353;
w8355 <= not w8352 and not w8353;
w8356 <= not w8354 and not w8355;
w8357 <= b(49) and w9;
w8358 <= b(47) and w27;
w8359 <= b(48) and w4;
w8360 <= not w8358 and not w8359;
w8361 <= not w8357 and w8360;
w8362 <= not w7748 and not w7750;
w8363 <= not b(48) and not b(49);
w8364 <= b(48) and b(49);
w8365 <= not w8363 and not w8364;
w8366 <= not w8362 and w8365;
w8367 <= w8362 and not w8365;
w8368 <= not w8366 and not w8367;
w8369 <= w12 and w8368;
w8370 <= w8361 and not w8369;
w8371 <= a(2) and not w8370;
w8372 <= a(2) and not w8371;
w8373 <= not w8370 and not w8371;
w8374 <= not w8372 and not w8373;
w8375 <= not w8356 and w8374;
w8376 <= w8356 and not w8374;
w8377 <= not w8375 and not w8376;
w8378 <= not w8045 and w8377;
w8379 <= w8045 and not w8377;
w8380 <= not w8378 and not w8379;
w8381 <= not w8329 and not w8336;
w8382 <= b(35) and w1045;
w8383 <= b(33) and w1134;
w8384 <= b(34) and w1040;
w8385 <= not w8383 and not w8384;
w8386 <= not w8382 and w8385;
w8387 <= w1048 and w4439;
w8388 <= w8386 and not w8387;
w8389 <= a(17) and not w8388;
w8390 <= a(17) and not w8389;
w8391 <= not w8388 and not w8389;
w8392 <= not w8390 and not w8391;
w8393 <= not w8252 and not w8258;
w8394 <= b(32) and w1370;
w8395 <= b(30) and w1506;
w8396 <= b(31) and w1365;
w8397 <= not w8395 and not w8396;
w8398 <= not w8394 and w8397;
w8399 <= w1373 and w3756;
w8400 <= w8398 and not w8399;
w8401 <= a(20) and not w8400;
w8402 <= a(20) and not w8401;
w8403 <= not w8400 and not w8401;
w8404 <= not w8402 and not w8403;
w8405 <= not w8233 and not w8237;
w8406 <= b(29) and w1791;
w8407 <= b(27) and w1941;
w8408 <= b(28) and w1786;
w8409 <= not w8407 and not w8408;
w8410 <= not w8406 and w8409;
w8411 <= w1794 and w3126;
w8412 <= w8410 and not w8411;
w8413 <= a(23) and not w8412;
w8414 <= a(23) and not w8413;
w8415 <= not w8412 and not w8413;
w8416 <= not w8414 and not w8415;
w8417 <= not w8225 and not w8230;
w8418 <= not w8206 and not w8212;
w8419 <= not w8168 and not w8174;
w8420 <= b(17) and w4030;
w8421 <= b(15) and w4275;
w8422 <= b(16) and w4025;
w8423 <= not w8421 and not w8422;
w8424 <= not w8420 and w8423;
w8425 <= w1099 and w4033;
w8426 <= w8424 and not w8425;
w8427 <= a(35) and not w8426;
w8428 <= a(35) and not w8427;
w8429 <= not w8426 and not w8427;
w8430 <= not w8428 and not w8429;
w8431 <= not w8163 and not w8165;
w8432 <= b(14) and w4778;
w8433 <= b(12) and w5020;
w8434 <= b(13) and w4773;
w8435 <= not w8433 and not w8434;
w8436 <= not w8432 and w8435;
w8437 <= w777 and w4781;
w8438 <= w8436 and not w8437;
w8439 <= a(38) and not w8438;
w8440 <= a(38) and not w8439;
w8441 <= not w8438 and not w8439;
w8442 <= not w8440 and not w8441;
w8443 <= not w8124 and not w8130;
w8444 <= b(8) and w6338;
w8445 <= b(6) and w6645;
w8446 <= b(7) and w6333;
w8447 <= not w8445 and not w8446;
w8448 <= not w8444 and w8447;
w8449 <= w328 and w6341;
w8450 <= w8448 and not w8449;
w8451 <= a(44) and not w8450;
w8452 <= a(44) and not w8451;
w8453 <= not w8450 and not w8451;
w8454 <= not w8452 and not w8453;
w8455 <= not w8119 and not w8121;
w8456 <= b(2) and w8105;
w8457 <= w7824 and not w8104;
w8458 <= w8099 and w8457;
w8459 <= b(0) and w8458;
w8460 <= b(1) and w8100;
w8461 <= not w8459 and not w8460;
w8462 <= not w8456 and w8461;
w8463 <= w39 and w8108;
w8464 <= w8462 and not w8463;
w8465 <= a(50) and not w8464;
w8466 <= a(50) and not w8465;
w8467 <= not w8464 and not w8465;
w8468 <= not w8466 and not w8467;
w8469 <= not w8115 and w8468;
w8470 <= w8115 and not w8468;
w8471 <= not w8469 and not w8470;
w8472 <= b(5) and w7189;
w8473 <= b(3) and w7530;
w8474 <= b(4) and w7184;
w8475 <= not w8473 and not w8474;
w8476 <= not w8472 and w8475;
w8477 <= w137 and w7192;
w8478 <= w8476 and not w8477;
w8479 <= a(47) and not w8478;
w8480 <= a(47) and not w8479;
w8481 <= not w8478 and not w8479;
w8482 <= not w8480 and not w8481;
w8483 <= w8471 and not w8482;
w8484 <= w8471 and not w8483;
w8485 <= not w8482 and not w8483;
w8486 <= not w8484 and not w8485;
w8487 <= not w8455 and not w8486;
w8488 <= w8455 and w8486;
w8489 <= not w8487 and not w8488;
w8490 <= not w8454 and w8489;
w8491 <= not w8454 and not w8490;
w8492 <= w8489 and not w8490;
w8493 <= not w8491 and not w8492;
w8494 <= not w8443 and not w8493;
w8495 <= not w8443 and not w8494;
w8496 <= not w8493 and not w8494;
w8497 <= not w8495 and not w8496;
w8498 <= b(11) and w5520;
w8499 <= b(9) and w5802;
w8500 <= b(10) and w5515;
w8501 <= not w8499 and not w8500;
w8502 <= not w8498 and w8501;
w8503 <= w561 and w5523;
w8504 <= w8502 and not w8503;
w8505 <= a(41) and not w8504;
w8506 <= a(41) and not w8505;
w8507 <= not w8504 and not w8505;
w8508 <= not w8506 and not w8507;
w8509 <= w8497 and w8508;
w8510 <= not w8497 and not w8508;
w8511 <= not w8509 and not w8510;
w8512 <= not w8148 and w8511;
w8513 <= w8148 and not w8511;
w8514 <= not w8512 and not w8513;
w8515 <= not w8442 and w8514;
w8516 <= w8514 and not w8515;
w8517 <= not w8442 and not w8515;
w8518 <= not w8516 and not w8517;
w8519 <= not w8431 and not w8518;
w8520 <= w8431 and w8518;
w8521 <= not w8519 and not w8520;
w8522 <= not w8430 and w8521;
w8523 <= not w8430 and not w8522;
w8524 <= w8521 and not w8522;
w8525 <= not w8523 and not w8524;
w8526 <= not w8419 and not w8525;
w8527 <= not w8419 and not w8526;
w8528 <= not w8525 and not w8526;
w8529 <= not w8527 and not w8528;
w8530 <= b(20) and w3381;
w8531 <= b(18) and w3586;
w8532 <= b(19) and w3376;
w8533 <= not w8531 and not w8532;
w8534 <= not w8530 and w8533;
w8535 <= w1589 and w3384;
w8536 <= w8534 and not w8535;
w8537 <= a(32) and not w8536;
w8538 <= a(32) and not w8537;
w8539 <= not w8536 and not w8537;
w8540 <= not w8538 and not w8539;
w8541 <= not w8529 and not w8540;
w8542 <= not w8529 and not w8541;
w8543 <= not w8540 and not w8541;
w8544 <= not w8542 and not w8543;
w8545 <= not w8187 and not w8193;
w8546 <= w8544 and w8545;
w8547 <= not w8544 and not w8545;
w8548 <= not w8546 and not w8547;
w8549 <= b(23) and w2793;
w8550 <= b(21) and w2986;
w8551 <= b(22) and w2788;
w8552 <= not w8550 and not w8551;
w8553 <= not w8549 and w8552;
w8554 <= w2043 and w2796;
w8555 <= w8553 and not w8554;
w8556 <= a(29) and not w8555;
w8557 <= a(29) and not w8556;
w8558 <= not w8555 and not w8556;
w8559 <= not w8557 and not w8558;
w8560 <= w8548 and not w8559;
w8561 <= not w8548 and w8559;
w8562 <= not w8418 and not w8561;
w8563 <= not w8560 and w8562;
w8564 <= not w8418 and not w8563;
w8565 <= not w8560 and not w8563;
w8566 <= not w8561 and w8565;
w8567 <= not w8564 and not w8566;
w8568 <= b(26) and w2282;
w8569 <= b(24) and w2428;
w8570 <= b(25) and w2277;
w8571 <= not w8569 and not w8570;
w8572 <= not w8568 and w8571;
w8573 <= w2285 and w2556;
w8574 <= w8572 and not w8573;
w8575 <= a(26) and not w8574;
w8576 <= a(26) and not w8575;
w8577 <= not w8574 and not w8575;
w8578 <= not w8576 and not w8577;
w8579 <= w8567 and w8578;
w8580 <= not w8567 and not w8578;
w8581 <= not w8579 and not w8580;
w8582 <= not w8417 and w8581;
w8583 <= w8417 and not w8581;
w8584 <= not w8582 and not w8583;
w8585 <= w8416 and not w8584;
w8586 <= not w8416 and w8584;
w8587 <= not w8585 and not w8586;
w8588 <= not w8405 and w8587;
w8589 <= w8405 and not w8587;
w8590 <= not w8588 and not w8589;
w8591 <= w8404 and not w8590;
w8592 <= not w8404 and w8590;
w8593 <= not w8591 and not w8592;
w8594 <= not w8393 and w8593;
w8595 <= w8393 and not w8593;
w8596 <= not w8594 and not w8595;
w8597 <= not w8392 and w8596;
w8598 <= w8596 and not w8597;
w8599 <= not w8392 and not w8597;
w8600 <= not w8598 and not w8599;
w8601 <= not w8271 and not w8278;
w8602 <= w8600 and w8601;
w8603 <= not w8600 and not w8601;
w8604 <= not w8602 and not w8603;
w8605 <= b(38) and w694;
w8606 <= b(36) and w799;
w8607 <= b(37) and w689;
w8608 <= not w8606 and not w8607;
w8609 <= not w8605 and w8608;
w8610 <= w697 and w4948;
w8611 <= w8609 and not w8610;
w8612 <= a(14) and not w8611;
w8613 <= a(14) and not w8612;
w8614 <= not w8611 and not w8612;
w8615 <= not w8613 and not w8614;
w8616 <= w8604 and not w8615;
w8617 <= w8604 and not w8616;
w8618 <= not w8615 and not w8616;
w8619 <= not w8617 and not w8618;
w8620 <= not w8291 and not w8297;
w8621 <= w8619 and w8620;
w8622 <= not w8619 and not w8620;
w8623 <= not w8621 and not w8622;
w8624 <= b(41) and w443;
w8625 <= b(39) and w510;
w8626 <= b(40) and w438;
w8627 <= not w8625 and not w8626;
w8628 <= not w8624 and w8627;
w8629 <= w446 and w5962;
w8630 <= w8628 and not w8629;
w8631 <= a(11) and not w8630;
w8632 <= a(11) and not w8631;
w8633 <= not w8630 and not w8631;
w8634 <= not w8632 and not w8633;
w8635 <= w8623 and not w8634;
w8636 <= w8623 and not w8635;
w8637 <= not w8634 and not w8635;
w8638 <= not w8636 and not w8637;
w8639 <= not w8310 and not w8316;
w8640 <= w8638 and w8639;
w8641 <= not w8638 and not w8639;
w8642 <= not w8640 and not w8641;
w8643 <= b(44) and w254;
w8644 <= b(42) and w284;
w8645 <= b(43) and w249;
w8646 <= not w8644 and not w8645;
w8647 <= not w8643 and w8646;
w8648 <= w257 and w6815;
w8649 <= w8647 and not w8648;
w8650 <= a(8) and not w8649;
w8651 <= a(8) and not w8650;
w8652 <= not w8649 and not w8650;
w8653 <= not w8651 and not w8652;
w8654 <= w8642 and not w8653;
w8655 <= not w8642 and w8653;
w8656 <= not w8381 and not w8655;
w8657 <= not w8654 and w8656;
w8658 <= not w8381 and not w8657;
w8659 <= not w8654 and not w8657;
w8660 <= not w8655 and w8659;
w8661 <= not w8658 and not w8660;
w8662 <= b(47) and w105;
w8663 <= b(45) and w146;
w8664 <= b(46) and w100;
w8665 <= not w8663 and not w8664;
w8666 <= not w8662 and w8665;
w8667 <= w108 and w7446;
w8668 <= w8666 and not w8667;
w8669 <= a(5) and not w8668;
w8670 <= a(5) and not w8669;
w8671 <= not w8668 and not w8669;
w8672 <= not w8670 and not w8671;
w8673 <= not w8661 and not w8672;
w8674 <= not w8661 and not w8673;
w8675 <= not w8672 and not w8673;
w8676 <= not w8674 and not w8675;
w8677 <= not w8349 and not w8355;
w8678 <= w8676 and w8677;
w8679 <= not w8676 and not w8677;
w8680 <= not w8678 and not w8679;
w8681 <= b(50) and w9;
w8682 <= b(48) and w27;
w8683 <= b(49) and w4;
w8684 <= not w8682 and not w8683;
w8685 <= not w8681 and w8684;
w8686 <= not w8364 and not w8366;
w8687 <= not b(49) and not b(50);
w8688 <= b(49) and b(50);
w8689 <= not w8687 and not w8688;
w8690 <= not w8686 and w8689;
w8691 <= w8686 and not w8689;
w8692 <= not w8690 and not w8691;
w8693 <= w12 and w8692;
w8694 <= w8685 and not w8693;
w8695 <= a(2) and not w8694;
w8696 <= a(2) and not w8695;
w8697 <= not w8694 and not w8695;
w8698 <= not w8696 and not w8697;
w8699 <= w8680 and not w8698;
w8700 <= w8680 and not w8699;
w8701 <= not w8698 and not w8699;
w8702 <= not w8700 and not w8701;
w8703 <= not w8376 and not w8378;
w8704 <= not w8702 and not w8703;
w8705 <= w8702 and w8703;
w8706 <= not w8704 and not w8705;
w8707 <= not w8699 and not w8704;
w8708 <= b(51) and w9;
w8709 <= b(49) and w27;
w8710 <= b(50) and w4;
w8711 <= not w8709 and not w8710;
w8712 <= not w8708 and w8711;
w8713 <= not w8688 and not w8690;
w8714 <= not b(50) and not b(51);
w8715 <= b(50) and b(51);
w8716 <= not w8714 and not w8715;
w8717 <= not w8713 and w8716;
w8718 <= w8713 and not w8716;
w8719 <= not w8717 and not w8718;
w8720 <= w12 and w8719;
w8721 <= w8712 and not w8720;
w8722 <= a(2) and not w8721;
w8723 <= a(2) and not w8722;
w8724 <= not w8721 and not w8722;
w8725 <= not w8723 and not w8724;
w8726 <= not w8673 and not w8679;
w8727 <= b(45) and w254;
w8728 <= b(43) and w284;
w8729 <= b(44) and w249;
w8730 <= not w8728 and not w8729;
w8731 <= not w8727 and w8730;
w8732 <= w257 and w7104;
w8733 <= w8731 and not w8732;
w8734 <= a(8) and not w8733;
w8735 <= a(8) and not w8734;
w8736 <= not w8733 and not w8734;
w8737 <= not w8735 and not w8736;
w8738 <= not w8597 and not w8603;
w8739 <= not w8592 and not w8594;
w8740 <= b(33) and w1370;
w8741 <= b(31) and w1506;
w8742 <= b(32) and w1365;
w8743 <= not w8741 and not w8742;
w8744 <= not w8740 and w8743;
w8745 <= w1373 and w3966;
w8746 <= w8744 and not w8745;
w8747 <= a(20) and not w8746;
w8748 <= a(20) and not w8747;
w8749 <= not w8746 and not w8747;
w8750 <= not w8748 and not w8749;
w8751 <= not w8586 and not w8588;
w8752 <= not w8580 and not w8582;
w8753 <= b(27) and w2282;
w8754 <= b(25) and w2428;
w8755 <= b(26) and w2277;
w8756 <= not w8754 and not w8755;
w8757 <= not w8753 and w8756;
w8758 <= w2285 and w2733;
w8759 <= w8757 and not w8758;
w8760 <= a(26) and not w8759;
w8761 <= a(26) and not w8760;
w8762 <= not w8759 and not w8760;
w8763 <= not w8761 and not w8762;
w8764 <= not w8522 and not w8526;
w8765 <= b(18) and w4030;
w8766 <= b(16) and w4275;
w8767 <= b(17) and w4025;
w8768 <= not w8766 and not w8767;
w8769 <= not w8765 and w8768;
w8770 <= w1309 and w4033;
w8771 <= w8769 and not w8770;
w8772 <= a(35) and not w8771;
w8773 <= a(35) and not w8772;
w8774 <= not w8771 and not w8772;
w8775 <= not w8773 and not w8774;
w8776 <= not w8515 and not w8519;
w8777 <= b(15) and w4778;
w8778 <= b(13) and w5020;
w8779 <= b(14) and w4773;
w8780 <= not w8778 and not w8779;
w8781 <= not w8777 and w8780;
w8782 <= w874 and w4781;
w8783 <= w8781 and not w8782;
w8784 <= a(38) and not w8783;
w8785 <= a(38) and not w8784;
w8786 <= not w8783 and not w8784;
w8787 <= not w8785 and not w8786;
w8788 <= not w8510 and not w8512;
w8789 <= b(12) and w5520;
w8790 <= b(10) and w5802;
w8791 <= b(11) and w5515;
w8792 <= not w8790 and not w8791;
w8793 <= not w8789 and w8792;
w8794 <= w585 and w5523;
w8795 <= w8793 and not w8794;
w8796 <= a(41) and not w8795;
w8797 <= a(41) and not w8796;
w8798 <= not w8795 and not w8796;
w8799 <= not w8797 and not w8798;
w8800 <= not w8490 and not w8494;
w8801 <= b(6) and w7189;
w8802 <= b(4) and w7530;
w8803 <= b(5) and w7184;
w8804 <= not w8802 and not w8803;
w8805 <= not w8801 and w8804;
w8806 <= w202 and w7192;
w8807 <= w8805 and not w8806;
w8808 <= a(47) and not w8807;
w8809 <= a(47) and not w8808;
w8810 <= not w8807 and not w8808;
w8811 <= not w8809 and not w8810;
w8812 <= a(50) and not a(51);
w8813 <= not a(50) and a(51);
w8814 <= not w8812 and not w8813;
w8815 <= b(0) and not w8814;
w8816 <= not w8470 and w8815;
w8817 <= w8470 and not w8815;
w8818 <= not w8816 and not w8817;
w8819 <= b(3) and w8105;
w8820 <= b(1) and w8458;
w8821 <= b(2) and w8100;
w8822 <= not w8820 and not w8821;
w8823 <= not w8819 and w8822;
w8824 <= w61 and w8108;
w8825 <= w8823 and not w8824;
w8826 <= a(50) and not w8825;
w8827 <= a(50) and not w8826;
w8828 <= not w8825 and not w8826;
w8829 <= not w8827 and not w8828;
w8830 <= not w8818 and not w8829;
w8831 <= w8818 and w8829;
w8832 <= not w8830 and not w8831;
w8833 <= not w8811 and w8832;
w8834 <= w8832 and not w8833;
w8835 <= not w8811 and not w8833;
w8836 <= not w8834 and not w8835;
w8837 <= not w8483 and not w8487;
w8838 <= w8836 and w8837;
w8839 <= not w8836 and not w8837;
w8840 <= not w8838 and not w8839;
w8841 <= b(9) and w6338;
w8842 <= b(7) and w6645;
w8843 <= b(8) and w6333;
w8844 <= not w8842 and not w8843;
w8845 <= not w8841 and w8844;
w8846 <= w394 and w6341;
w8847 <= w8845 and not w8846;
w8848 <= a(44) and not w8847;
w8849 <= a(44) and not w8848;
w8850 <= not w8847 and not w8848;
w8851 <= not w8849 and not w8850;
w8852 <= not w8840 and w8851;
w8853 <= w8840 and not w8851;
w8854 <= not w8852 and not w8853;
w8855 <= not w8800 and w8854;
w8856 <= w8800 and not w8854;
w8857 <= not w8855 and not w8856;
w8858 <= not w8799 and w8857;
w8859 <= not w8799 and not w8858;
w8860 <= w8857 and not w8858;
w8861 <= not w8859 and not w8860;
w8862 <= not w8788 and not w8861;
w8863 <= w8788 and not w8860;
w8864 <= not w8859 and w8863;
w8865 <= not w8862 and not w8864;
w8866 <= not w8787 and w8865;
w8867 <= w8787 and not w8865;
w8868 <= not w8866 and not w8867;
w8869 <= not w8776 and w8868;
w8870 <= w8776 and not w8868;
w8871 <= not w8869 and not w8870;
w8872 <= not w8775 and w8871;
w8873 <= w8775 and not w8871;
w8874 <= not w8872 and not w8873;
w8875 <= not w8764 and w8874;
w8876 <= w8764 and not w8874;
w8877 <= not w8875 and not w8876;
w8878 <= b(21) and w3381;
w8879 <= b(19) and w3586;
w8880 <= b(20) and w3376;
w8881 <= not w8879 and not w8880;
w8882 <= not w8878 and w8881;
w8883 <= w1727 and w3384;
w8884 <= w8882 and not w8883;
w8885 <= a(32) and not w8884;
w8886 <= a(32) and not w8885;
w8887 <= not w8884 and not w8885;
w8888 <= not w8886 and not w8887;
w8889 <= w8877 and not w8888;
w8890 <= w8877 and not w8889;
w8891 <= not w8888 and not w8889;
w8892 <= not w8890 and not w8891;
w8893 <= not w8541 and not w8547;
w8894 <= w8892 and w8893;
w8895 <= not w8892 and not w8893;
w8896 <= not w8894 and not w8895;
w8897 <= b(24) and w2793;
w8898 <= b(22) and w2986;
w8899 <= b(23) and w2788;
w8900 <= not w8898 and not w8899;
w8901 <= not w8897 and w8900;
w8902 <= w2201 and w2796;
w8903 <= w8901 and not w8902;
w8904 <= a(29) and not w8903;
w8905 <= a(29) and not w8904;
w8906 <= not w8903 and not w8904;
w8907 <= not w8905 and not w8906;
w8908 <= not w8896 and w8907;
w8909 <= w8896 and not w8907;
w8910 <= not w8908 and not w8909;
w8911 <= not w8565 and w8910;
w8912 <= w8565 and not w8910;
w8913 <= not w8911 and not w8912;
w8914 <= not w8763 and w8913;
w8915 <= w8913 and not w8914;
w8916 <= not w8763 and not w8914;
w8917 <= not w8915 and not w8916;
w8918 <= not w8752 and w8917;
w8919 <= w8752 and not w8917;
w8920 <= not w8918 and not w8919;
w8921 <= b(30) and w1791;
w8922 <= b(28) and w1941;
w8923 <= b(29) and w1786;
w8924 <= not w8922 and not w8923;
w8925 <= not w8921 and w8924;
w8926 <= w1794 and w3320;
w8927 <= w8925 and not w8926;
w8928 <= a(23) and not w8927;
w8929 <= a(23) and not w8928;
w8930 <= not w8927 and not w8928;
w8931 <= not w8929 and not w8930;
w8932 <= not w8920 and not w8931;
w8933 <= w8920 and w8931;
w8934 <= not w8932 and not w8933;
w8935 <= not w8751 and w8934;
w8936 <= w8751 and not w8934;
w8937 <= not w8935 and not w8936;
w8938 <= not w8750 and w8937;
w8939 <= w8937 and not w8938;
w8940 <= not w8750 and not w8938;
w8941 <= not w8939 and not w8940;
w8942 <= not w8739 and w8941;
w8943 <= w8739 and not w8941;
w8944 <= not w8942 and not w8943;
w8945 <= b(36) and w1045;
w8946 <= b(34) and w1134;
w8947 <= b(35) and w1040;
w8948 <= not w8946 and not w8947;
w8949 <= not w8945 and w8948;
w8950 <= w1048 and w4665;
w8951 <= w8949 and not w8950;
w8952 <= a(17) and not w8951;
w8953 <= a(17) and not w8952;
w8954 <= not w8951 and not w8952;
w8955 <= not w8953 and not w8954;
w8956 <= not w8944 and not w8955;
w8957 <= w8944 and w8955;
w8958 <= not w8956 and not w8957;
w8959 <= w8738 and not w8958;
w8960 <= not w8738 and w8958;
w8961 <= not w8959 and not w8960;
w8962 <= b(39) and w694;
w8963 <= b(37) and w799;
w8964 <= b(38) and w689;
w8965 <= not w8963 and not w8964;
w8966 <= not w8962 and w8965;
w8967 <= w697 and w5194;
w8968 <= w8966 and not w8967;
w8969 <= a(14) and not w8968;
w8970 <= a(14) and not w8969;
w8971 <= not w8968 and not w8969;
w8972 <= not w8970 and not w8971;
w8973 <= w8961 and not w8972;
w8974 <= w8961 and not w8973;
w8975 <= not w8972 and not w8973;
w8976 <= not w8974 and not w8975;
w8977 <= not w8616 and not w8622;
w8978 <= w8976 and w8977;
w8979 <= not w8976 and not w8977;
w8980 <= not w8978 and not w8979;
w8981 <= b(42) and w443;
w8982 <= b(40) and w510;
w8983 <= b(41) and w438;
w8984 <= not w8982 and not w8983;
w8985 <= not w8981 and w8984;
w8986 <= w446 and w6232;
w8987 <= w8985 and not w8986;
w8988 <= a(11) and not w8987;
w8989 <= a(11) and not w8988;
w8990 <= not w8987 and not w8988;
w8991 <= not w8989 and not w8990;
w8992 <= not w8980 and w8991;
w8993 <= w8980 and not w8991;
w8994 <= not w8992 and not w8993;
w8995 <= not w8635 and not w8641;
w8996 <= w8994 and not w8995;
w8997 <= not w8994 and w8995;
w8998 <= not w8996 and not w8997;
w8999 <= not w8737 and w8998;
w9000 <= w8998 and not w8999;
w9001 <= not w8737 and not w8999;
w9002 <= not w9000 and not w9001;
w9003 <= not w8659 and w9002;
w9004 <= w8659 and not w9002;
w9005 <= not w9003 and not w9004;
w9006 <= b(48) and w105;
w9007 <= b(46) and w146;
w9008 <= b(47) and w100;
w9009 <= not w9007 and not w9008;
w9010 <= not w9006 and w9009;
w9011 <= w108 and w7752;
w9012 <= w9010 and not w9011;
w9013 <= a(5) and not w9012;
w9014 <= a(5) and not w9013;
w9015 <= not w9012 and not w9013;
w9016 <= not w9014 and not w9015;
w9017 <= w9005 and w9016;
w9018 <= not w9005 and not w9016;
w9019 <= not w9017 and not w9018;
w9020 <= not w8726 and w9019;
w9021 <= w8726 and not w9019;
w9022 <= not w9020 and not w9021;
w9023 <= not w8725 and w9022;
w9024 <= w8725 and not w9022;
w9025 <= not w9023 and not w9024;
w9026 <= not w8707 and w9025;
w9027 <= w8707 and not w9025;
w9028 <= not w9026 and not w9027;
w9029 <= not w9023 and not w9026;
w9030 <= not w9018 and not w9020;
w9031 <= not w8993 and not w8996;
w9032 <= not w8752 and not w8917;
w9033 <= not w8914 and not w9032;
w9034 <= not w8909 and not w8911;
w9035 <= not w8872 and not w8875;
w9036 <= b(16) and w4778;
w9037 <= b(14) and w5020;
w9038 <= b(15) and w4773;
w9039 <= not w9037 and not w9038;
w9040 <= not w9036 and w9039;
w9041 <= w980 and w4781;
w9042 <= w9040 and not w9041;
w9043 <= a(38) and not w9042;
w9044 <= a(38) and not w9043;
w9045 <= not w9042 and not w9043;
w9046 <= not w9044 and not w9045;
w9047 <= not w8858 and not w8862;
w9048 <= not w8853 and not w8855;
w9049 <= b(7) and w7189;
w9050 <= b(5) and w7530;
w9051 <= b(6) and w7184;
w9052 <= not w9050 and not w9051;
w9053 <= not w9049 and w9052;
w9054 <= w227 and w7192;
w9055 <= w9053 and not w9054;
w9056 <= a(47) and not w9055;
w9057 <= a(47) and not w9056;
w9058 <= not w9055 and not w9056;
w9059 <= not w9057 and not w9058;
w9060 <= w8470 and w8815;
w9061 <= not w8830 and not w9060;
w9062 <= b(4) and w8105;
w9063 <= b(2) and w8458;
w9064 <= b(3) and w8100;
w9065 <= not w9063 and not w9064;
w9066 <= not w9062 and w9065;
w9067 <= w89 and w8108;
w9068 <= w9066 and not w9067;
w9069 <= a(50) and not w9068;
w9070 <= a(50) and not w9069;
w9071 <= not w9068 and not w9069;
w9072 <= not w9070 and not w9071;
w9073 <= a(53) and not w8815;
w9074 <= not a(51) and a(52);
w9075 <= a(51) and not a(52);
w9076 <= not w9074 and not w9075;
w9077 <= w8814 and not w9076;
w9078 <= b(0) and w9077;
w9079 <= not a(52) and a(53);
w9080 <= a(52) and not a(53);
w9081 <= not w9079 and not w9080;
w9082 <= not w8814 and w9081;
w9083 <= b(1) and w9082;
w9084 <= not w9078 and not w9083;
w9085 <= not w8814 and not w9081;
w9086 <= not w15 and w9085;
w9087 <= w9084 and not w9086;
w9088 <= a(53) and not w9087;
w9089 <= a(53) and not w9088;
w9090 <= not w9087 and not w9088;
w9091 <= not w9089 and not w9090;
w9092 <= w9073 and not w9091;
w9093 <= not w9073 and w9091;
w9094 <= not w9092 and not w9093;
w9095 <= w9072 and not w9094;
w9096 <= not w9072 and w9094;
w9097 <= not w9095 and not w9096;
w9098 <= not w9061 and w9097;
w9099 <= w9061 and not w9097;
w9100 <= not w9098 and not w9099;
w9101 <= not w9059 and w9100;
w9102 <= w9100 and not w9101;
w9103 <= not w9059 and not w9101;
w9104 <= not w9102 and not w9103;
w9105 <= not w8833 and not w8839;
w9106 <= w9104 and w9105;
w9107 <= not w9104 and not w9105;
w9108 <= not w9106 and not w9107;
w9109 <= b(10) and w6338;
w9110 <= b(8) and w6645;
w9111 <= b(9) and w6333;
w9112 <= not w9110 and not w9111;
w9113 <= not w9109 and w9112;
w9114 <= w481 and w6341;
w9115 <= w9113 and not w9114;
w9116 <= a(44) and not w9115;
w9117 <= a(44) and not w9116;
w9118 <= not w9115 and not w9116;
w9119 <= not w9117 and not w9118;
w9120 <= w9108 and not w9119;
w9121 <= not w9108 and w9119;
w9122 <= not w9048 and not w9121;
w9123 <= not w9120 and w9122;
w9124 <= not w9048 and not w9123;
w9125 <= not w9120 and not w9123;
w9126 <= not w9121 and w9125;
w9127 <= not w9124 and not w9126;
w9128 <= b(13) and w5520;
w9129 <= b(11) and w5802;
w9130 <= b(12) and w5515;
w9131 <= not w9129 and not w9130;
w9132 <= not w9128 and w9131;
w9133 <= w751 and w5523;
w9134 <= w9132 and not w9133;
w9135 <= a(41) and not w9134;
w9136 <= a(41) and not w9135;
w9137 <= not w9134 and not w9135;
w9138 <= not w9136 and not w9137;
w9139 <= w9127 and w9138;
w9140 <= not w9127 and not w9138;
w9141 <= not w9139 and not w9140;
w9142 <= not w9047 and w9141;
w9143 <= w9047 and not w9141;
w9144 <= not w9142 and not w9143;
w9145 <= not w9046 and w9144;
w9146 <= w9144 and not w9145;
w9147 <= not w9046 and not w9145;
w9148 <= not w9146 and not w9147;
w9149 <= not w8866 and not w8869;
w9150 <= w9148 and w9149;
w9151 <= not w9148 and not w9149;
w9152 <= not w9150 and not w9151;
w9153 <= b(19) and w4030;
w9154 <= b(17) and w4275;
w9155 <= b(18) and w4025;
w9156 <= not w9154 and not w9155;
w9157 <= not w9153 and w9156;
w9158 <= w1451 and w4033;
w9159 <= w9157 and not w9158;
w9160 <= a(35) and not w9159;
w9161 <= a(35) and not w9160;
w9162 <= not w9159 and not w9160;
w9163 <= not w9161 and not w9162;
w9164 <= w9152 and not w9163;
w9165 <= not w9152 and w9163;
w9166 <= not w9035 and not w9165;
w9167 <= not w9164 and w9166;
w9168 <= not w9035 and not w9167;
w9169 <= not w9164 and not w9167;
w9170 <= not w9165 and w9169;
w9171 <= not w9168 and not w9170;
w9172 <= b(22) and w3381;
w9173 <= b(20) and w3586;
w9174 <= b(21) and w3376;
w9175 <= not w9173 and not w9174;
w9176 <= not w9172 and w9175;
w9177 <= w1888 and w3384;
w9178 <= w9176 and not w9177;
w9179 <= a(32) and not w9178;
w9180 <= a(32) and not w9179;
w9181 <= not w9178 and not w9179;
w9182 <= not w9180 and not w9181;
w9183 <= not w9171 and not w9182;
w9184 <= not w9171 and not w9183;
w9185 <= not w9182 and not w9183;
w9186 <= not w9184 and not w9185;
w9187 <= not w8889 and not w8895;
w9188 <= w9186 and w9187;
w9189 <= not w9186 and not w9187;
w9190 <= not w9188 and not w9189;
w9191 <= b(25) and w2793;
w9192 <= b(23) and w2986;
w9193 <= b(24) and w2788;
w9194 <= not w9192 and not w9193;
w9195 <= not w9191 and w9194;
w9196 <= w2228 and w2796;
w9197 <= w9195 and not w9196;
w9198 <= a(29) and not w9197;
w9199 <= a(29) and not w9198;
w9200 <= not w9197 and not w9198;
w9201 <= not w9199 and not w9200;
w9202 <= w9190 and not w9201;
w9203 <= w9190 and not w9202;
w9204 <= not w9201 and not w9202;
w9205 <= not w9203 and not w9204;
w9206 <= not w9034 and w9205;
w9207 <= w9034 and not w9205;
w9208 <= not w9206 and not w9207;
w9209 <= b(28) and w2282;
w9210 <= b(26) and w2428;
w9211 <= b(27) and w2277;
w9212 <= not w9210 and not w9211;
w9213 <= not w9209 and w9212;
w9214 <= w2285 and w2932;
w9215 <= w9213 and not w9214;
w9216 <= a(26) and not w9215;
w9217 <= a(26) and not w9216;
w9218 <= not w9215 and not w9216;
w9219 <= not w9217 and not w9218;
w9220 <= not w9208 and not w9219;
w9221 <= w9208 and w9219;
w9222 <= not w9220 and not w9221;
w9223 <= w9033 and not w9222;
w9224 <= not w9033 and w9222;
w9225 <= not w9223 and not w9224;
w9226 <= b(31) and w1791;
w9227 <= b(29) and w1941;
w9228 <= b(30) and w1786;
w9229 <= not w9227 and not w9228;
w9230 <= not w9226 and w9229;
w9231 <= w1794 and w3539;
w9232 <= w9230 and not w9231;
w9233 <= a(23) and not w9232;
w9234 <= a(23) and not w9233;
w9235 <= not w9232 and not w9233;
w9236 <= not w9234 and not w9235;
w9237 <= w9225 and not w9236;
w9238 <= w9225 and not w9237;
w9239 <= not w9236 and not w9237;
w9240 <= not w9238 and not w9239;
w9241 <= not w8932 and not w8935;
w9242 <= w9240 and w9241;
w9243 <= not w9240 and not w9241;
w9244 <= not w9242 and not w9243;
w9245 <= b(34) and w1370;
w9246 <= b(32) and w1506;
w9247 <= b(33) and w1365;
w9248 <= not w9246 and not w9247;
w9249 <= not w9245 and w9248;
w9250 <= w1373 and w4209;
w9251 <= w9249 and not w9250;
w9252 <= a(20) and not w9251;
w9253 <= a(20) and not w9252;
w9254 <= not w9251 and not w9252;
w9255 <= not w9253 and not w9254;
w9256 <= w9244 and not w9255;
w9257 <= w9244 and not w9256;
w9258 <= not w9255 and not w9256;
w9259 <= not w9257 and not w9258;
w9260 <= not w8739 and not w8941;
w9261 <= not w8938 and not w9260;
w9262 <= w9259 and w9261;
w9263 <= not w9259 and not w9261;
w9264 <= not w9262 and not w9263;
w9265 <= b(37) and w1045;
w9266 <= b(35) and w1134;
w9267 <= b(36) and w1040;
w9268 <= not w9266 and not w9267;
w9269 <= not w9265 and w9268;
w9270 <= w1048 and w4924;
w9271 <= w9269 and not w9270;
w9272 <= a(17) and not w9271;
w9273 <= a(17) and not w9272;
w9274 <= not w9271 and not w9272;
w9275 <= not w9273 and not w9274;
w9276 <= w9264 and not w9275;
w9277 <= w9264 and not w9276;
w9278 <= not w9275 and not w9276;
w9279 <= not w9277 and not w9278;
w9280 <= not w8956 and not w8960;
w9281 <= w9279 and w9280;
w9282 <= not w9279 and not w9280;
w9283 <= not w9281 and not w9282;
w9284 <= b(40) and w694;
w9285 <= b(38) and w799;
w9286 <= b(39) and w689;
w9287 <= not w9285 and not w9286;
w9288 <= not w9284 and w9287;
w9289 <= w697 and w5698;
w9290 <= w9288 and not w9289;
w9291 <= a(14) and not w9290;
w9292 <= a(14) and not w9291;
w9293 <= not w9290 and not w9291;
w9294 <= not w9292 and not w9293;
w9295 <= w9283 and not w9294;
w9296 <= w9283 and not w9295;
w9297 <= not w9294 and not w9295;
w9298 <= not w9296 and not w9297;
w9299 <= not w8973 and not w8979;
w9300 <= w9298 and w9299;
w9301 <= not w9298 and not w9299;
w9302 <= not w9300 and not w9301;
w9303 <= b(43) and w443;
w9304 <= b(41) and w510;
w9305 <= b(42) and w438;
w9306 <= not w9304 and not w9305;
w9307 <= not w9303 and w9306;
w9308 <= w446 and w6258;
w9309 <= w9307 and not w9308;
w9310 <= a(11) and not w9309;
w9311 <= a(11) and not w9310;
w9312 <= not w9309 and not w9310;
w9313 <= not w9311 and not w9312;
w9314 <= w9302 and not w9313;
w9315 <= not w9302 and w9313;
w9316 <= not w9031 and not w9315;
w9317 <= not w9314 and w9316;
w9318 <= not w9031 and not w9317;
w9319 <= not w9314 and not w9317;
w9320 <= not w9315 and w9319;
w9321 <= not w9318 and not w9320;
w9322 <= b(46) and w254;
w9323 <= b(44) and w284;
w9324 <= b(45) and w249;
w9325 <= not w9323 and not w9324;
w9326 <= not w9322 and w9325;
w9327 <= w257 and w7420;
w9328 <= w9326 and not w9327;
w9329 <= a(8) and not w9328;
w9330 <= a(8) and not w9329;
w9331 <= not w9328 and not w9329;
w9332 <= not w9330 and not w9331;
w9333 <= not w9321 and not w9332;
w9334 <= not w9321 and not w9333;
w9335 <= not w9332 and not w9333;
w9336 <= not w9334 and not w9335;
w9337 <= not w8659 and not w9002;
w9338 <= not w8999 and not w9337;
w9339 <= w9336 and w9338;
w9340 <= not w9336 and not w9338;
w9341 <= not w9339 and not w9340;
w9342 <= b(49) and w105;
w9343 <= b(47) and w146;
w9344 <= b(48) and w100;
w9345 <= not w9343 and not w9344;
w9346 <= not w9342 and w9345;
w9347 <= w108 and w8368;
w9348 <= w9346 and not w9347;
w9349 <= a(5) and not w9348;
w9350 <= a(5) and not w9349;
w9351 <= not w9348 and not w9349;
w9352 <= not w9350 and not w9351;
w9353 <= w9341 and not w9352;
w9354 <= w9341 and not w9353;
w9355 <= not w9352 and not w9353;
w9356 <= not w9354 and not w9355;
w9357 <= not w9030 and w9356;
w9358 <= w9030 and not w9356;
w9359 <= not w9357 and not w9358;
w9360 <= b(52) and w9;
w9361 <= b(50) and w27;
w9362 <= b(51) and w4;
w9363 <= not w9361 and not w9362;
w9364 <= not w9360 and w9363;
w9365 <= not w8715 and not w8717;
w9366 <= not b(51) and not b(52);
w9367 <= b(51) and b(52);
w9368 <= not w9366 and not w9367;
w9369 <= not w9365 and w9368;
w9370 <= w9365 and not w9368;
w9371 <= not w9369 and not w9370;
w9372 <= w12 and w9371;
w9373 <= w9364 and not w9372;
w9374 <= a(2) and not w9373;
w9375 <= a(2) and not w9374;
w9376 <= not w9373 and not w9374;
w9377 <= not w9375 and not w9376;
w9378 <= not w9359 and not w9377;
w9379 <= w9359 and w9377;
w9380 <= not w9378 and not w9379;
w9381 <= not w9029 and w9380;
w9382 <= w9029 and not w9380;
w9383 <= not w9381 and not w9382;
w9384 <= not w9378 and not w9381;
w9385 <= not w9030 and not w9356;
w9386 <= not w9353 and not w9385;
w9387 <= b(35) and w1370;
w9388 <= b(33) and w1506;
w9389 <= b(34) and w1365;
w9390 <= not w9388 and not w9389;
w9391 <= not w9387 and w9390;
w9392 <= w1373 and w4439;
w9393 <= w9391 and not w9392;
w9394 <= a(20) and not w9393;
w9395 <= a(20) and not w9394;
w9396 <= not w9393 and not w9394;
w9397 <= not w9395 and not w9396;
w9398 <= not w9237 and not w9243;
w9399 <= b(32) and w1791;
w9400 <= b(30) and w1941;
w9401 <= b(31) and w1786;
w9402 <= not w9400 and not w9401;
w9403 <= not w9399 and w9402;
w9404 <= w1794 and w3756;
w9405 <= w9403 and not w9404;
w9406 <= a(23) and not w9405;
w9407 <= a(23) and not w9406;
w9408 <= not w9405 and not w9406;
w9409 <= not w9407 and not w9408;
w9410 <= not w9220 and not w9224;
w9411 <= b(29) and w2282;
w9412 <= b(27) and w2428;
w9413 <= b(28) and w2277;
w9414 <= not w9412 and not w9413;
w9415 <= not w9411 and w9414;
w9416 <= w2285 and w3126;
w9417 <= w9415 and not w9416;
w9418 <= a(26) and not w9417;
w9419 <= a(26) and not w9418;
w9420 <= not w9417 and not w9418;
w9421 <= not w9419 and not w9420;
w9422 <= not w9034 and not w9205;
w9423 <= not w9202 and not w9422;
w9424 <= not w9183 and not w9189;
w9425 <= b(23) and w3381;
w9426 <= b(21) and w3586;
w9427 <= b(22) and w3376;
w9428 <= not w9426 and not w9427;
w9429 <= not w9425 and w9428;
w9430 <= w2043 and w3384;
w9431 <= w9429 and not w9430;
w9432 <= a(32) and not w9431;
w9433 <= a(32) and not w9432;
w9434 <= not w9431 and not w9432;
w9435 <= not w9433 and not w9434;
w9436 <= not w9145 and not w9151;
w9437 <= b(17) and w4778;
w9438 <= b(15) and w5020;
w9439 <= b(16) and w4773;
w9440 <= not w9438 and not w9439;
w9441 <= not w9437 and w9440;
w9442 <= w1099 and w4781;
w9443 <= w9441 and not w9442;
w9444 <= a(38) and not w9443;
w9445 <= a(38) and not w9444;
w9446 <= not w9443 and not w9444;
w9447 <= not w9445 and not w9446;
w9448 <= not w9140 and not w9142;
w9449 <= b(14) and w5520;
w9450 <= b(12) and w5802;
w9451 <= b(13) and w5515;
w9452 <= not w9450 and not w9451;
w9453 <= not w9449 and w9452;
w9454 <= w777 and w5523;
w9455 <= w9453 and not w9454;
w9456 <= a(41) and not w9455;
w9457 <= a(41) and not w9456;
w9458 <= not w9455 and not w9456;
w9459 <= not w9457 and not w9458;
w9460 <= b(11) and w6338;
w9461 <= b(9) and w6645;
w9462 <= b(10) and w6333;
w9463 <= not w9461 and not w9462;
w9464 <= not w9460 and w9463;
w9465 <= w561 and w6341;
w9466 <= w9464 and not w9465;
w9467 <= a(44) and not w9466;
w9468 <= a(44) and not w9467;
w9469 <= not w9466 and not w9467;
w9470 <= not w9468 and not w9469;
w9471 <= not w9101 and not w9107;
w9472 <= not w9096 and not w9098;
w9473 <= b(2) and w9082;
w9474 <= w8814 and not w9081;
w9475 <= w9076 and w9474;
w9476 <= b(0) and w9475;
w9477 <= b(1) and w9077;
w9478 <= not w9476 and not w9477;
w9479 <= not w9473 and w9478;
w9480 <= w39 and w9085;
w9481 <= w9479 and not w9480;
w9482 <= a(53) and not w9481;
w9483 <= a(53) and not w9482;
w9484 <= not w9481 and not w9482;
w9485 <= not w9483 and not w9484;
w9486 <= not w9092 and w9485;
w9487 <= w9092 and not w9485;
w9488 <= not w9486 and not w9487;
w9489 <= b(5) and w8105;
w9490 <= b(3) and w8458;
w9491 <= b(4) and w8100;
w9492 <= not w9490 and not w9491;
w9493 <= not w9489 and w9492;
w9494 <= w137 and w8108;
w9495 <= w9493 and not w9494;
w9496 <= a(50) and not w9495;
w9497 <= a(50) and not w9496;
w9498 <= not w9495 and not w9496;
w9499 <= not w9497 and not w9498;
w9500 <= w9488 and not w9499;
w9501 <= not w9488 and w9499;
w9502 <= not w9472 and not w9501;
w9503 <= not w9500 and w9502;
w9504 <= not w9472 and not w9503;
w9505 <= not w9500 and not w9503;
w9506 <= not w9501 and w9505;
w9507 <= not w9504 and not w9506;
w9508 <= b(8) and w7189;
w9509 <= b(6) and w7530;
w9510 <= b(7) and w7184;
w9511 <= not w9509 and not w9510;
w9512 <= not w9508 and w9511;
w9513 <= w328 and w7192;
w9514 <= w9512 and not w9513;
w9515 <= a(47) and not w9514;
w9516 <= a(47) and not w9515;
w9517 <= not w9514 and not w9515;
w9518 <= not w9516 and not w9517;
w9519 <= w9507 and w9518;
w9520 <= not w9507 and not w9518;
w9521 <= not w9519 and not w9520;
w9522 <= not w9471 and w9521;
w9523 <= w9471 and not w9521;
w9524 <= not w9522 and not w9523;
w9525 <= w9470 and not w9524;
w9526 <= not w9470 and w9524;
w9527 <= not w9525 and not w9526;
w9528 <= not w9125 and w9527;
w9529 <= w9125 and not w9527;
w9530 <= not w9528 and not w9529;
w9531 <= not w9459 and w9530;
w9532 <= w9530 and not w9531;
w9533 <= not w9459 and not w9531;
w9534 <= not w9532 and not w9533;
w9535 <= not w9448 and not w9534;
w9536 <= w9448 and w9534;
w9537 <= not w9535 and not w9536;
w9538 <= not w9447 and w9537;
w9539 <= not w9447 and not w9538;
w9540 <= w9537 and not w9538;
w9541 <= not w9539 and not w9540;
w9542 <= not w9436 and not w9541;
w9543 <= not w9436 and not w9542;
w9544 <= not w9541 and not w9542;
w9545 <= not w9543 and not w9544;
w9546 <= b(20) and w4030;
w9547 <= b(18) and w4275;
w9548 <= b(19) and w4025;
w9549 <= not w9547 and not w9548;
w9550 <= not w9546 and w9549;
w9551 <= w1589 and w4033;
w9552 <= w9550 and not w9551;
w9553 <= a(35) and not w9552;
w9554 <= a(35) and not w9553;
w9555 <= not w9552 and not w9553;
w9556 <= not w9554 and not w9555;
w9557 <= not w9545 and not w9556;
w9558 <= not w9545 and not w9557;
w9559 <= not w9556 and not w9557;
w9560 <= not w9558 and not w9559;
w9561 <= not w9169 and not w9560;
w9562 <= w9169 and w9560;
w9563 <= not w9561 and not w9562;
w9564 <= not w9435 and w9563;
w9565 <= not w9435 and not w9564;
w9566 <= w9563 and not w9564;
w9567 <= not w9565 and not w9566;
w9568 <= not w9424 and not w9567;
w9569 <= not w9424 and not w9568;
w9570 <= not w9567 and not w9568;
w9571 <= not w9569 and not w9570;
w9572 <= b(26) and w2793;
w9573 <= b(24) and w2986;
w9574 <= b(25) and w2788;
w9575 <= not w9573 and not w9574;
w9576 <= not w9572 and w9575;
w9577 <= w2556 and w2796;
w9578 <= w9576 and not w9577;
w9579 <= a(29) and not w9578;
w9580 <= a(29) and not w9579;
w9581 <= not w9578 and not w9579;
w9582 <= not w9580 and not w9581;
w9583 <= w9571 and w9582;
w9584 <= not w9571 and not w9582;
w9585 <= not w9583 and not w9584;
w9586 <= not w9423 and w9585;
w9587 <= w9423 and not w9585;
w9588 <= not w9586 and not w9587;
w9589 <= w9421 and not w9588;
w9590 <= not w9421 and w9588;
w9591 <= not w9589 and not w9590;
w9592 <= not w9410 and w9591;
w9593 <= w9410 and not w9591;
w9594 <= not w9592 and not w9593;
w9595 <= w9409 and not w9594;
w9596 <= not w9409 and w9594;
w9597 <= not w9595 and not w9596;
w9598 <= not w9398 and w9597;
w9599 <= w9398 and not w9597;
w9600 <= not w9598 and not w9599;
w9601 <= not w9397 and w9600;
w9602 <= w9600 and not w9601;
w9603 <= not w9397 and not w9601;
w9604 <= not w9602 and not w9603;
w9605 <= not w9256 and not w9263;
w9606 <= w9604 and w9605;
w9607 <= not w9604 and not w9605;
w9608 <= not w9606 and not w9607;
w9609 <= b(38) and w1045;
w9610 <= b(36) and w1134;
w9611 <= b(37) and w1040;
w9612 <= not w9610 and not w9611;
w9613 <= not w9609 and w9612;
w9614 <= w1048 and w4948;
w9615 <= w9613 and not w9614;
w9616 <= a(17) and not w9615;
w9617 <= a(17) and not w9616;
w9618 <= not w9615 and not w9616;
w9619 <= not w9617 and not w9618;
w9620 <= w9608 and not w9619;
w9621 <= w9608 and not w9620;
w9622 <= not w9619 and not w9620;
w9623 <= not w9621 and not w9622;
w9624 <= not w9276 and not w9282;
w9625 <= w9623 and w9624;
w9626 <= not w9623 and not w9624;
w9627 <= not w9625 and not w9626;
w9628 <= b(41) and w694;
w9629 <= b(39) and w799;
w9630 <= b(40) and w689;
w9631 <= not w9629 and not w9630;
w9632 <= not w9628 and w9631;
w9633 <= w697 and w5962;
w9634 <= w9632 and not w9633;
w9635 <= a(14) and not w9634;
w9636 <= a(14) and not w9635;
w9637 <= not w9634 and not w9635;
w9638 <= not w9636 and not w9637;
w9639 <= w9627 and not w9638;
w9640 <= w9627 and not w9639;
w9641 <= not w9638 and not w9639;
w9642 <= not w9640 and not w9641;
w9643 <= not w9295 and not w9301;
w9644 <= w9642 and w9643;
w9645 <= not w9642 and not w9643;
w9646 <= not w9644 and not w9645;
w9647 <= b(44) and w443;
w9648 <= b(42) and w510;
w9649 <= b(43) and w438;
w9650 <= not w9648 and not w9649;
w9651 <= not w9647 and w9650;
w9652 <= w446 and w6815;
w9653 <= w9651 and not w9652;
w9654 <= a(11) and not w9653;
w9655 <= a(11) and not w9654;
w9656 <= not w9653 and not w9654;
w9657 <= not w9655 and not w9656;
w9658 <= w9646 and not w9657;
w9659 <= not w9646 and w9657;
w9660 <= not w9319 and not w9659;
w9661 <= not w9658 and w9660;
w9662 <= not w9319 and not w9661;
w9663 <= not w9658 and not w9661;
w9664 <= not w9659 and w9663;
w9665 <= not w9662 and not w9664;
w9666 <= b(47) and w254;
w9667 <= b(45) and w284;
w9668 <= b(46) and w249;
w9669 <= not w9667 and not w9668;
w9670 <= not w9666 and w9669;
w9671 <= w257 and w7446;
w9672 <= w9670 and not w9671;
w9673 <= a(8) and not w9672;
w9674 <= a(8) and not w9673;
w9675 <= not w9672 and not w9673;
w9676 <= not w9674 and not w9675;
w9677 <= not w9665 and not w9676;
w9678 <= not w9665 and not w9677;
w9679 <= not w9676 and not w9677;
w9680 <= not w9678 and not w9679;
w9681 <= not w9333 and not w9340;
w9682 <= w9680 and w9681;
w9683 <= not w9680 and not w9681;
w9684 <= not w9682 and not w9683;
w9685 <= b(50) and w105;
w9686 <= b(48) and w146;
w9687 <= b(49) and w100;
w9688 <= not w9686 and not w9687;
w9689 <= not w9685 and w9688;
w9690 <= w108 and w8692;
w9691 <= w9689 and not w9690;
w9692 <= a(5) and not w9691;
w9693 <= a(5) and not w9692;
w9694 <= not w9691 and not w9692;
w9695 <= not w9693 and not w9694;
w9696 <= w9684 and not w9695;
w9697 <= not w9684 and w9695;
w9698 <= not w9386 and not w9697;
w9699 <= not w9696 and w9698;
w9700 <= not w9386 and not w9699;
w9701 <= not w9696 and not w9699;
w9702 <= not w9697 and w9701;
w9703 <= not w9700 and not w9702;
w9704 <= b(53) and w9;
w9705 <= b(51) and w27;
w9706 <= b(52) and w4;
w9707 <= not w9705 and not w9706;
w9708 <= not w9704 and w9707;
w9709 <= not w9367 and not w9369;
w9710 <= not b(52) and not b(53);
w9711 <= b(52) and b(53);
w9712 <= not w9710 and not w9711;
w9713 <= not w9709 and w9712;
w9714 <= w9709 and not w9712;
w9715 <= not w9713 and not w9714;
w9716 <= w12 and w9715;
w9717 <= w9708 and not w9716;
w9718 <= a(2) and not w9717;
w9719 <= a(2) and not w9718;
w9720 <= not w9717 and not w9718;
w9721 <= not w9719 and not w9720;
w9722 <= not w9703 and w9721;
w9723 <= w9703 and not w9721;
w9724 <= not w9722 and not w9723;
w9725 <= not w9384 and not w9724;
w9726 <= w9384 and w9724;
w9727 <= not w9725 and not w9726;
w9728 <= not w9703 and not w9721;
w9729 <= not w9725 and not w9728;
w9730 <= b(54) and w9;
w9731 <= b(52) and w27;
w9732 <= b(53) and w4;
w9733 <= not w9731 and not w9732;
w9734 <= not w9730 and w9733;
w9735 <= not w9711 and not w9713;
w9736 <= not b(53) and not b(54);
w9737 <= b(53) and b(54);
w9738 <= not w9736 and not w9737;
w9739 <= not w9735 and w9738;
w9740 <= w9735 and not w9738;
w9741 <= not w9739 and not w9740;
w9742 <= w12 and w9741;
w9743 <= w9734 and not w9742;
w9744 <= a(2) and not w9743;
w9745 <= a(2) and not w9744;
w9746 <= not w9743 and not w9744;
w9747 <= not w9745 and not w9746;
w9748 <= b(45) and w443;
w9749 <= b(43) and w510;
w9750 <= b(44) and w438;
w9751 <= not w9749 and not w9750;
w9752 <= not w9748 and w9751;
w9753 <= w446 and w7104;
w9754 <= w9752 and not w9753;
w9755 <= a(11) and not w9754;
w9756 <= a(11) and not w9755;
w9757 <= not w9754 and not w9755;
w9758 <= not w9756 and not w9757;
w9759 <= not w9639 and not w9645;
w9760 <= not w9601 and not w9607;
w9761 <= not w9596 and not w9598;
w9762 <= not w9590 and not w9592;
w9763 <= b(30) and w2282;
w9764 <= b(28) and w2428;
w9765 <= b(29) and w2277;
w9766 <= not w9764 and not w9765;
w9767 <= not w9763 and w9766;
w9768 <= w2285 and w3320;
w9769 <= w9767 and not w9768;
w9770 <= a(26) and not w9769;
w9771 <= a(26) and not w9770;
w9772 <= not w9769 and not w9770;
w9773 <= not w9771 and not w9772;
w9774 <= not w9584 and not w9586;
w9775 <= b(27) and w2793;
w9776 <= b(25) and w2986;
w9777 <= b(26) and w2788;
w9778 <= not w9776 and not w9777;
w9779 <= not w9775 and w9778;
w9780 <= w2733 and w2796;
w9781 <= w9779 and not w9780;
w9782 <= a(29) and not w9781;
w9783 <= a(29) and not w9782;
w9784 <= not w9781 and not w9782;
w9785 <= not w9783 and not w9784;
w9786 <= not w9564 and not w9568;
w9787 <= b(24) and w3381;
w9788 <= b(22) and w3586;
w9789 <= b(23) and w3376;
w9790 <= not w9788 and not w9789;
w9791 <= not w9787 and w9790;
w9792 <= w2201 and w3384;
w9793 <= w9791 and not w9792;
w9794 <= a(32) and not w9793;
w9795 <= a(32) and not w9794;
w9796 <= not w9793 and not w9794;
w9797 <= not w9795 and not w9796;
w9798 <= not w9557 and not w9561;
w9799 <= b(21) and w4030;
w9800 <= b(19) and w4275;
w9801 <= b(20) and w4025;
w9802 <= not w9800 and not w9801;
w9803 <= not w9799 and w9802;
w9804 <= w1727 and w4033;
w9805 <= w9803 and not w9804;
w9806 <= a(35) and not w9805;
w9807 <= a(35) and not w9806;
w9808 <= not w9805 and not w9806;
w9809 <= not w9807 and not w9808;
w9810 <= not w9538 and not w9542;
w9811 <= b(18) and w4778;
w9812 <= b(16) and w5020;
w9813 <= b(17) and w4773;
w9814 <= not w9812 and not w9813;
w9815 <= not w9811 and w9814;
w9816 <= w1309 and w4781;
w9817 <= w9815 and not w9816;
w9818 <= a(38) and not w9817;
w9819 <= a(38) and not w9818;
w9820 <= not w9817 and not w9818;
w9821 <= not w9819 and not w9820;
w9822 <= not w9531 and not w9535;
w9823 <= b(15) and w5520;
w9824 <= b(13) and w5802;
w9825 <= b(14) and w5515;
w9826 <= not w9824 and not w9825;
w9827 <= not w9823 and w9826;
w9828 <= w874 and w5523;
w9829 <= w9827 and not w9828;
w9830 <= a(41) and not w9829;
w9831 <= a(41) and not w9830;
w9832 <= not w9829 and not w9830;
w9833 <= not w9831 and not w9832;
w9834 <= not w9526 and not w9528;
w9835 <= b(12) and w6338;
w9836 <= b(10) and w6645;
w9837 <= b(11) and w6333;
w9838 <= not w9836 and not w9837;
w9839 <= not w9835 and w9838;
w9840 <= w585 and w6341;
w9841 <= w9839 and not w9840;
w9842 <= a(44) and not w9841;
w9843 <= a(44) and not w9842;
w9844 <= not w9841 and not w9842;
w9845 <= not w9843 and not w9844;
w9846 <= not w9520 and not w9522;
w9847 <= b(9) and w7189;
w9848 <= b(7) and w7530;
w9849 <= b(8) and w7184;
w9850 <= not w9848 and not w9849;
w9851 <= not w9847 and w9850;
w9852 <= w394 and w7192;
w9853 <= w9851 and not w9852;
w9854 <= a(47) and not w9853;
w9855 <= a(47) and not w9854;
w9856 <= not w9853 and not w9854;
w9857 <= not w9855 and not w9856;
w9858 <= b(6) and w8105;
w9859 <= b(4) and w8458;
w9860 <= b(5) and w8100;
w9861 <= not w9859 and not w9860;
w9862 <= not w9858 and w9861;
w9863 <= w202 and w8108;
w9864 <= w9862 and not w9863;
w9865 <= a(50) and not w9864;
w9866 <= a(50) and not w9865;
w9867 <= not w9864 and not w9865;
w9868 <= not w9866 and not w9867;
w9869 <= a(53) and not a(54);
w9870 <= not a(53) and a(54);
w9871 <= not w9869 and not w9870;
w9872 <= b(0) and not w9871;
w9873 <= not w9487 and w9872;
w9874 <= w9487 and not w9872;
w9875 <= not w9873 and not w9874;
w9876 <= b(3) and w9082;
w9877 <= b(1) and w9475;
w9878 <= b(2) and w9077;
w9879 <= not w9877 and not w9878;
w9880 <= not w9876 and w9879;
w9881 <= w61 and w9085;
w9882 <= w9880 and not w9881;
w9883 <= a(53) and not w9882;
w9884 <= a(53) and not w9883;
w9885 <= not w9882 and not w9883;
w9886 <= not w9884 and not w9885;
w9887 <= not w9875 and not w9886;
w9888 <= w9875 and w9886;
w9889 <= not w9887 and not w9888;
w9890 <= not w9868 and w9889;
w9891 <= w9889 and not w9890;
w9892 <= not w9868 and not w9890;
w9893 <= not w9891 and not w9892;
w9894 <= not w9505 and not w9893;
w9895 <= w9505 and w9893;
w9896 <= not w9894 and not w9895;
w9897 <= not w9857 and w9896;
w9898 <= not w9857 and not w9897;
w9899 <= w9896 and not w9897;
w9900 <= not w9898 and not w9899;
w9901 <= not w9846 and not w9900;
w9902 <= w9846 and not w9899;
w9903 <= not w9898 and w9902;
w9904 <= not w9901 and not w9903;
w9905 <= not w9845 and w9904;
w9906 <= not w9845 and not w9905;
w9907 <= w9904 and not w9905;
w9908 <= not w9906 and not w9907;
w9909 <= not w9834 and not w9908;
w9910 <= w9834 and not w9907;
w9911 <= not w9906 and w9910;
w9912 <= not w9909 and not w9911;
w9913 <= not w9833 and w9912;
w9914 <= w9833 and not w9912;
w9915 <= not w9913 and not w9914;
w9916 <= not w9822 and w9915;
w9917 <= w9822 and not w9915;
w9918 <= not w9916 and not w9917;
w9919 <= not w9821 and w9918;
w9920 <= not w9821 and not w9919;
w9921 <= w9918 and not w9919;
w9922 <= not w9920 and not w9921;
w9923 <= not w9810 and not w9922;
w9924 <= w9810 and not w9921;
w9925 <= not w9920 and w9924;
w9926 <= not w9923 and not w9925;
w9927 <= not w9809 and w9926;
w9928 <= w9809 and not w9926;
w9929 <= not w9927 and not w9928;
w9930 <= not w9798 and w9929;
w9931 <= w9798 and not w9929;
w9932 <= not w9930 and not w9931;
w9933 <= not w9797 and w9932;
w9934 <= w9797 and not w9932;
w9935 <= not w9933 and not w9934;
w9936 <= not w9786 and w9935;
w9937 <= w9786 and not w9935;
w9938 <= not w9936 and not w9937;
w9939 <= not w9785 and w9938;
w9940 <= w9785 and not w9938;
w9941 <= not w9939 and not w9940;
w9942 <= not w9774 and w9941;
w9943 <= w9774 and not w9941;
w9944 <= not w9942 and not w9943;
w9945 <= not w9773 and w9944;
w9946 <= w9773 and not w9944;
w9947 <= not w9945 and not w9946;
w9948 <= not w9762 and w9947;
w9949 <= w9762 and not w9947;
w9950 <= not w9948 and not w9949;
w9951 <= b(33) and w1791;
w9952 <= b(31) and w1941;
w9953 <= b(32) and w1786;
w9954 <= not w9952 and not w9953;
w9955 <= not w9951 and w9954;
w9956 <= w1794 and w3966;
w9957 <= w9955 and not w9956;
w9958 <= a(23) and not w9957;
w9959 <= a(23) and not w9958;
w9960 <= not w9957 and not w9958;
w9961 <= not w9959 and not w9960;
w9962 <= w9950 and not w9961;
w9963 <= w9950 and not w9962;
w9964 <= not w9961 and not w9962;
w9965 <= not w9963 and not w9964;
w9966 <= not w9761 and w9965;
w9967 <= w9761 and not w9965;
w9968 <= not w9966 and not w9967;
w9969 <= b(36) and w1370;
w9970 <= b(34) and w1506;
w9971 <= b(35) and w1365;
w9972 <= not w9970 and not w9971;
w9973 <= not w9969 and w9972;
w9974 <= w1373 and w4665;
w9975 <= w9973 and not w9974;
w9976 <= a(20) and not w9975;
w9977 <= a(20) and not w9976;
w9978 <= not w9975 and not w9976;
w9979 <= not w9977 and not w9978;
w9980 <= not w9968 and not w9979;
w9981 <= w9968 and w9979;
w9982 <= not w9980 and not w9981;
w9983 <= w9760 and not w9982;
w9984 <= not w9760 and w9982;
w9985 <= not w9983 and not w9984;
w9986 <= b(39) and w1045;
w9987 <= b(37) and w1134;
w9988 <= b(38) and w1040;
w9989 <= not w9987 and not w9988;
w9990 <= not w9986 and w9989;
w9991 <= w1048 and w5194;
w9992 <= w9990 and not w9991;
w9993 <= a(17) and not w9992;
w9994 <= a(17) and not w9993;
w9995 <= not w9992 and not w9993;
w9996 <= not w9994 and not w9995;
w9997 <= w9985 and not w9996;
w9998 <= w9985 and not w9997;
w9999 <= not w9996 and not w9997;
w10000 <= not w9998 and not w9999;
w10001 <= not w9620 and not w9626;
w10002 <= w10000 and w10001;
w10003 <= not w10000 and not w10001;
w10004 <= not w10002 and not w10003;
w10005 <= b(42) and w694;
w10006 <= b(40) and w799;
w10007 <= b(41) and w689;
w10008 <= not w10006 and not w10007;
w10009 <= not w10005 and w10008;
w10010 <= w697 and w6232;
w10011 <= w10009 and not w10010;
w10012 <= a(14) and not w10011;
w10013 <= a(14) and not w10012;
w10014 <= not w10011 and not w10012;
w10015 <= not w10013 and not w10014;
w10016 <= not w10004 and w10015;
w10017 <= w10004 and not w10015;
w10018 <= not w10016 and not w10017;
w10019 <= not w9759 and w10018;
w10020 <= w9759 and not w10018;
w10021 <= not w10019 and not w10020;
w10022 <= not w9758 and w10021;
w10023 <= not w9758 and not w10022;
w10024 <= w10021 and not w10022;
w10025 <= not w10023 and not w10024;
w10026 <= not w9663 and not w10025;
w10027 <= not w9663 and not w10026;
w10028 <= not w10025 and not w10026;
w10029 <= not w10027 and not w10028;
w10030 <= b(48) and w254;
w10031 <= b(46) and w284;
w10032 <= b(47) and w249;
w10033 <= not w10031 and not w10032;
w10034 <= not w10030 and w10033;
w10035 <= w257 and w7752;
w10036 <= w10034 and not w10035;
w10037 <= a(8) and not w10036;
w10038 <= a(8) and not w10037;
w10039 <= not w10036 and not w10037;
w10040 <= not w10038 and not w10039;
w10041 <= not w10029 and not w10040;
w10042 <= not w10029 and not w10041;
w10043 <= not w10040 and not w10041;
w10044 <= not w10042 and not w10043;
w10045 <= not w9677 and not w9683;
w10046 <= w10044 and w10045;
w10047 <= not w10044 and not w10045;
w10048 <= not w10046 and not w10047;
w10049 <= b(51) and w105;
w10050 <= b(49) and w146;
w10051 <= b(50) and w100;
w10052 <= not w10050 and not w10051;
w10053 <= not w10049 and w10052;
w10054 <= w108 and w8719;
w10055 <= w10053 and not w10054;
w10056 <= a(5) and not w10055;
w10057 <= a(5) and not w10056;
w10058 <= not w10055 and not w10056;
w10059 <= not w10057 and not w10058;
w10060 <= not w10048 and w10059;
w10061 <= w10048 and not w10059;
w10062 <= not w10060 and not w10061;
w10063 <= not w9701 and w10062;
w10064 <= w9701 and not w10062;
w10065 <= not w10063 and not w10064;
w10066 <= not w9747 and w10065;
w10067 <= w9747 and not w10065;
w10068 <= not w10066 and not w10067;
w10069 <= not w9729 and w10068;
w10070 <= w9729 and not w10068;
w10071 <= not w10069 and not w10070;
w10072 <= not w10066 and not w10069;
w10073 <= not w10061 and not w10063;
w10074 <= b(52) and w105;
w10075 <= b(50) and w146;
w10076 <= b(51) and w100;
w10077 <= not w10075 and not w10076;
w10078 <= not w10074 and w10077;
w10079 <= w108 and w9371;
w10080 <= w10078 and not w10079;
w10081 <= a(5) and not w10080;
w10082 <= a(5) and not w10081;
w10083 <= not w10080 and not w10081;
w10084 <= not w10082 and not w10083;
w10085 <= not w10041 and not w10047;
w10086 <= b(49) and w254;
w10087 <= b(47) and w284;
w10088 <= b(48) and w249;
w10089 <= not w10087 and not w10088;
w10090 <= not w10086 and w10089;
w10091 <= w257 and w8368;
w10092 <= w10090 and not w10091;
w10093 <= a(8) and not w10092;
w10094 <= a(8) and not w10093;
w10095 <= not w10092 and not w10093;
w10096 <= not w10094 and not w10095;
w10097 <= not w10022 and not w10026;
w10098 <= not w10017 and not w10019;
w10099 <= not w9919 and not w9923;
w10100 <= b(16) and w5520;
w10101 <= b(14) and w5802;
w10102 <= b(15) and w5515;
w10103 <= not w10101 and not w10102;
w10104 <= not w10100 and w10103;
w10105 <= w980 and w5523;
w10106 <= w10104 and not w10105;
w10107 <= a(41) and not w10106;
w10108 <= a(41) and not w10107;
w10109 <= not w10106 and not w10107;
w10110 <= not w10108 and not w10109;
w10111 <= not w9905 and not w9909;
w10112 <= b(13) and w6338;
w10113 <= b(11) and w6645;
w10114 <= b(12) and w6333;
w10115 <= not w10113 and not w10114;
w10116 <= not w10112 and w10115;
w10117 <= w751 and w6341;
w10118 <= w10116 and not w10117;
w10119 <= a(44) and not w10118;
w10120 <= a(44) and not w10119;
w10121 <= not w10118 and not w10119;
w10122 <= not w10120 and not w10121;
w10123 <= not w9897 and not w9901;
w10124 <= b(10) and w7189;
w10125 <= b(8) and w7530;
w10126 <= b(9) and w7184;
w10127 <= not w10125 and not w10126;
w10128 <= not w10124 and w10127;
w10129 <= w481 and w7192;
w10130 <= w10128 and not w10129;
w10131 <= a(47) and not w10130;
w10132 <= a(47) and not w10131;
w10133 <= not w10130 and not w10131;
w10134 <= not w10132 and not w10133;
w10135 <= not w9890 and not w9894;
w10136 <= b(7) and w8105;
w10137 <= b(5) and w8458;
w10138 <= b(6) and w8100;
w10139 <= not w10137 and not w10138;
w10140 <= not w10136 and w10139;
w10141 <= w227 and w8108;
w10142 <= w10140 and not w10141;
w10143 <= a(50) and not w10142;
w10144 <= a(50) and not w10143;
w10145 <= not w10142 and not w10143;
w10146 <= not w10144 and not w10145;
w10147 <= w9487 and w9872;
w10148 <= not w9887 and not w10147;
w10149 <= b(4) and w9082;
w10150 <= b(2) and w9475;
w10151 <= b(3) and w9077;
w10152 <= not w10150 and not w10151;
w10153 <= not w10149 and w10152;
w10154 <= w89 and w9085;
w10155 <= w10153 and not w10154;
w10156 <= a(53) and not w10155;
w10157 <= a(53) and not w10156;
w10158 <= not w10155 and not w10156;
w10159 <= not w10157 and not w10158;
w10160 <= a(56) and not w9872;
w10161 <= not a(54) and a(55);
w10162 <= a(54) and not a(55);
w10163 <= not w10161 and not w10162;
w10164 <= w9871 and not w10163;
w10165 <= b(0) and w10164;
w10166 <= not a(55) and a(56);
w10167 <= a(55) and not a(56);
w10168 <= not w10166 and not w10167;
w10169 <= not w9871 and w10168;
w10170 <= b(1) and w10169;
w10171 <= not w10165 and not w10170;
w10172 <= not w9871 and not w10168;
w10173 <= not w15 and w10172;
w10174 <= w10171 and not w10173;
w10175 <= a(56) and not w10174;
w10176 <= a(56) and not w10175;
w10177 <= not w10174 and not w10175;
w10178 <= not w10176 and not w10177;
w10179 <= w10160 and not w10178;
w10180 <= not w10160 and w10178;
w10181 <= not w10179 and not w10180;
w10182 <= w10159 and not w10181;
w10183 <= not w10159 and w10181;
w10184 <= not w10182 and not w10183;
w10185 <= not w10148 and w10184;
w10186 <= w10148 and not w10184;
w10187 <= not w10185 and not w10186;
w10188 <= w10146 and not w10187;
w10189 <= not w10146 and w10187;
w10190 <= not w10188 and not w10189;
w10191 <= not w10135 and w10190;
w10192 <= w10135 and not w10190;
w10193 <= not w10191 and not w10192;
w10194 <= w10134 and not w10193;
w10195 <= not w10134 and w10193;
w10196 <= not w10194 and not w10195;
w10197 <= not w10123 and w10196;
w10198 <= w10123 and not w10196;
w10199 <= not w10197 and not w10198;
w10200 <= w10122 and not w10199;
w10201 <= not w10122 and w10199;
w10202 <= not w10200 and not w10201;
w10203 <= not w10111 and w10202;
w10204 <= w10111 and not w10202;
w10205 <= not w10203 and not w10204;
w10206 <= not w10110 and w10205;
w10207 <= w10205 and not w10206;
w10208 <= not w10110 and not w10206;
w10209 <= not w10207 and not w10208;
w10210 <= not w9913 and not w9916;
w10211 <= w10209 and w10210;
w10212 <= not w10209 and not w10210;
w10213 <= not w10211 and not w10212;
w10214 <= b(19) and w4778;
w10215 <= b(17) and w5020;
w10216 <= b(18) and w4773;
w10217 <= not w10215 and not w10216;
w10218 <= not w10214 and w10217;
w10219 <= w1451 and w4781;
w10220 <= w10218 and not w10219;
w10221 <= a(38) and not w10220;
w10222 <= a(38) and not w10221;
w10223 <= not w10220 and not w10221;
w10224 <= not w10222 and not w10223;
w10225 <= w10213 and not w10224;
w10226 <= not w10213 and w10224;
w10227 <= not w10099 and not w10226;
w10228 <= not w10225 and w10227;
w10229 <= not w10099 and not w10228;
w10230 <= not w10225 and not w10228;
w10231 <= not w10226 and w10230;
w10232 <= not w10229 and not w10231;
w10233 <= b(22) and w4030;
w10234 <= b(20) and w4275;
w10235 <= b(21) and w4025;
w10236 <= not w10234 and not w10235;
w10237 <= not w10233 and w10236;
w10238 <= w1888 and w4033;
w10239 <= w10237 and not w10238;
w10240 <= a(35) and not w10239;
w10241 <= a(35) and not w10240;
w10242 <= not w10239 and not w10240;
w10243 <= not w10241 and not w10242;
w10244 <= not w10232 and not w10243;
w10245 <= not w10232 and not w10244;
w10246 <= not w10243 and not w10244;
w10247 <= not w10245 and not w10246;
w10248 <= not w9927 and not w9930;
w10249 <= w10247 and w10248;
w10250 <= not w10247 and not w10248;
w10251 <= not w10249 and not w10250;
w10252 <= b(25) and w3381;
w10253 <= b(23) and w3586;
w10254 <= b(24) and w3376;
w10255 <= not w10253 and not w10254;
w10256 <= not w10252 and w10255;
w10257 <= w2228 and w3384;
w10258 <= w10256 and not w10257;
w10259 <= a(32) and not w10258;
w10260 <= a(32) and not w10259;
w10261 <= not w10258 and not w10259;
w10262 <= not w10260 and not w10261;
w10263 <= w10251 and not w10262;
w10264 <= w10251 and not w10263;
w10265 <= not w10262 and not w10263;
w10266 <= not w10264 and not w10265;
w10267 <= not w9933 and not w9936;
w10268 <= w10266 and w10267;
w10269 <= not w10266 and not w10267;
w10270 <= not w10268 and not w10269;
w10271 <= b(28) and w2793;
w10272 <= b(26) and w2986;
w10273 <= b(27) and w2788;
w10274 <= not w10272 and not w10273;
w10275 <= not w10271 and w10274;
w10276 <= w2796 and w2932;
w10277 <= w10275 and not w10276;
w10278 <= a(29) and not w10277;
w10279 <= a(29) and not w10278;
w10280 <= not w10277 and not w10278;
w10281 <= not w10279 and not w10280;
w10282 <= w10270 and not w10281;
w10283 <= w10270 and not w10282;
w10284 <= not w10281 and not w10282;
w10285 <= not w10283 and not w10284;
w10286 <= not w9939 and not w9942;
w10287 <= w10285 and w10286;
w10288 <= not w10285 and not w10286;
w10289 <= not w10287 and not w10288;
w10290 <= b(31) and w2282;
w10291 <= b(29) and w2428;
w10292 <= b(30) and w2277;
w10293 <= not w10291 and not w10292;
w10294 <= not w10290 and w10293;
w10295 <= w2285 and w3539;
w10296 <= w10294 and not w10295;
w10297 <= a(26) and not w10296;
w10298 <= a(26) and not w10297;
w10299 <= not w10296 and not w10297;
w10300 <= not w10298 and not w10299;
w10301 <= w10289 and not w10300;
w10302 <= w10289 and not w10301;
w10303 <= not w10300 and not w10301;
w10304 <= not w10302 and not w10303;
w10305 <= not w9945 and not w9948;
w10306 <= w10304 and w10305;
w10307 <= not w10304 and not w10305;
w10308 <= not w10306 and not w10307;
w10309 <= b(34) and w1791;
w10310 <= b(32) and w1941;
w10311 <= b(33) and w1786;
w10312 <= not w10310 and not w10311;
w10313 <= not w10309 and w10312;
w10314 <= w1794 and w4209;
w10315 <= w10313 and not w10314;
w10316 <= a(23) and not w10315;
w10317 <= a(23) and not w10316;
w10318 <= not w10315 and not w10316;
w10319 <= not w10317 and not w10318;
w10320 <= w10308 and not w10319;
w10321 <= w10308 and not w10320;
w10322 <= not w10319 and not w10320;
w10323 <= not w10321 and not w10322;
w10324 <= not w9761 and not w9965;
w10325 <= not w9962 and not w10324;
w10326 <= w10323 and w10325;
w10327 <= not w10323 and not w10325;
w10328 <= not w10326 and not w10327;
w10329 <= b(37) and w1370;
w10330 <= b(35) and w1506;
w10331 <= b(36) and w1365;
w10332 <= not w10330 and not w10331;
w10333 <= not w10329 and w10332;
w10334 <= w1373 and w4924;
w10335 <= w10333 and not w10334;
w10336 <= a(20) and not w10335;
w10337 <= a(20) and not w10336;
w10338 <= not w10335 and not w10336;
w10339 <= not w10337 and not w10338;
w10340 <= w10328 and not w10339;
w10341 <= w10328 and not w10340;
w10342 <= not w10339 and not w10340;
w10343 <= not w10341 and not w10342;
w10344 <= not w9980 and not w9984;
w10345 <= w10343 and w10344;
w10346 <= not w10343 and not w10344;
w10347 <= not w10345 and not w10346;
w10348 <= b(40) and w1045;
w10349 <= b(38) and w1134;
w10350 <= b(39) and w1040;
w10351 <= not w10349 and not w10350;
w10352 <= not w10348 and w10351;
w10353 <= w1048 and w5698;
w10354 <= w10352 and not w10353;
w10355 <= a(17) and not w10354;
w10356 <= a(17) and not w10355;
w10357 <= not w10354 and not w10355;
w10358 <= not w10356 and not w10357;
w10359 <= w10347 and not w10358;
w10360 <= w10347 and not w10359;
w10361 <= not w10358 and not w10359;
w10362 <= not w10360 and not w10361;
w10363 <= not w9997 and not w10003;
w10364 <= w10362 and w10363;
w10365 <= not w10362 and not w10363;
w10366 <= not w10364 and not w10365;
w10367 <= b(43) and w694;
w10368 <= b(41) and w799;
w10369 <= b(42) and w689;
w10370 <= not w10368 and not w10369;
w10371 <= not w10367 and w10370;
w10372 <= w697 and w6258;
w10373 <= w10371 and not w10372;
w10374 <= a(14) and not w10373;
w10375 <= a(14) and not w10374;
w10376 <= not w10373 and not w10374;
w10377 <= not w10375 and not w10376;
w10378 <= w10366 and not w10377;
w10379 <= not w10366 and w10377;
w10380 <= not w10098 and not w10379;
w10381 <= not w10378 and w10380;
w10382 <= not w10098 and not w10381;
w10383 <= not w10378 and not w10381;
w10384 <= not w10379 and w10383;
w10385 <= not w10382 and not w10384;
w10386 <= b(46) and w443;
w10387 <= b(44) and w510;
w10388 <= b(45) and w438;
w10389 <= not w10387 and not w10388;
w10390 <= not w10386 and w10389;
w10391 <= w446 and w7420;
w10392 <= w10390 and not w10391;
w10393 <= a(11) and not w10392;
w10394 <= a(11) and not w10393;
w10395 <= not w10392 and not w10393;
w10396 <= not w10394 and not w10395;
w10397 <= w10385 and w10396;
w10398 <= not w10385 and not w10396;
w10399 <= not w10397 and not w10398;
w10400 <= not w10097 and w10399;
w10401 <= w10097 and not w10399;
w10402 <= not w10400 and not w10401;
w10403 <= w10096 and not w10402;
w10404 <= not w10096 and w10402;
w10405 <= not w10403 and not w10404;
w10406 <= not w10085 and w10405;
w10407 <= w10085 and not w10405;
w10408 <= not w10406 and not w10407;
w10409 <= not w10084 and w10408;
w10410 <= w10408 and not w10409;
w10411 <= not w10084 and not w10409;
w10412 <= not w10410 and not w10411;
w10413 <= not w10073 and w10412;
w10414 <= w10073 and not w10412;
w10415 <= not w10413 and not w10414;
w10416 <= b(55) and w9;
w10417 <= b(53) and w27;
w10418 <= b(54) and w4;
w10419 <= not w10417 and not w10418;
w10420 <= not w10416 and w10419;
w10421 <= not w9737 and not w9739;
w10422 <= not b(54) and not b(55);
w10423 <= b(54) and b(55);
w10424 <= not w10422 and not w10423;
w10425 <= not w10421 and w10424;
w10426 <= w10421 and not w10424;
w10427 <= not w10425 and not w10426;
w10428 <= w12 and w10427;
w10429 <= w10420 and not w10428;
w10430 <= a(2) and not w10429;
w10431 <= a(2) and not w10430;
w10432 <= not w10429 and not w10430;
w10433 <= not w10431 and not w10432;
w10434 <= not w10415 and not w10433;
w10435 <= w10415 and w10433;
w10436 <= not w10434 and not w10435;
w10437 <= not w10072 and w10436;
w10438 <= w10072 and not w10436;
w10439 <= not w10437 and not w10438;
w10440 <= b(56) and w9;
w10441 <= b(54) and w27;
w10442 <= b(55) and w4;
w10443 <= not w10441 and not w10442;
w10444 <= not w10440 and w10443;
w10445 <= not w10423 and not w10425;
w10446 <= not b(55) and not b(56);
w10447 <= b(55) and b(56);
w10448 <= not w10446 and not w10447;
w10449 <= not w10445 and w10448;
w10450 <= w10445 and not w10448;
w10451 <= not w10449 and not w10450;
w10452 <= w12 and w10451;
w10453 <= w10444 and not w10452;
w10454 <= a(2) and not w10453;
w10455 <= a(2) and not w10454;
w10456 <= not w10453 and not w10454;
w10457 <= not w10455 and not w10456;
w10458 <= not w10073 and not w10412;
w10459 <= not w10409 and not w10458;
w10460 <= not w10404 and not w10406;
w10461 <= b(50) and w254;
w10462 <= b(48) and w284;
w10463 <= b(49) and w249;
w10464 <= not w10462 and not w10463;
w10465 <= not w10461 and w10464;
w10466 <= w257 and w8692;
w10467 <= w10465 and not w10466;
w10468 <= a(8) and not w10467;
w10469 <= a(8) and not w10468;
w10470 <= not w10467 and not w10468;
w10471 <= not w10469 and not w10470;
w10472 <= not w10398 and not w10400;
w10473 <= b(35) and w1791;
w10474 <= b(33) and w1941;
w10475 <= b(34) and w1786;
w10476 <= not w10474 and not w10475;
w10477 <= not w10473 and w10476;
w10478 <= w1794 and w4439;
w10479 <= w10477 and not w10478;
w10480 <= a(23) and not w10479;
w10481 <= a(23) and not w10480;
w10482 <= not w10479 and not w10480;
w10483 <= not w10481 and not w10482;
w10484 <= not w10301 and not w10307;
w10485 <= b(32) and w2282;
w10486 <= b(30) and w2428;
w10487 <= b(31) and w2277;
w10488 <= not w10486 and not w10487;
w10489 <= not w10485 and w10488;
w10490 <= w2285 and w3756;
w10491 <= w10489 and not w10490;
w10492 <= a(26) and not w10491;
w10493 <= a(26) and not w10492;
w10494 <= not w10491 and not w10492;
w10495 <= not w10493 and not w10494;
w10496 <= not w10282 and not w10288;
w10497 <= not w10263 and not w10269;
w10498 <= not w10244 and not w10250;
w10499 <= not w10206 and not w10212;
w10500 <= b(17) and w5520;
w10501 <= b(15) and w5802;
w10502 <= b(16) and w5515;
w10503 <= not w10501 and not w10502;
w10504 <= not w10500 and w10503;
w10505 <= w1099 and w5523;
w10506 <= w10504 and not w10505;
w10507 <= a(41) and not w10506;
w10508 <= a(41) and not w10507;
w10509 <= not w10506 and not w10507;
w10510 <= not w10508 and not w10509;
w10511 <= not w10201 and not w10203;
w10512 <= b(14) and w6338;
w10513 <= b(12) and w6645;
w10514 <= b(13) and w6333;
w10515 <= not w10513 and not w10514;
w10516 <= not w10512 and w10515;
w10517 <= w777 and w6341;
w10518 <= w10516 and not w10517;
w10519 <= a(44) and not w10518;
w10520 <= a(44) and not w10519;
w10521 <= not w10518 and not w10519;
w10522 <= not w10520 and not w10521;
w10523 <= not w10195 and not w10197;
w10524 <= b(11) and w7189;
w10525 <= b(9) and w7530;
w10526 <= b(10) and w7184;
w10527 <= not w10525 and not w10526;
w10528 <= not w10524 and w10527;
w10529 <= w561 and w7192;
w10530 <= w10528 and not w10529;
w10531 <= a(47) and not w10530;
w10532 <= a(47) and not w10531;
w10533 <= not w10530 and not w10531;
w10534 <= not w10532 and not w10533;
w10535 <= not w10189 and not w10191;
w10536 <= not w10183 and not w10185;
w10537 <= b(2) and w10169;
w10538 <= w9871 and not w10168;
w10539 <= w10163 and w10538;
w10540 <= b(0) and w10539;
w10541 <= b(1) and w10164;
w10542 <= not w10540 and not w10541;
w10543 <= not w10537 and w10542;
w10544 <= w39 and w10172;
w10545 <= w10543 and not w10544;
w10546 <= a(56) and not w10545;
w10547 <= a(56) and not w10546;
w10548 <= not w10545 and not w10546;
w10549 <= not w10547 and not w10548;
w10550 <= not w10179 and w10549;
w10551 <= w10179 and not w10549;
w10552 <= not w10550 and not w10551;
w10553 <= b(5) and w9082;
w10554 <= b(3) and w9475;
w10555 <= b(4) and w9077;
w10556 <= not w10554 and not w10555;
w10557 <= not w10553 and w10556;
w10558 <= w137 and w9085;
w10559 <= w10557 and not w10558;
w10560 <= a(53) and not w10559;
w10561 <= a(53) and not w10560;
w10562 <= not w10559 and not w10560;
w10563 <= not w10561 and not w10562;
w10564 <= w10552 and not w10563;
w10565 <= not w10552 and w10563;
w10566 <= not w10536 and not w10565;
w10567 <= not w10564 and w10566;
w10568 <= not w10536 and not w10567;
w10569 <= not w10564 and not w10567;
w10570 <= not w10565 and w10569;
w10571 <= not w10568 and not w10570;
w10572 <= b(8) and w8105;
w10573 <= b(6) and w8458;
w10574 <= b(7) and w8100;
w10575 <= not w10573 and not w10574;
w10576 <= not w10572 and w10575;
w10577 <= w328 and w8108;
w10578 <= w10576 and not w10577;
w10579 <= a(50) and not w10578;
w10580 <= a(50) and not w10579;
w10581 <= not w10578 and not w10579;
w10582 <= not w10580 and not w10581;
w10583 <= w10571 and w10582;
w10584 <= not w10571 and not w10582;
w10585 <= not w10583 and not w10584;
w10586 <= not w10535 and w10585;
w10587 <= w10535 and not w10585;
w10588 <= not w10586 and not w10587;
w10589 <= w10534 and not w10588;
w10590 <= not w10534 and w10588;
w10591 <= not w10589 and not w10590;
w10592 <= not w10523 and w10591;
w10593 <= w10523 and not w10591;
w10594 <= not w10592 and not w10593;
w10595 <= not w10522 and w10594;
w10596 <= w10594 and not w10595;
w10597 <= not w10522 and not w10595;
w10598 <= not w10596 and not w10597;
w10599 <= not w10511 and not w10598;
w10600 <= w10511 and w10598;
w10601 <= not w10599 and not w10600;
w10602 <= not w10510 and w10601;
w10603 <= not w10510 and not w10602;
w10604 <= w10601 and not w10602;
w10605 <= not w10603 and not w10604;
w10606 <= not w10499 and not w10605;
w10607 <= not w10499 and not w10606;
w10608 <= not w10605 and not w10606;
w10609 <= not w10607 and not w10608;
w10610 <= b(20) and w4778;
w10611 <= b(18) and w5020;
w10612 <= b(19) and w4773;
w10613 <= not w10611 and not w10612;
w10614 <= not w10610 and w10613;
w10615 <= w1589 and w4781;
w10616 <= w10614 and not w10615;
w10617 <= a(38) and not w10616;
w10618 <= a(38) and not w10617;
w10619 <= not w10616 and not w10617;
w10620 <= not w10618 and not w10619;
w10621 <= not w10609 and not w10620;
w10622 <= not w10609 and not w10621;
w10623 <= not w10620 and not w10621;
w10624 <= not w10622 and not w10623;
w10625 <= not w10230 and w10624;
w10626 <= w10230 and not w10624;
w10627 <= not w10625 and not w10626;
w10628 <= b(23) and w4030;
w10629 <= b(21) and w4275;
w10630 <= b(22) and w4025;
w10631 <= not w10629 and not w10630;
w10632 <= not w10628 and w10631;
w10633 <= w2043 and w4033;
w10634 <= w10632 and not w10633;
w10635 <= a(35) and not w10634;
w10636 <= a(35) and not w10635;
w10637 <= not w10634 and not w10635;
w10638 <= not w10636 and not w10637;
w10639 <= not w10627 and not w10638;
w10640 <= w10627 and w10638;
w10641 <= not w10639 and not w10640;
w10642 <= w10498 and not w10641;
w10643 <= not w10498 and w10641;
w10644 <= not w10642 and not w10643;
w10645 <= b(26) and w3381;
w10646 <= b(24) and w3586;
w10647 <= b(25) and w3376;
w10648 <= not w10646 and not w10647;
w10649 <= not w10645 and w10648;
w10650 <= w2556 and w3384;
w10651 <= w10649 and not w10650;
w10652 <= a(32) and not w10651;
w10653 <= a(32) and not w10652;
w10654 <= not w10651 and not w10652;
w10655 <= not w10653 and not w10654;
w10656 <= w10644 and not w10655;
w10657 <= not w10644 and w10655;
w10658 <= not w10497 and not w10657;
w10659 <= not w10656 and w10658;
w10660 <= not w10497 and not w10659;
w10661 <= not w10656 and not w10659;
w10662 <= not w10657 and w10661;
w10663 <= not w10660 and not w10662;
w10664 <= b(29) and w2793;
w10665 <= b(27) and w2986;
w10666 <= b(28) and w2788;
w10667 <= not w10665 and not w10666;
w10668 <= not w10664 and w10667;
w10669 <= w2796 and w3126;
w10670 <= w10668 and not w10669;
w10671 <= a(29) and not w10670;
w10672 <= a(29) and not w10671;
w10673 <= not w10670 and not w10671;
w10674 <= not w10672 and not w10673;
w10675 <= w10663 and w10674;
w10676 <= not w10663 and not w10674;
w10677 <= not w10675 and not w10676;
w10678 <= not w10496 and w10677;
w10679 <= w10496 and not w10677;
w10680 <= not w10678 and not w10679;
w10681 <= w10495 and not w10680;
w10682 <= not w10495 and w10680;
w10683 <= not w10681 and not w10682;
w10684 <= not w10484 and w10683;
w10685 <= w10484 and not w10683;
w10686 <= not w10684 and not w10685;
w10687 <= not w10483 and w10686;
w10688 <= w10686 and not w10687;
w10689 <= not w10483 and not w10687;
w10690 <= not w10688 and not w10689;
w10691 <= not w10320 and not w10327;
w10692 <= w10690 and w10691;
w10693 <= not w10690 and not w10691;
w10694 <= not w10692 and not w10693;
w10695 <= b(38) and w1370;
w10696 <= b(36) and w1506;
w10697 <= b(37) and w1365;
w10698 <= not w10696 and not w10697;
w10699 <= not w10695 and w10698;
w10700 <= w1373 and w4948;
w10701 <= w10699 and not w10700;
w10702 <= a(20) and not w10701;
w10703 <= a(20) and not w10702;
w10704 <= not w10701 and not w10702;
w10705 <= not w10703 and not w10704;
w10706 <= w10694 and not w10705;
w10707 <= w10694 and not w10706;
w10708 <= not w10705 and not w10706;
w10709 <= not w10707 and not w10708;
w10710 <= not w10340 and not w10346;
w10711 <= w10709 and w10710;
w10712 <= not w10709 and not w10710;
w10713 <= not w10711 and not w10712;
w10714 <= b(41) and w1045;
w10715 <= b(39) and w1134;
w10716 <= b(40) and w1040;
w10717 <= not w10715 and not w10716;
w10718 <= not w10714 and w10717;
w10719 <= w1048 and w5962;
w10720 <= w10718 and not w10719;
w10721 <= a(17) and not w10720;
w10722 <= a(17) and not w10721;
w10723 <= not w10720 and not w10721;
w10724 <= not w10722 and not w10723;
w10725 <= w10713 and not w10724;
w10726 <= w10713 and not w10725;
w10727 <= not w10724 and not w10725;
w10728 <= not w10726 and not w10727;
w10729 <= not w10359 and not w10365;
w10730 <= w10728 and w10729;
w10731 <= not w10728 and not w10729;
w10732 <= not w10730 and not w10731;
w10733 <= b(44) and w694;
w10734 <= b(42) and w799;
w10735 <= b(43) and w689;
w10736 <= not w10734 and not w10735;
w10737 <= not w10733 and w10736;
w10738 <= w697 and w6815;
w10739 <= w10737 and not w10738;
w10740 <= a(14) and not w10739;
w10741 <= a(14) and not w10740;
w10742 <= not w10739 and not w10740;
w10743 <= not w10741 and not w10742;
w10744 <= w10732 and not w10743;
w10745 <= not w10732 and w10743;
w10746 <= not w10383 and not w10745;
w10747 <= not w10744 and w10746;
w10748 <= not w10383 and not w10747;
w10749 <= not w10744 and not w10747;
w10750 <= not w10745 and w10749;
w10751 <= not w10748 and not w10750;
w10752 <= b(47) and w443;
w10753 <= b(45) and w510;
w10754 <= b(46) and w438;
w10755 <= not w10753 and not w10754;
w10756 <= not w10752 and w10755;
w10757 <= w446 and w7446;
w10758 <= w10756 and not w10757;
w10759 <= a(11) and not w10758;
w10760 <= a(11) and not w10759;
w10761 <= not w10758 and not w10759;
w10762 <= not w10760 and not w10761;
w10763 <= not w10751 and not w10762;
w10764 <= not w10751 and not w10763;
w10765 <= not w10762 and not w10763;
w10766 <= not w10764 and not w10765;
w10767 <= not w10472 and not w10766;
w10768 <= w10472 and w10766;
w10769 <= not w10767 and not w10768;
w10770 <= not w10471 and w10769;
w10771 <= not w10471 and not w10770;
w10772 <= w10769 and not w10770;
w10773 <= not w10771 and not w10772;
w10774 <= not w10460 and not w10773;
w10775 <= not w10460 and not w10774;
w10776 <= not w10773 and not w10774;
w10777 <= not w10775 and not w10776;
w10778 <= b(53) and w105;
w10779 <= b(51) and w146;
w10780 <= b(52) and w100;
w10781 <= not w10779 and not w10780;
w10782 <= not w10778 and w10781;
w10783 <= w108 and w9715;
w10784 <= w10782 and not w10783;
w10785 <= a(5) and not w10784;
w10786 <= a(5) and not w10785;
w10787 <= not w10784 and not w10785;
w10788 <= not w10786 and not w10787;
w10789 <= w10777 and w10788;
w10790 <= not w10777 and not w10788;
w10791 <= not w10789 and not w10790;
w10792 <= not w10459 and w10791;
w10793 <= w10459 and not w10791;
w10794 <= not w10792 and not w10793;
w10795 <= not w10457 and w10794;
w10796 <= w10794 and not w10795;
w10797 <= not w10457 and not w10795;
w10798 <= not w10796 and not w10797;
w10799 <= not w10434 and not w10437;
w10800 <= not w10798 and not w10799;
w10801 <= w10798 and w10799;
w10802 <= not w10800 and not w10801;
w10803 <= not w10790 and not w10792;
w10804 <= b(54) and w105;
w10805 <= b(52) and w146;
w10806 <= b(53) and w100;
w10807 <= not w10805 and not w10806;
w10808 <= not w10804 and w10807;
w10809 <= w108 and w9741;
w10810 <= w10808 and not w10809;
w10811 <= a(5) and not w10810;
w10812 <= a(5) and not w10811;
w10813 <= not w10810 and not w10811;
w10814 <= not w10812 and not w10813;
w10815 <= not w10770 and not w10774;
w10816 <= b(51) and w254;
w10817 <= b(49) and w284;
w10818 <= b(50) and w249;
w10819 <= not w10817 and not w10818;
w10820 <= not w10816 and w10819;
w10821 <= w257 and w8719;
w10822 <= w10820 and not w10821;
w10823 <= a(8) and not w10822;
w10824 <= a(8) and not w10823;
w10825 <= not w10822 and not w10823;
w10826 <= not w10824 and not w10825;
w10827 <= not w10763 and not w10767;
w10828 <= b(48) and w443;
w10829 <= b(46) and w510;
w10830 <= b(47) and w438;
w10831 <= not w10829 and not w10830;
w10832 <= not w10828 and w10831;
w10833 <= w446 and w7752;
w10834 <= w10832 and not w10833;
w10835 <= a(11) and not w10834;
w10836 <= a(11) and not w10835;
w10837 <= not w10834 and not w10835;
w10838 <= not w10836 and not w10837;
w10839 <= b(45) and w694;
w10840 <= b(43) and w799;
w10841 <= b(44) and w689;
w10842 <= not w10840 and not w10841;
w10843 <= not w10839 and w10842;
w10844 <= w697 and w7104;
w10845 <= w10843 and not w10844;
w10846 <= a(14) and not w10845;
w10847 <= a(14) and not w10846;
w10848 <= not w10845 and not w10846;
w10849 <= not w10847 and not w10848;
w10850 <= not w10725 and not w10731;
w10851 <= not w10687 and not w10693;
w10852 <= not w10682 and not w10684;
w10853 <= not w10676 and not w10678;
w10854 <= b(30) and w2793;
w10855 <= b(28) and w2986;
w10856 <= b(29) and w2788;
w10857 <= not w10855 and not w10856;
w10858 <= not w10854 and w10857;
w10859 <= w2796 and w3320;
w10860 <= w10858 and not w10859;
w10861 <= a(29) and not w10860;
w10862 <= a(29) and not w10861;
w10863 <= not w10860 and not w10861;
w10864 <= not w10862 and not w10863;
w10865 <= not w10230 and not w10624;
w10866 <= not w10621 and not w10865;
w10867 <= b(21) and w4778;
w10868 <= b(19) and w5020;
w10869 <= b(20) and w4773;
w10870 <= not w10868 and not w10869;
w10871 <= not w10867 and w10870;
w10872 <= w1727 and w4781;
w10873 <= w10871 and not w10872;
w10874 <= a(38) and not w10873;
w10875 <= a(38) and not w10874;
w10876 <= not w10873 and not w10874;
w10877 <= not w10875 and not w10876;
w10878 <= not w10602 and not w10606;
w10879 <= b(18) and w5520;
w10880 <= b(16) and w5802;
w10881 <= b(17) and w5515;
w10882 <= not w10880 and not w10881;
w10883 <= not w10879 and w10882;
w10884 <= w1309 and w5523;
w10885 <= w10883 and not w10884;
w10886 <= a(41) and not w10885;
w10887 <= a(41) and not w10886;
w10888 <= not w10885 and not w10886;
w10889 <= not w10887 and not w10888;
w10890 <= not w10595 and not w10599;
w10891 <= b(15) and w6338;
w10892 <= b(13) and w6645;
w10893 <= b(14) and w6333;
w10894 <= not w10892 and not w10893;
w10895 <= not w10891 and w10894;
w10896 <= w874 and w6341;
w10897 <= w10895 and not w10896;
w10898 <= a(44) and not w10897;
w10899 <= a(44) and not w10898;
w10900 <= not w10897 and not w10898;
w10901 <= not w10899 and not w10900;
w10902 <= not w10590 and not w10592;
w10903 <= b(12) and w7189;
w10904 <= b(10) and w7530;
w10905 <= b(11) and w7184;
w10906 <= not w10904 and not w10905;
w10907 <= not w10903 and w10906;
w10908 <= w585 and w7192;
w10909 <= w10907 and not w10908;
w10910 <= a(47) and not w10909;
w10911 <= a(47) and not w10910;
w10912 <= not w10909 and not w10910;
w10913 <= not w10911 and not w10912;
w10914 <= not w10584 and not w10586;
w10915 <= b(6) and w9082;
w10916 <= b(4) and w9475;
w10917 <= b(5) and w9077;
w10918 <= not w10916 and not w10917;
w10919 <= not w10915 and w10918;
w10920 <= w202 and w9085;
w10921 <= w10919 and not w10920;
w10922 <= a(53) and not w10921;
w10923 <= a(53) and not w10922;
w10924 <= not w10921 and not w10922;
w10925 <= not w10923 and not w10924;
w10926 <= a(56) and not a(57);
w10927 <= not a(56) and a(57);
w10928 <= not w10926 and not w10927;
w10929 <= b(0) and not w10928;
w10930 <= not w10551 and w10929;
w10931 <= w10551 and not w10929;
w10932 <= not w10930 and not w10931;
w10933 <= b(3) and w10169;
w10934 <= b(1) and w10539;
w10935 <= b(2) and w10164;
w10936 <= not w10934 and not w10935;
w10937 <= not w10933 and w10936;
w10938 <= w61 and w10172;
w10939 <= w10937 and not w10938;
w10940 <= a(56) and not w10939;
w10941 <= a(56) and not w10940;
w10942 <= not w10939 and not w10940;
w10943 <= not w10941 and not w10942;
w10944 <= not w10932 and not w10943;
w10945 <= w10932 and w10943;
w10946 <= not w10944 and not w10945;
w10947 <= not w10925 and w10946;
w10948 <= w10946 and not w10947;
w10949 <= not w10925 and not w10947;
w10950 <= not w10948 and not w10949;
w10951 <= not w10569 and w10950;
w10952 <= w10569 and not w10950;
w10953 <= not w10951 and not w10952;
w10954 <= b(9) and w8105;
w10955 <= b(7) and w8458;
w10956 <= b(8) and w8100;
w10957 <= not w10955 and not w10956;
w10958 <= not w10954 and w10957;
w10959 <= w394 and w8108;
w10960 <= w10958 and not w10959;
w10961 <= a(50) and not w10960;
w10962 <= a(50) and not w10961;
w10963 <= not w10960 and not w10961;
w10964 <= not w10962 and not w10963;
w10965 <= not w10953 and not w10964;
w10966 <= w10953 and w10964;
w10967 <= not w10965 and not w10966;
w10968 <= not w10914 and w10967;
w10969 <= w10914 and not w10967;
w10970 <= not w10968 and not w10969;
w10971 <= w10913 and not w10970;
w10972 <= not w10913 and w10970;
w10973 <= not w10971 and not w10972;
w10974 <= not w10902 and w10973;
w10975 <= w10902 and not w10973;
w10976 <= not w10974 and not w10975;
w10977 <= not w10901 and w10976;
w10978 <= w10901 and not w10976;
w10979 <= not w10977 and not w10978;
w10980 <= not w10890 and w10979;
w10981 <= w10890 and not w10979;
w10982 <= not w10980 and not w10981;
w10983 <= not w10889 and w10982;
w10984 <= not w10889 and not w10983;
w10985 <= w10982 and not w10983;
w10986 <= not w10984 and not w10985;
w10987 <= not w10878 and not w10986;
w10988 <= w10878 and not w10985;
w10989 <= not w10984 and w10988;
w10990 <= not w10987 and not w10989;
w10991 <= not w10877 and w10990;
w10992 <= w10877 and not w10990;
w10993 <= not w10991 and not w10992;
w10994 <= not w10866 and w10993;
w10995 <= w10866 and not w10993;
w10996 <= not w10994 and not w10995;
w10997 <= b(24) and w4030;
w10998 <= b(22) and w4275;
w10999 <= b(23) and w4025;
w11000 <= not w10998 and not w10999;
w11001 <= not w10997 and w11000;
w11002 <= w2201 and w4033;
w11003 <= w11001 and not w11002;
w11004 <= a(35) and not w11003;
w11005 <= a(35) and not w11004;
w11006 <= not w11003 and not w11004;
w11007 <= not w11005 and not w11006;
w11008 <= w10996 and not w11007;
w11009 <= w10996 and not w11008;
w11010 <= not w11007 and not w11008;
w11011 <= not w11009 and not w11010;
w11012 <= not w10639 and not w10643;
w11013 <= w11011 and w11012;
w11014 <= not w11011 and not w11012;
w11015 <= not w11013 and not w11014;
w11016 <= b(27) and w3381;
w11017 <= b(25) and w3586;
w11018 <= b(26) and w3376;
w11019 <= not w11017 and not w11018;
w11020 <= not w11016 and w11019;
w11021 <= w2733 and w3384;
w11022 <= w11020 and not w11021;
w11023 <= a(32) and not w11022;
w11024 <= a(32) and not w11023;
w11025 <= not w11022 and not w11023;
w11026 <= not w11024 and not w11025;
w11027 <= not w11015 and w11026;
w11028 <= w11015 and not w11026;
w11029 <= not w11027 and not w11028;
w11030 <= not w10661 and w11029;
w11031 <= w10661 and not w11029;
w11032 <= not w11030 and not w11031;
w11033 <= not w10864 and w11032;
w11034 <= w10864 and not w11032;
w11035 <= not w11033 and not w11034;
w11036 <= not w10853 and w11035;
w11037 <= w10853 and not w11035;
w11038 <= not w11036 and not w11037;
w11039 <= b(33) and w2282;
w11040 <= b(31) and w2428;
w11041 <= b(32) and w2277;
w11042 <= not w11040 and not w11041;
w11043 <= not w11039 and w11042;
w11044 <= w2285 and w3966;
w11045 <= w11043 and not w11044;
w11046 <= a(26) and not w11045;
w11047 <= a(26) and not w11046;
w11048 <= not w11045 and not w11046;
w11049 <= not w11047 and not w11048;
w11050 <= w11038 and not w11049;
w11051 <= w11038 and not w11050;
w11052 <= not w11049 and not w11050;
w11053 <= not w11051 and not w11052;
w11054 <= not w10852 and w11053;
w11055 <= w10852 and not w11053;
w11056 <= not w11054 and not w11055;
w11057 <= b(36) and w1791;
w11058 <= b(34) and w1941;
w11059 <= b(35) and w1786;
w11060 <= not w11058 and not w11059;
w11061 <= not w11057 and w11060;
w11062 <= w1794 and w4665;
w11063 <= w11061 and not w11062;
w11064 <= a(23) and not w11063;
w11065 <= a(23) and not w11064;
w11066 <= not w11063 and not w11064;
w11067 <= not w11065 and not w11066;
w11068 <= not w11056 and not w11067;
w11069 <= w11056 and w11067;
w11070 <= not w11068 and not w11069;
w11071 <= w10851 and not w11070;
w11072 <= not w10851 and w11070;
w11073 <= not w11071 and not w11072;
w11074 <= b(39) and w1370;
w11075 <= b(37) and w1506;
w11076 <= b(38) and w1365;
w11077 <= not w11075 and not w11076;
w11078 <= not w11074 and w11077;
w11079 <= w1373 and w5194;
w11080 <= w11078 and not w11079;
w11081 <= a(20) and not w11080;
w11082 <= a(20) and not w11081;
w11083 <= not w11080 and not w11081;
w11084 <= not w11082 and not w11083;
w11085 <= w11073 and not w11084;
w11086 <= w11073 and not w11085;
w11087 <= not w11084 and not w11085;
w11088 <= not w11086 and not w11087;
w11089 <= not w10706 and not w10712;
w11090 <= w11088 and w11089;
w11091 <= not w11088 and not w11089;
w11092 <= not w11090 and not w11091;
w11093 <= b(42) and w1045;
w11094 <= b(40) and w1134;
w11095 <= b(41) and w1040;
w11096 <= not w11094 and not w11095;
w11097 <= not w11093 and w11096;
w11098 <= w1048 and w6232;
w11099 <= w11097 and not w11098;
w11100 <= a(17) and not w11099;
w11101 <= a(17) and not w11100;
w11102 <= not w11099 and not w11100;
w11103 <= not w11101 and not w11102;
w11104 <= not w11092 and w11103;
w11105 <= w11092 and not w11103;
w11106 <= not w11104 and not w11105;
w11107 <= not w10850 and w11106;
w11108 <= w10850 and not w11106;
w11109 <= not w11107 and not w11108;
w11110 <= not w10849 and w11109;
w11111 <= not w10849 and not w11110;
w11112 <= w11109 and not w11110;
w11113 <= not w11111 and not w11112;
w11114 <= not w10749 and not w11113;
w11115 <= w10749 and not w11112;
w11116 <= not w11111 and w11115;
w11117 <= not w11114 and not w11116;
w11118 <= not w10838 and w11117;
w11119 <= not w10838 and not w11118;
w11120 <= w11117 and not w11118;
w11121 <= not w11119 and not w11120;
w11122 <= not w10827 and not w11121;
w11123 <= w10827 and not w11120;
w11124 <= not w11119 and w11123;
w11125 <= not w11122 and not w11124;
w11126 <= not w10826 and w11125;
w11127 <= not w10826 and not w11126;
w11128 <= w11125 and not w11126;
w11129 <= not w11127 and not w11128;
w11130 <= not w10815 and not w11129;
w11131 <= w10815 and not w11128;
w11132 <= not w11127 and w11131;
w11133 <= not w11130 and not w11132;
w11134 <= not w10814 and w11133;
w11135 <= not w10814 and not w11134;
w11136 <= w11133 and not w11134;
w11137 <= not w11135 and not w11136;
w11138 <= not w10803 and not w11137;
w11139 <= not w10803 and not w11138;
w11140 <= not w11137 and not w11138;
w11141 <= not w11139 and not w11140;
w11142 <= b(57) and w9;
w11143 <= b(55) and w27;
w11144 <= b(56) and w4;
w11145 <= not w11143 and not w11144;
w11146 <= not w11142 and w11145;
w11147 <= not w10447 and not w10449;
w11148 <= not b(56) and not b(57);
w11149 <= b(56) and b(57);
w11150 <= not w11148 and not w11149;
w11151 <= not w11147 and w11150;
w11152 <= w11147 and not w11150;
w11153 <= not w11151 and not w11152;
w11154 <= w12 and w11153;
w11155 <= w11146 and not w11154;
w11156 <= a(2) and not w11155;
w11157 <= a(2) and not w11156;
w11158 <= not w11155 and not w11156;
w11159 <= not w11157 and not w11158;
w11160 <= not w11141 and not w11159;
w11161 <= not w11141 and not w11160;
w11162 <= not w11159 and not w11160;
w11163 <= not w11161 and not w11162;
w11164 <= not w10795 and not w10800;
w11165 <= not w11163 and not w11164;
w11166 <= w11163 and w11164;
w11167 <= not w11165 and not w11166;
w11168 <= b(58) and w9;
w11169 <= b(56) and w27;
w11170 <= b(57) and w4;
w11171 <= not w11169 and not w11170;
w11172 <= not w11168 and w11171;
w11173 <= not w11149 and not w11151;
w11174 <= not b(57) and not b(58);
w11175 <= b(57) and b(58);
w11176 <= not w11174 and not w11175;
w11177 <= not w11173 and w11176;
w11178 <= w11173 and not w11176;
w11179 <= not w11177 and not w11178;
w11180 <= w12 and w11179;
w11181 <= w11172 and not w11180;
w11182 <= a(2) and not w11181;
w11183 <= a(2) and not w11182;
w11184 <= not w11181 and not w11182;
w11185 <= not w11183 and not w11184;
w11186 <= not w11134 and not w11138;
w11187 <= b(55) and w105;
w11188 <= b(53) and w146;
w11189 <= b(54) and w100;
w11190 <= not w11188 and not w11189;
w11191 <= not w11187 and w11190;
w11192 <= w108 and w10427;
w11193 <= w11191 and not w11192;
w11194 <= a(5) and not w11193;
w11195 <= a(5) and not w11194;
w11196 <= not w11193 and not w11194;
w11197 <= not w11195 and not w11196;
w11198 <= not w11126 and not w11130;
w11199 <= b(52) and w254;
w11200 <= b(50) and w284;
w11201 <= b(51) and w249;
w11202 <= not w11200 and not w11201;
w11203 <= not w11199 and w11202;
w11204 <= w257 and w9371;
w11205 <= w11203 and not w11204;
w11206 <= a(8) and not w11205;
w11207 <= a(8) and not w11206;
w11208 <= not w11205 and not w11206;
w11209 <= not w11207 and not w11208;
w11210 <= not w11118 and not w11122;
w11211 <= b(49) and w443;
w11212 <= b(47) and w510;
w11213 <= b(48) and w438;
w11214 <= not w11212 and not w11213;
w11215 <= not w11211 and w11214;
w11216 <= w446 and w8368;
w11217 <= w11215 and not w11216;
w11218 <= a(11) and not w11217;
w11219 <= a(11) and not w11218;
w11220 <= not w11217 and not w11218;
w11221 <= not w11219 and not w11220;
w11222 <= not w11110 and not w11114;
w11223 <= not w11105 and not w11107;
w11224 <= not w11033 and not w11036;
w11225 <= not w11028 and not w11030;
w11226 <= not w10983 and not w10987;
w11227 <= not w10972 and not w10974;
w11228 <= b(10) and w8105;
w11229 <= b(8) and w8458;
w11230 <= b(9) and w8100;
w11231 <= not w11229 and not w11230;
w11232 <= not w11228 and w11231;
w11233 <= w481 and w8108;
w11234 <= w11232 and not w11233;
w11235 <= a(50) and not w11234;
w11236 <= a(50) and not w11235;
w11237 <= not w11234 and not w11235;
w11238 <= not w11236 and not w11237;
w11239 <= not w10569 and not w10950;
w11240 <= not w10947 and not w11239;
w11241 <= b(7) and w9082;
w11242 <= b(5) and w9475;
w11243 <= b(6) and w9077;
w11244 <= not w11242 and not w11243;
w11245 <= not w11241 and w11244;
w11246 <= w227 and w9085;
w11247 <= w11245 and not w11246;
w11248 <= a(53) and not w11247;
w11249 <= a(53) and not w11248;
w11250 <= not w11247 and not w11248;
w11251 <= not w11249 and not w11250;
w11252 <= w10551 and w10929;
w11253 <= not w10944 and not w11252;
w11254 <= b(4) and w10169;
w11255 <= b(2) and w10539;
w11256 <= b(3) and w10164;
w11257 <= not w11255 and not w11256;
w11258 <= not w11254 and w11257;
w11259 <= w89 and w10172;
w11260 <= w11258 and not w11259;
w11261 <= a(56) and not w11260;
w11262 <= a(56) and not w11261;
w11263 <= not w11260 and not w11261;
w11264 <= not w11262 and not w11263;
w11265 <= a(59) and not w10929;
w11266 <= not a(57) and a(58);
w11267 <= a(57) and not a(58);
w11268 <= not w11266 and not w11267;
w11269 <= w10928 and not w11268;
w11270 <= b(0) and w11269;
w11271 <= not a(58) and a(59);
w11272 <= a(58) and not a(59);
w11273 <= not w11271 and not w11272;
w11274 <= not w10928 and w11273;
w11275 <= b(1) and w11274;
w11276 <= not w11270 and not w11275;
w11277 <= not w10928 and not w11273;
w11278 <= not w15 and w11277;
w11279 <= w11276 and not w11278;
w11280 <= a(59) and not w11279;
w11281 <= a(59) and not w11280;
w11282 <= not w11279 and not w11280;
w11283 <= not w11281 and not w11282;
w11284 <= w11265 and not w11283;
w11285 <= not w11265 and w11283;
w11286 <= not w11284 and not w11285;
w11287 <= w11264 and not w11286;
w11288 <= not w11264 and w11286;
w11289 <= not w11287 and not w11288;
w11290 <= not w11253 and w11289;
w11291 <= w11253 and not w11289;
w11292 <= not w11290 and not w11291;
w11293 <= w11251 and not w11292;
w11294 <= not w11251 and w11292;
w11295 <= not w11293 and not w11294;
w11296 <= not w11240 and w11295;
w11297 <= w11240 and not w11295;
w11298 <= not w11296 and not w11297;
w11299 <= not w11238 and w11298;
w11300 <= w11298 and not w11299;
w11301 <= not w11238 and not w11299;
w11302 <= not w11300 and not w11301;
w11303 <= not w10965 and not w10968;
w11304 <= w11302 and w11303;
w11305 <= not w11302 and not w11303;
w11306 <= not w11304 and not w11305;
w11307 <= b(13) and w7189;
w11308 <= b(11) and w7530;
w11309 <= b(12) and w7184;
w11310 <= not w11308 and not w11309;
w11311 <= not w11307 and w11310;
w11312 <= w751 and w7192;
w11313 <= w11311 and not w11312;
w11314 <= a(47) and not w11313;
w11315 <= a(47) and not w11314;
w11316 <= not w11313 and not w11314;
w11317 <= not w11315 and not w11316;
w11318 <= w11306 and not w11317;
w11319 <= not w11306 and w11317;
w11320 <= not w11227 and not w11319;
w11321 <= not w11318 and w11320;
w11322 <= not w11227 and not w11321;
w11323 <= not w11318 and not w11321;
w11324 <= not w11319 and w11323;
w11325 <= not w11322 and not w11324;
w11326 <= b(16) and w6338;
w11327 <= b(14) and w6645;
w11328 <= b(15) and w6333;
w11329 <= not w11327 and not w11328;
w11330 <= not w11326 and w11329;
w11331 <= w980 and w6341;
w11332 <= w11330 and not w11331;
w11333 <= a(44) and not w11332;
w11334 <= a(44) and not w11333;
w11335 <= not w11332 and not w11333;
w11336 <= not w11334 and not w11335;
w11337 <= not w11325 and not w11336;
w11338 <= not w11325 and not w11337;
w11339 <= not w11336 and not w11337;
w11340 <= not w11338 and not w11339;
w11341 <= not w10977 and not w10980;
w11342 <= w11340 and w11341;
w11343 <= not w11340 and not w11341;
w11344 <= not w11342 and not w11343;
w11345 <= b(19) and w5520;
w11346 <= b(17) and w5802;
w11347 <= b(18) and w5515;
w11348 <= not w11346 and not w11347;
w11349 <= not w11345 and w11348;
w11350 <= w1451 and w5523;
w11351 <= w11349 and not w11350;
w11352 <= a(41) and not w11351;
w11353 <= a(41) and not w11352;
w11354 <= not w11351 and not w11352;
w11355 <= not w11353 and not w11354;
w11356 <= w11344 and not w11355;
w11357 <= not w11344 and w11355;
w11358 <= not w11226 and not w11357;
w11359 <= not w11356 and w11358;
w11360 <= not w11226 and not w11359;
w11361 <= not w11356 and not w11359;
w11362 <= not w11357 and w11361;
w11363 <= not w11360 and not w11362;
w11364 <= b(22) and w4778;
w11365 <= b(20) and w5020;
w11366 <= b(21) and w4773;
w11367 <= not w11365 and not w11366;
w11368 <= not w11364 and w11367;
w11369 <= w1888 and w4781;
w11370 <= w11368 and not w11369;
w11371 <= a(38) and not w11370;
w11372 <= a(38) and not w11371;
w11373 <= not w11370 and not w11371;
w11374 <= not w11372 and not w11373;
w11375 <= not w11363 and not w11374;
w11376 <= not w11363 and not w11375;
w11377 <= not w11374 and not w11375;
w11378 <= not w11376 and not w11377;
w11379 <= not w10991 and not w10994;
w11380 <= w11378 and w11379;
w11381 <= not w11378 and not w11379;
w11382 <= not w11380 and not w11381;
w11383 <= b(25) and w4030;
w11384 <= b(23) and w4275;
w11385 <= b(24) and w4025;
w11386 <= not w11384 and not w11385;
w11387 <= not w11383 and w11386;
w11388 <= w2228 and w4033;
w11389 <= w11387 and not w11388;
w11390 <= a(35) and not w11389;
w11391 <= a(35) and not w11390;
w11392 <= not w11389 and not w11390;
w11393 <= not w11391 and not w11392;
w11394 <= w11382 and not w11393;
w11395 <= w11382 and not w11394;
w11396 <= not w11393 and not w11394;
w11397 <= not w11395 and not w11396;
w11398 <= not w11008 and not w11014;
w11399 <= w11397 and w11398;
w11400 <= not w11397 and not w11398;
w11401 <= not w11399 and not w11400;
w11402 <= b(28) and w3381;
w11403 <= b(26) and w3586;
w11404 <= b(27) and w3376;
w11405 <= not w11403 and not w11404;
w11406 <= not w11402 and w11405;
w11407 <= w2932 and w3384;
w11408 <= w11406 and not w11407;
w11409 <= a(32) and not w11408;
w11410 <= a(32) and not w11409;
w11411 <= not w11408 and not w11409;
w11412 <= not w11410 and not w11411;
w11413 <= w11401 and not w11412;
w11414 <= w11401 and not w11413;
w11415 <= not w11412 and not w11413;
w11416 <= not w11414 and not w11415;
w11417 <= not w11225 and w11416;
w11418 <= w11225 and not w11416;
w11419 <= not w11417 and not w11418;
w11420 <= b(31) and w2793;
w11421 <= b(29) and w2986;
w11422 <= b(30) and w2788;
w11423 <= not w11421 and not w11422;
w11424 <= not w11420 and w11423;
w11425 <= w2796 and w3539;
w11426 <= w11424 and not w11425;
w11427 <= a(29) and not w11426;
w11428 <= a(29) and not w11427;
w11429 <= not w11426 and not w11427;
w11430 <= not w11428 and not w11429;
w11431 <= not w11419 and not w11430;
w11432 <= w11419 and w11430;
w11433 <= not w11431 and not w11432;
w11434 <= w11224 and not w11433;
w11435 <= not w11224 and w11433;
w11436 <= not w11434 and not w11435;
w11437 <= b(34) and w2282;
w11438 <= b(32) and w2428;
w11439 <= b(33) and w2277;
w11440 <= not w11438 and not w11439;
w11441 <= not w11437 and w11440;
w11442 <= w2285 and w4209;
w11443 <= w11441 and not w11442;
w11444 <= a(26) and not w11443;
w11445 <= a(26) and not w11444;
w11446 <= not w11443 and not w11444;
w11447 <= not w11445 and not w11446;
w11448 <= w11436 and not w11447;
w11449 <= w11436 and not w11448;
w11450 <= not w11447 and not w11448;
w11451 <= not w11449 and not w11450;
w11452 <= not w10852 and not w11053;
w11453 <= not w11050 and not w11452;
w11454 <= w11451 and w11453;
w11455 <= not w11451 and not w11453;
w11456 <= not w11454 and not w11455;
w11457 <= b(37) and w1791;
w11458 <= b(35) and w1941;
w11459 <= b(36) and w1786;
w11460 <= not w11458 and not w11459;
w11461 <= not w11457 and w11460;
w11462 <= w1794 and w4924;
w11463 <= w11461 and not w11462;
w11464 <= a(23) and not w11463;
w11465 <= a(23) and not w11464;
w11466 <= not w11463 and not w11464;
w11467 <= not w11465 and not w11466;
w11468 <= w11456 and not w11467;
w11469 <= w11456 and not w11468;
w11470 <= not w11467 and not w11468;
w11471 <= not w11469 and not w11470;
w11472 <= not w11068 and not w11072;
w11473 <= w11471 and w11472;
w11474 <= not w11471 and not w11472;
w11475 <= not w11473 and not w11474;
w11476 <= b(40) and w1370;
w11477 <= b(38) and w1506;
w11478 <= b(39) and w1365;
w11479 <= not w11477 and not w11478;
w11480 <= not w11476 and w11479;
w11481 <= w1373 and w5698;
w11482 <= w11480 and not w11481;
w11483 <= a(20) and not w11482;
w11484 <= a(20) and not w11483;
w11485 <= not w11482 and not w11483;
w11486 <= not w11484 and not w11485;
w11487 <= w11475 and not w11486;
w11488 <= w11475 and not w11487;
w11489 <= not w11486 and not w11487;
w11490 <= not w11488 and not w11489;
w11491 <= not w11085 and not w11091;
w11492 <= w11490 and w11491;
w11493 <= not w11490 and not w11491;
w11494 <= not w11492 and not w11493;
w11495 <= b(43) and w1045;
w11496 <= b(41) and w1134;
w11497 <= b(42) and w1040;
w11498 <= not w11496 and not w11497;
w11499 <= not w11495 and w11498;
w11500 <= w1048 and w6258;
w11501 <= w11499 and not w11500;
w11502 <= a(17) and not w11501;
w11503 <= a(17) and not w11502;
w11504 <= not w11501 and not w11502;
w11505 <= not w11503 and not w11504;
w11506 <= w11494 and not w11505;
w11507 <= not w11494 and w11505;
w11508 <= not w11223 and not w11507;
w11509 <= not w11506 and w11508;
w11510 <= not w11223 and not w11509;
w11511 <= not w11506 and not w11509;
w11512 <= not w11507 and w11511;
w11513 <= not w11510 and not w11512;
w11514 <= b(46) and w694;
w11515 <= b(44) and w799;
w11516 <= b(45) and w689;
w11517 <= not w11515 and not w11516;
w11518 <= not w11514 and w11517;
w11519 <= w697 and w7420;
w11520 <= w11518 and not w11519;
w11521 <= a(14) and not w11520;
w11522 <= a(14) and not w11521;
w11523 <= not w11520 and not w11521;
w11524 <= not w11522 and not w11523;
w11525 <= w11513 and w11524;
w11526 <= not w11513 and not w11524;
w11527 <= not w11525 and not w11526;
w11528 <= not w11222 and w11527;
w11529 <= w11222 and not w11527;
w11530 <= not w11528 and not w11529;
w11531 <= w11221 and not w11530;
w11532 <= not w11221 and w11530;
w11533 <= not w11531 and not w11532;
w11534 <= not w11210 and w11533;
w11535 <= w11210 and not w11533;
w11536 <= not w11534 and not w11535;
w11537 <= w11209 and not w11536;
w11538 <= not w11209 and w11536;
w11539 <= not w11537 and not w11538;
w11540 <= not w11198 and w11539;
w11541 <= w11198 and not w11539;
w11542 <= not w11540 and not w11541;
w11543 <= w11197 and not w11542;
w11544 <= not w11197 and w11542;
w11545 <= not w11543 and not w11544;
w11546 <= not w11186 and w11545;
w11547 <= w11186 and not w11545;
w11548 <= not w11546 and not w11547;
w11549 <= not w11185 and w11548;
w11550 <= w11548 and not w11549;
w11551 <= not w11185 and not w11549;
w11552 <= not w11550 and not w11551;
w11553 <= not w11160 and not w11165;
w11554 <= not w11552 and not w11553;
w11555 <= w11552 and w11553;
w11556 <= not w11554 and not w11555;
w11557 <= not w11549 and not w11554;
w11558 <= not w11544 and not w11546;
w11559 <= not w11538 and not w11540;
w11560 <= b(53) and w254;
w11561 <= b(51) and w284;
w11562 <= b(52) and w249;
w11563 <= not w11561 and not w11562;
w11564 <= not w11560 and w11563;
w11565 <= w257 and w9715;
w11566 <= w11564 and not w11565;
w11567 <= a(8) and not w11566;
w11568 <= a(8) and not w11567;
w11569 <= not w11566 and not w11567;
w11570 <= not w11568 and not w11569;
w11571 <= not w11532 and not w11534;
w11572 <= b(50) and w443;
w11573 <= b(48) and w510;
w11574 <= b(49) and w438;
w11575 <= not w11573 and not w11574;
w11576 <= not w11572 and w11575;
w11577 <= w446 and w8692;
w11578 <= w11576 and not w11577;
w11579 <= a(11) and not w11578;
w11580 <= a(11) and not w11579;
w11581 <= not w11578 and not w11579;
w11582 <= not w11580 and not w11581;
w11583 <= not w11526 and not w11528;
w11584 <= not w11487 and not w11493;
w11585 <= b(35) and w2282;
w11586 <= b(33) and w2428;
w11587 <= b(34) and w2277;
w11588 <= not w11586 and not w11587;
w11589 <= not w11585 and w11588;
w11590 <= w2285 and w4439;
w11591 <= w11589 and not w11590;
w11592 <= a(26) and not w11591;
w11593 <= a(26) and not w11592;
w11594 <= not w11591 and not w11592;
w11595 <= not w11593 and not w11594;
w11596 <= not w11431 and not w11435;
w11597 <= not w11225 and not w11416;
w11598 <= not w11413 and not w11597;
w11599 <= not w11375 and not w11381;
w11600 <= not w11337 and not w11343;
w11601 <= b(17) and w6338;
w11602 <= b(15) and w6645;
w11603 <= b(16) and w6333;
w11604 <= not w11602 and not w11603;
w11605 <= not w11601 and w11604;
w11606 <= w1099 and w6341;
w11607 <= w11605 and not w11606;
w11608 <= a(44) and not w11607;
w11609 <= a(44) and not w11608;
w11610 <= not w11607 and not w11608;
w11611 <= not w11609 and not w11610;
w11612 <= b(14) and w7189;
w11613 <= b(12) and w7530;
w11614 <= b(13) and w7184;
w11615 <= not w11613 and not w11614;
w11616 <= not w11612 and w11615;
w11617 <= w777 and w7192;
w11618 <= w11616 and not w11617;
w11619 <= a(47) and not w11618;
w11620 <= a(47) and not w11619;
w11621 <= not w11618 and not w11619;
w11622 <= not w11620 and not w11621;
w11623 <= not w11299 and not w11305;
w11624 <= b(11) and w8105;
w11625 <= b(9) and w8458;
w11626 <= b(10) and w8100;
w11627 <= not w11625 and not w11626;
w11628 <= not w11624 and w11627;
w11629 <= w561 and w8108;
w11630 <= w11628 and not w11629;
w11631 <= a(50) and not w11630;
w11632 <= a(50) and not w11631;
w11633 <= not w11630 and not w11631;
w11634 <= not w11632 and not w11633;
w11635 <= not w11294 and not w11296;
w11636 <= not w11288 and not w11290;
w11637 <= b(2) and w11274;
w11638 <= w10928 and not w11273;
w11639 <= w11268 and w11638;
w11640 <= b(0) and w11639;
w11641 <= b(1) and w11269;
w11642 <= not w11640 and not w11641;
w11643 <= not w11637 and w11642;
w11644 <= w39 and w11277;
w11645 <= w11643 and not w11644;
w11646 <= a(59) and not w11645;
w11647 <= a(59) and not w11646;
w11648 <= not w11645 and not w11646;
w11649 <= not w11647 and not w11648;
w11650 <= not w11284 and w11649;
w11651 <= w11284 and not w11649;
w11652 <= not w11650 and not w11651;
w11653 <= b(5) and w10169;
w11654 <= b(3) and w10539;
w11655 <= b(4) and w10164;
w11656 <= not w11654 and not w11655;
w11657 <= not w11653 and w11656;
w11658 <= w137 and w10172;
w11659 <= w11657 and not w11658;
w11660 <= a(56) and not w11659;
w11661 <= a(56) and not w11660;
w11662 <= not w11659 and not w11660;
w11663 <= not w11661 and not w11662;
w11664 <= w11652 and not w11663;
w11665 <= not w11652 and w11663;
w11666 <= not w11636 and not w11665;
w11667 <= not w11664 and w11666;
w11668 <= not w11636 and not w11667;
w11669 <= not w11664 and not w11667;
w11670 <= not w11665 and w11669;
w11671 <= not w11668 and not w11670;
w11672 <= b(8) and w9082;
w11673 <= b(6) and w9475;
w11674 <= b(7) and w9077;
w11675 <= not w11673 and not w11674;
w11676 <= not w11672 and w11675;
w11677 <= w328 and w9085;
w11678 <= w11676 and not w11677;
w11679 <= a(53) and not w11678;
w11680 <= a(53) and not w11679;
w11681 <= not w11678 and not w11679;
w11682 <= not w11680 and not w11681;
w11683 <= w11671 and w11682;
w11684 <= not w11671 and not w11682;
w11685 <= not w11683 and not w11684;
w11686 <= not w11635 and w11685;
w11687 <= w11635 and not w11685;
w11688 <= not w11686 and not w11687;
w11689 <= w11634 and not w11688;
w11690 <= not w11634 and w11688;
w11691 <= not w11689 and not w11690;
w11692 <= not w11623 and w11691;
w11693 <= w11623 and not w11691;
w11694 <= not w11692 and not w11693;
w11695 <= not w11622 and w11694;
w11696 <= w11694 and not w11695;
w11697 <= not w11622 and not w11695;
w11698 <= not w11696 and not w11697;
w11699 <= not w11323 and not w11698;
w11700 <= w11323 and w11698;
w11701 <= not w11699 and not w11700;
w11702 <= not w11611 and w11701;
w11703 <= not w11611 and not w11702;
w11704 <= w11701 and not w11702;
w11705 <= not w11703 and not w11704;
w11706 <= not w11600 and not w11705;
w11707 <= not w11600 and not w11706;
w11708 <= not w11705 and not w11706;
w11709 <= not w11707 and not w11708;
w11710 <= b(20) and w5520;
w11711 <= b(18) and w5802;
w11712 <= b(19) and w5515;
w11713 <= not w11711 and not w11712;
w11714 <= not w11710 and w11713;
w11715 <= w1589 and w5523;
w11716 <= w11714 and not w11715;
w11717 <= a(41) and not w11716;
w11718 <= a(41) and not w11717;
w11719 <= not w11716 and not w11717;
w11720 <= not w11718 and not w11719;
w11721 <= not w11709 and not w11720;
w11722 <= not w11709 and not w11721;
w11723 <= not w11720 and not w11721;
w11724 <= not w11722 and not w11723;
w11725 <= not w11361 and w11724;
w11726 <= w11361 and not w11724;
w11727 <= not w11725 and not w11726;
w11728 <= b(23) and w4778;
w11729 <= b(21) and w5020;
w11730 <= b(22) and w4773;
w11731 <= not w11729 and not w11730;
w11732 <= not w11728 and w11731;
w11733 <= w2043 and w4781;
w11734 <= w11732 and not w11733;
w11735 <= a(38) and not w11734;
w11736 <= a(38) and not w11735;
w11737 <= not w11734 and not w11735;
w11738 <= not w11736 and not w11737;
w11739 <= not w11727 and not w11738;
w11740 <= w11727 and w11738;
w11741 <= not w11739 and not w11740;
w11742 <= w11599 and not w11741;
w11743 <= not w11599 and w11741;
w11744 <= not w11742 and not w11743;
w11745 <= b(26) and w4030;
w11746 <= b(24) and w4275;
w11747 <= b(25) and w4025;
w11748 <= not w11746 and not w11747;
w11749 <= not w11745 and w11748;
w11750 <= w2556 and w4033;
w11751 <= w11749 and not w11750;
w11752 <= a(35) and not w11751;
w11753 <= a(35) and not w11752;
w11754 <= not w11751 and not w11752;
w11755 <= not w11753 and not w11754;
w11756 <= w11744 and not w11755;
w11757 <= w11744 and not w11756;
w11758 <= not w11755 and not w11756;
w11759 <= not w11757 and not w11758;
w11760 <= not w11394 and not w11400;
w11761 <= w11759 and w11760;
w11762 <= not w11759 and not w11760;
w11763 <= not w11761 and not w11762;
w11764 <= b(29) and w3381;
w11765 <= b(27) and w3586;
w11766 <= b(28) and w3376;
w11767 <= not w11765 and not w11766;
w11768 <= not w11764 and w11767;
w11769 <= w3126 and w3384;
w11770 <= w11768 and not w11769;
w11771 <= a(32) and not w11770;
w11772 <= a(32) and not w11771;
w11773 <= not w11770 and not w11771;
w11774 <= not w11772 and not w11773;
w11775 <= w11763 and not w11774;
w11776 <= not w11763 and w11774;
w11777 <= not w11598 and not w11776;
w11778 <= not w11775 and w11777;
w11779 <= not w11598 and not w11778;
w11780 <= not w11775 and not w11778;
w11781 <= not w11776 and w11780;
w11782 <= not w11779 and not w11781;
w11783 <= b(32) and w2793;
w11784 <= b(30) and w2986;
w11785 <= b(31) and w2788;
w11786 <= not w11784 and not w11785;
w11787 <= not w11783 and w11786;
w11788 <= w2796 and w3756;
w11789 <= w11787 and not w11788;
w11790 <= a(29) and not w11789;
w11791 <= a(29) and not w11790;
w11792 <= not w11789 and not w11790;
w11793 <= not w11791 and not w11792;
w11794 <= w11782 and w11793;
w11795 <= not w11782 and not w11793;
w11796 <= not w11794 and not w11795;
w11797 <= not w11596 and w11796;
w11798 <= w11596 and not w11796;
w11799 <= not w11797 and not w11798;
w11800 <= not w11595 and w11799;
w11801 <= w11799 and not w11800;
w11802 <= not w11595 and not w11800;
w11803 <= not w11801 and not w11802;
w11804 <= not w11448 and not w11455;
w11805 <= w11803 and w11804;
w11806 <= not w11803 and not w11804;
w11807 <= not w11805 and not w11806;
w11808 <= b(38) and w1791;
w11809 <= b(36) and w1941;
w11810 <= b(37) and w1786;
w11811 <= not w11809 and not w11810;
w11812 <= not w11808 and w11811;
w11813 <= w1794 and w4948;
w11814 <= w11812 and not w11813;
w11815 <= a(23) and not w11814;
w11816 <= a(23) and not w11815;
w11817 <= not w11814 and not w11815;
w11818 <= not w11816 and not w11817;
w11819 <= w11807 and not w11818;
w11820 <= w11807 and not w11819;
w11821 <= not w11818 and not w11819;
w11822 <= not w11820 and not w11821;
w11823 <= not w11468 and not w11474;
w11824 <= w11822 and w11823;
w11825 <= not w11822 and not w11823;
w11826 <= not w11824 and not w11825;
w11827 <= b(41) and w1370;
w11828 <= b(39) and w1506;
w11829 <= b(40) and w1365;
w11830 <= not w11828 and not w11829;
w11831 <= not w11827 and w11830;
w11832 <= w1373 and w5962;
w11833 <= w11831 and not w11832;
w11834 <= a(20) and not w11833;
w11835 <= a(20) and not w11834;
w11836 <= not w11833 and not w11834;
w11837 <= not w11835 and not w11836;
w11838 <= w11826 and not w11837;
w11839 <= not w11826 and w11837;
w11840 <= not w11584 and not w11839;
w11841 <= not w11838 and w11840;
w11842 <= not w11584 and not w11841;
w11843 <= not w11838 and not w11841;
w11844 <= not w11839 and w11843;
w11845 <= not w11842 and not w11844;
w11846 <= b(44) and w1045;
w11847 <= b(42) and w1134;
w11848 <= b(43) and w1040;
w11849 <= not w11847 and not w11848;
w11850 <= not w11846 and w11849;
w11851 <= w1048 and w6815;
w11852 <= w11850 and not w11851;
w11853 <= a(17) and not w11852;
w11854 <= a(17) and not w11853;
w11855 <= not w11852 and not w11853;
w11856 <= not w11854 and not w11855;
w11857 <= not w11845 and not w11856;
w11858 <= not w11845 and not w11857;
w11859 <= not w11856 and not w11857;
w11860 <= not w11858 and not w11859;
w11861 <= not w11511 and w11860;
w11862 <= w11511 and not w11860;
w11863 <= not w11861 and not w11862;
w11864 <= b(47) and w694;
w11865 <= b(45) and w799;
w11866 <= b(46) and w689;
w11867 <= not w11865 and not w11866;
w11868 <= not w11864 and w11867;
w11869 <= w697 and w7446;
w11870 <= w11868 and not w11869;
w11871 <= a(14) and not w11870;
w11872 <= a(14) and not w11871;
w11873 <= not w11870 and not w11871;
w11874 <= not w11872 and not w11873;
w11875 <= not w11863 and not w11874;
w11876 <= w11863 and w11874;
w11877 <= not w11875 and not w11876;
w11878 <= not w11583 and w11877;
w11879 <= w11583 and not w11877;
w11880 <= not w11878 and not w11879;
w11881 <= not w11582 and w11880;
w11882 <= w11880 and not w11881;
w11883 <= not w11582 and not w11881;
w11884 <= not w11882 and not w11883;
w11885 <= not w11571 and not w11884;
w11886 <= w11571 and w11884;
w11887 <= not w11885 and not w11886;
w11888 <= not w11570 and w11887;
w11889 <= not w11570 and not w11888;
w11890 <= w11887 and not w11888;
w11891 <= not w11889 and not w11890;
w11892 <= not w11559 and not w11891;
w11893 <= not w11559 and not w11892;
w11894 <= not w11891 and not w11892;
w11895 <= not w11893 and not w11894;
w11896 <= b(56) and w105;
w11897 <= b(54) and w146;
w11898 <= b(55) and w100;
w11899 <= not w11897 and not w11898;
w11900 <= not w11896 and w11899;
w11901 <= w108 and w10451;
w11902 <= w11900 and not w11901;
w11903 <= a(5) and not w11902;
w11904 <= a(5) and not w11903;
w11905 <= not w11902 and not w11903;
w11906 <= not w11904 and not w11905;
w11907 <= not w11895 and not w11906;
w11908 <= not w11895 and not w11907;
w11909 <= not w11906 and not w11907;
w11910 <= not w11908 and not w11909;
w11911 <= b(59) and w9;
w11912 <= b(57) and w27;
w11913 <= b(58) and w4;
w11914 <= not w11912 and not w11913;
w11915 <= not w11911 and w11914;
w11916 <= not w11175 and not w11177;
w11917 <= not b(58) and not b(59);
w11918 <= b(58) and b(59);
w11919 <= not w11917 and not w11918;
w11920 <= not w11916 and w11919;
w11921 <= w11916 and not w11919;
w11922 <= not w11920 and not w11921;
w11923 <= w12 and w11922;
w11924 <= w11915 and not w11923;
w11925 <= a(2) and not w11924;
w11926 <= a(2) and not w11925;
w11927 <= not w11924 and not w11925;
w11928 <= not w11926 and not w11927;
w11929 <= not w11910 and w11928;
w11930 <= w11910 and not w11928;
w11931 <= not w11929 and not w11930;
w11932 <= not w11558 and not w11931;
w11933 <= not w11558 and not w11932;
w11934 <= not w11931 and not w11932;
w11935 <= not w11933 and not w11934;
w11936 <= not w11557 and not w11935;
w11937 <= w11557 and not w11934;
w11938 <= not w11933 and w11937;
w11939 <= not w11936 and not w11938;
w11940 <= not w11932 and not w11936;
w11941 <= not w11910 and not w11928;
w11942 <= not w11907 and not w11941;
w11943 <= b(60) and w9;
w11944 <= b(58) and w27;
w11945 <= b(59) and w4;
w11946 <= not w11944 and not w11945;
w11947 <= not w11943 and w11946;
w11948 <= not w11918 and not w11920;
w11949 <= not b(59) and not b(60);
w11950 <= b(59) and b(60);
w11951 <= not w11949 and not w11950;
w11952 <= not w11948 and w11951;
w11953 <= w11948 and not w11951;
w11954 <= not w11952 and not w11953;
w11955 <= w12 and w11954;
w11956 <= w11947 and not w11955;
w11957 <= a(2) and not w11956;
w11958 <= a(2) and not w11957;
w11959 <= not w11956 and not w11957;
w11960 <= not w11958 and not w11959;
w11961 <= b(57) and w105;
w11962 <= b(55) and w146;
w11963 <= b(56) and w100;
w11964 <= not w11962 and not w11963;
w11965 <= not w11961 and w11964;
w11966 <= w108 and w11153;
w11967 <= w11965 and not w11966;
w11968 <= a(5) and not w11967;
w11969 <= a(5) and not w11968;
w11970 <= not w11967 and not w11968;
w11971 <= not w11969 and not w11970;
w11972 <= not w11888 and not w11892;
w11973 <= b(54) and w254;
w11974 <= b(52) and w284;
w11975 <= b(53) and w249;
w11976 <= not w11974 and not w11975;
w11977 <= not w11973 and w11976;
w11978 <= w257 and w9741;
w11979 <= w11977 and not w11978;
w11980 <= a(8) and not w11979;
w11981 <= a(8) and not w11980;
w11982 <= not w11979 and not w11980;
w11983 <= not w11981 and not w11982;
w11984 <= not w11881 and not w11885;
w11985 <= b(51) and w443;
w11986 <= b(49) and w510;
w11987 <= b(50) and w438;
w11988 <= not w11986 and not w11987;
w11989 <= not w11985 and w11988;
w11990 <= w446 and w8719;
w11991 <= w11989 and not w11990;
w11992 <= a(11) and not w11991;
w11993 <= a(11) and not w11992;
w11994 <= not w11991 and not w11992;
w11995 <= not w11993 and not w11994;
w11996 <= not w11875 and not w11878;
w11997 <= b(48) and w694;
w11998 <= b(46) and w799;
w11999 <= b(47) and w689;
w12000 <= not w11998 and not w11999;
w12001 <= not w11997 and w12000;
w12002 <= w697 and w7752;
w12003 <= w12001 and not w12002;
w12004 <= a(14) and not w12003;
w12005 <= a(14) and not w12004;
w12006 <= not w12003 and not w12004;
w12007 <= not w12005 and not w12006;
w12008 <= not w11511 and not w11860;
w12009 <= not w11857 and not w12008;
w12010 <= b(45) and w1045;
w12011 <= b(43) and w1134;
w12012 <= b(44) and w1040;
w12013 <= not w12011 and not w12012;
w12014 <= not w12010 and w12013;
w12015 <= w1048 and w7104;
w12016 <= w12014 and not w12015;
w12017 <= a(17) and not w12016;
w12018 <= a(17) and not w12017;
w12019 <= not w12016 and not w12017;
w12020 <= not w12018 and not w12019;
w12021 <= not w11800 and not w11806;
w12022 <= not w11795 and not w11797;
w12023 <= b(33) and w2793;
w12024 <= b(31) and w2986;
w12025 <= b(32) and w2788;
w12026 <= not w12024 and not w12025;
w12027 <= not w12023 and w12026;
w12028 <= w2796 and w3966;
w12029 <= w12027 and not w12028;
w12030 <= a(29) and not w12029;
w12031 <= a(29) and not w12030;
w12032 <= not w12029 and not w12030;
w12033 <= not w12031 and not w12032;
w12034 <= not w11361 and not w11724;
w12035 <= not w11721 and not w12034;
w12036 <= b(21) and w5520;
w12037 <= b(19) and w5802;
w12038 <= b(20) and w5515;
w12039 <= not w12037 and not w12038;
w12040 <= not w12036 and w12039;
w12041 <= w1727 and w5523;
w12042 <= w12040 and not w12041;
w12043 <= a(41) and not w12042;
w12044 <= a(41) and not w12043;
w12045 <= not w12042 and not w12043;
w12046 <= not w12044 and not w12045;
w12047 <= not w11702 and not w11706;
w12048 <= b(18) and w6338;
w12049 <= b(16) and w6645;
w12050 <= b(17) and w6333;
w12051 <= not w12049 and not w12050;
w12052 <= not w12048 and w12051;
w12053 <= w1309 and w6341;
w12054 <= w12052 and not w12053;
w12055 <= a(44) and not w12054;
w12056 <= a(44) and not w12055;
w12057 <= not w12054 and not w12055;
w12058 <= not w12056 and not w12057;
w12059 <= not w11695 and not w11699;
w12060 <= b(15) and w7189;
w12061 <= b(13) and w7530;
w12062 <= b(14) and w7184;
w12063 <= not w12061 and not w12062;
w12064 <= not w12060 and w12063;
w12065 <= w874 and w7192;
w12066 <= w12064 and not w12065;
w12067 <= a(47) and not w12066;
w12068 <= a(47) and not w12067;
w12069 <= not w12066 and not w12067;
w12070 <= not w12068 and not w12069;
w12071 <= not w11690 and not w11692;
w12072 <= b(12) and w8105;
w12073 <= b(10) and w8458;
w12074 <= b(11) and w8100;
w12075 <= not w12073 and not w12074;
w12076 <= not w12072 and w12075;
w12077 <= w585 and w8108;
w12078 <= w12076 and not w12077;
w12079 <= a(50) and not w12078;
w12080 <= a(50) and not w12079;
w12081 <= not w12078 and not w12079;
w12082 <= not w12080 and not w12081;
w12083 <= not w11684 and not w11686;
w12084 <= b(6) and w10169;
w12085 <= b(4) and w10539;
w12086 <= b(5) and w10164;
w12087 <= not w12085 and not w12086;
w12088 <= not w12084 and w12087;
w12089 <= w202 and w10172;
w12090 <= w12088 and not w12089;
w12091 <= a(56) and not w12090;
w12092 <= a(56) and not w12091;
w12093 <= not w12090 and not w12091;
w12094 <= not w12092 and not w12093;
w12095 <= a(59) and not a(60);
w12096 <= not a(59) and a(60);
w12097 <= not w12095 and not w12096;
w12098 <= b(0) and not w12097;
w12099 <= not w11651 and w12098;
w12100 <= w11651 and not w12098;
w12101 <= not w12099 and not w12100;
w12102 <= b(3) and w11274;
w12103 <= b(1) and w11639;
w12104 <= b(2) and w11269;
w12105 <= not w12103 and not w12104;
w12106 <= not w12102 and w12105;
w12107 <= w61 and w11277;
w12108 <= w12106 and not w12107;
w12109 <= a(59) and not w12108;
w12110 <= a(59) and not w12109;
w12111 <= not w12108 and not w12109;
w12112 <= not w12110 and not w12111;
w12113 <= not w12101 and not w12112;
w12114 <= w12101 and w12112;
w12115 <= not w12113 and not w12114;
w12116 <= not w12094 and w12115;
w12117 <= w12115 and not w12116;
w12118 <= not w12094 and not w12116;
w12119 <= not w12117 and not w12118;
w12120 <= not w11669 and w12119;
w12121 <= w11669 and not w12119;
w12122 <= not w12120 and not w12121;
w12123 <= b(9) and w9082;
w12124 <= b(7) and w9475;
w12125 <= b(8) and w9077;
w12126 <= not w12124 and not w12125;
w12127 <= not w12123 and w12126;
w12128 <= w394 and w9085;
w12129 <= w12127 and not w12128;
w12130 <= a(53) and not w12129;
w12131 <= a(53) and not w12130;
w12132 <= not w12129 and not w12130;
w12133 <= not w12131 and not w12132;
w12134 <= not w12122 and not w12133;
w12135 <= w12122 and w12133;
w12136 <= not w12134 and not w12135;
w12137 <= not w12083 and w12136;
w12138 <= w12083 and not w12136;
w12139 <= not w12137 and not w12138;
w12140 <= w12082 and not w12139;
w12141 <= not w12082 and w12139;
w12142 <= not w12140 and not w12141;
w12143 <= not w12071 and w12142;
w12144 <= w12071 and not w12142;
w12145 <= not w12143 and not w12144;
w12146 <= not w12070 and w12145;
w12147 <= w12070 and not w12145;
w12148 <= not w12146 and not w12147;
w12149 <= not w12059 and w12148;
w12150 <= w12059 and not w12148;
w12151 <= not w12149 and not w12150;
w12152 <= not w12058 and w12151;
w12153 <= not w12058 and not w12152;
w12154 <= w12151 and not w12152;
w12155 <= not w12153 and not w12154;
w12156 <= not w12047 and not w12155;
w12157 <= w12047 and not w12154;
w12158 <= not w12153 and w12157;
w12159 <= not w12156 and not w12158;
w12160 <= not w12046 and w12159;
w12161 <= w12046 and not w12159;
w12162 <= not w12160 and not w12161;
w12163 <= not w12035 and w12162;
w12164 <= w12035 and not w12162;
w12165 <= not w12163 and not w12164;
w12166 <= b(24) and w4778;
w12167 <= b(22) and w5020;
w12168 <= b(23) and w4773;
w12169 <= not w12167 and not w12168;
w12170 <= not w12166 and w12169;
w12171 <= w2201 and w4781;
w12172 <= w12170 and not w12171;
w12173 <= a(38) and not w12172;
w12174 <= a(38) and not w12173;
w12175 <= not w12172 and not w12173;
w12176 <= not w12174 and not w12175;
w12177 <= w12165 and not w12176;
w12178 <= w12165 and not w12177;
w12179 <= not w12176 and not w12177;
w12180 <= not w12178 and not w12179;
w12181 <= not w11739 and not w11743;
w12182 <= w12180 and w12181;
w12183 <= not w12180 and not w12181;
w12184 <= not w12182 and not w12183;
w12185 <= b(27) and w4030;
w12186 <= b(25) and w4275;
w12187 <= b(26) and w4025;
w12188 <= not w12186 and not w12187;
w12189 <= not w12185 and w12188;
w12190 <= w2733 and w4033;
w12191 <= w12189 and not w12190;
w12192 <= a(35) and not w12191;
w12193 <= a(35) and not w12192;
w12194 <= not w12191 and not w12192;
w12195 <= not w12193 and not w12194;
w12196 <= w12184 and not w12195;
w12197 <= w12184 and not w12196;
w12198 <= not w12195 and not w12196;
w12199 <= not w12197 and not w12198;
w12200 <= not w11756 and not w11762;
w12201 <= w12199 and w12200;
w12202 <= not w12199 and not w12200;
w12203 <= not w12201 and not w12202;
w12204 <= b(30) and w3381;
w12205 <= b(28) and w3586;
w12206 <= b(29) and w3376;
w12207 <= not w12205 and not w12206;
w12208 <= not w12204 and w12207;
w12209 <= w3320 and w3384;
w12210 <= w12208 and not w12209;
w12211 <= a(32) and not w12210;
w12212 <= a(32) and not w12211;
w12213 <= not w12210 and not w12211;
w12214 <= not w12212 and not w12213;
w12215 <= not w12203 and w12214;
w12216 <= w12203 and not w12214;
w12217 <= not w12215 and not w12216;
w12218 <= not w11780 and w12217;
w12219 <= w11780 and not w12217;
w12220 <= not w12218 and not w12219;
w12221 <= not w12033 and w12220;
w12222 <= w12220 and not w12221;
w12223 <= not w12033 and not w12221;
w12224 <= not w12222 and not w12223;
w12225 <= not w12022 and w12224;
w12226 <= w12022 and not w12224;
w12227 <= not w12225 and not w12226;
w12228 <= b(36) and w2282;
w12229 <= b(34) and w2428;
w12230 <= b(35) and w2277;
w12231 <= not w12229 and not w12230;
w12232 <= not w12228 and w12231;
w12233 <= w2285 and w4665;
w12234 <= w12232 and not w12233;
w12235 <= a(26) and not w12234;
w12236 <= a(26) and not w12235;
w12237 <= not w12234 and not w12235;
w12238 <= not w12236 and not w12237;
w12239 <= not w12227 and not w12238;
w12240 <= w12227 and w12238;
w12241 <= not w12239 and not w12240;
w12242 <= w12021 and not w12241;
w12243 <= not w12021 and w12241;
w12244 <= not w12242 and not w12243;
w12245 <= b(39) and w1791;
w12246 <= b(37) and w1941;
w12247 <= b(38) and w1786;
w12248 <= not w12246 and not w12247;
w12249 <= not w12245 and w12248;
w12250 <= w1794 and w5194;
w12251 <= w12249 and not w12250;
w12252 <= a(23) and not w12251;
w12253 <= a(23) and not w12252;
w12254 <= not w12251 and not w12252;
w12255 <= not w12253 and not w12254;
w12256 <= w12244 and not w12255;
w12257 <= w12244 and not w12256;
w12258 <= not w12255 and not w12256;
w12259 <= not w12257 and not w12258;
w12260 <= not w11819 and not w11825;
w12261 <= w12259 and w12260;
w12262 <= not w12259 and not w12260;
w12263 <= not w12261 and not w12262;
w12264 <= b(42) and w1370;
w12265 <= b(40) and w1506;
w12266 <= b(41) and w1365;
w12267 <= not w12265 and not w12266;
w12268 <= not w12264 and w12267;
w12269 <= w1373 and w6232;
w12270 <= w12268 and not w12269;
w12271 <= a(20) and not w12270;
w12272 <= a(20) and not w12271;
w12273 <= not w12270 and not w12271;
w12274 <= not w12272 and not w12273;
w12275 <= not w12263 and w12274;
w12276 <= w12263 and not w12274;
w12277 <= not w12275 and not w12276;
w12278 <= not w11843 and w12277;
w12279 <= w11843 and not w12277;
w12280 <= not w12278 and not w12279;
w12281 <= not w12020 and w12280;
w12282 <= not w12020 and not w12281;
w12283 <= w12280 and not w12281;
w12284 <= not w12282 and not w12283;
w12285 <= not w12009 and not w12284;
w12286 <= w12009 and not w12283;
w12287 <= not w12282 and w12286;
w12288 <= not w12285 and not w12287;
w12289 <= not w12007 and w12288;
w12290 <= not w12007 and not w12289;
w12291 <= w12288 and not w12289;
w12292 <= not w12290 and not w12291;
w12293 <= not w11996 and not w12292;
w12294 <= w11996 and not w12291;
w12295 <= not w12290 and w12294;
w12296 <= not w12293 and not w12295;
w12297 <= not w11995 and w12296;
w12298 <= not w11995 and not w12297;
w12299 <= w12296 and not w12297;
w12300 <= not w12298 and not w12299;
w12301 <= not w11984 and not w12300;
w12302 <= w11984 and not w12299;
w12303 <= not w12298 and w12302;
w12304 <= not w12301 and not w12303;
w12305 <= not w11983 and w12304;
w12306 <= w11983 and not w12304;
w12307 <= not w12305 and not w12306;
w12308 <= not w11972 and w12307;
w12309 <= w11972 and not w12307;
w12310 <= not w12308 and not w12309;
w12311 <= not w11971 and w12310;
w12312 <= w11971 and not w12310;
w12313 <= not w12311 and not w12312;
w12314 <= not w11960 and w12313;
w12315 <= w11960 and not w12313;
w12316 <= not w12314 and not w12315;
w12317 <= not w11942 and w12316;
w12318 <= w11942 and not w12316;
w12319 <= not w12317 and not w12318;
w12320 <= not w11940 and w12319;
w12321 <= w11940 and not w12319;
w12322 <= not w12320 and not w12321;
w12323 <= b(55) and w254;
w12324 <= b(53) and w284;
w12325 <= b(54) and w249;
w12326 <= not w12324 and not w12325;
w12327 <= not w12323 and w12326;
w12328 <= w257 and w10427;
w12329 <= w12327 and not w12328;
w12330 <= a(8) and not w12329;
w12331 <= a(8) and not w12330;
w12332 <= not w12329 and not w12330;
w12333 <= not w12331 and not w12332;
w12334 <= not w12297 and not w12301;
w12335 <= b(52) and w443;
w12336 <= b(50) and w510;
w12337 <= b(51) and w438;
w12338 <= not w12336 and not w12337;
w12339 <= not w12335 and w12338;
w12340 <= w446 and w9371;
w12341 <= w12339 and not w12340;
w12342 <= a(11) and not w12341;
w12343 <= a(11) and not w12342;
w12344 <= not w12341 and not w12342;
w12345 <= not w12343 and not w12344;
w12346 <= not w12289 and not w12293;
w12347 <= b(49) and w694;
w12348 <= b(47) and w799;
w12349 <= b(48) and w689;
w12350 <= not w12348 and not w12349;
w12351 <= not w12347 and w12350;
w12352 <= w697 and w8368;
w12353 <= w12351 and not w12352;
w12354 <= a(14) and not w12353;
w12355 <= a(14) and not w12354;
w12356 <= not w12353 and not w12354;
w12357 <= not w12355 and not w12356;
w12358 <= not w12281 and not w12285;
w12359 <= not w12276 and not w12278;
w12360 <= not w12022 and not w12224;
w12361 <= not w12221 and not w12360;
w12362 <= not w12216 and not w12218;
w12363 <= not w12152 and not w12156;
w12364 <= not w12141 and not w12143;
w12365 <= b(10) and w9082;
w12366 <= b(8) and w9475;
w12367 <= b(9) and w9077;
w12368 <= not w12366 and not w12367;
w12369 <= not w12365 and w12368;
w12370 <= w481 and w9085;
w12371 <= w12369 and not w12370;
w12372 <= a(53) and not w12371;
w12373 <= a(53) and not w12372;
w12374 <= not w12371 and not w12372;
w12375 <= not w12373 and not w12374;
w12376 <= not w11669 and not w12119;
w12377 <= not w12116 and not w12376;
w12378 <= b(7) and w10169;
w12379 <= b(5) and w10539;
w12380 <= b(6) and w10164;
w12381 <= not w12379 and not w12380;
w12382 <= not w12378 and w12381;
w12383 <= w227 and w10172;
w12384 <= w12382 and not w12383;
w12385 <= a(56) and not w12384;
w12386 <= a(56) and not w12385;
w12387 <= not w12384 and not w12385;
w12388 <= not w12386 and not w12387;
w12389 <= w11651 and w12098;
w12390 <= not w12113 and not w12389;
w12391 <= b(4) and w11274;
w12392 <= b(2) and w11639;
w12393 <= b(3) and w11269;
w12394 <= not w12392 and not w12393;
w12395 <= not w12391 and w12394;
w12396 <= w89 and w11277;
w12397 <= w12395 and not w12396;
w12398 <= a(59) and not w12397;
w12399 <= a(59) and not w12398;
w12400 <= not w12397 and not w12398;
w12401 <= not w12399 and not w12400;
w12402 <= a(62) and not w12098;
w12403 <= not a(60) and a(61);
w12404 <= a(60) and not a(61);
w12405 <= not w12403 and not w12404;
w12406 <= w12097 and not w12405;
w12407 <= b(0) and w12406;
w12408 <= not a(61) and a(62);
w12409 <= a(61) and not a(62);
w12410 <= not w12408 and not w12409;
w12411 <= not w12097 and w12410;
w12412 <= b(1) and w12411;
w12413 <= not w12407 and not w12412;
w12414 <= not w12097 and not w12410;
w12415 <= not w15 and w12414;
w12416 <= w12413 and not w12415;
w12417 <= a(62) and not w12416;
w12418 <= a(62) and not w12417;
w12419 <= not w12416 and not w12417;
w12420 <= not w12418 and not w12419;
w12421 <= w12402 and not w12420;
w12422 <= not w12402 and w12420;
w12423 <= not w12421 and not w12422;
w12424 <= w12401 and not w12423;
w12425 <= not w12401 and w12423;
w12426 <= not w12424 and not w12425;
w12427 <= not w12390 and w12426;
w12428 <= w12390 and not w12426;
w12429 <= not w12427 and not w12428;
w12430 <= w12388 and not w12429;
w12431 <= not w12388 and w12429;
w12432 <= not w12430 and not w12431;
w12433 <= not w12377 and w12432;
w12434 <= w12377 and not w12432;
w12435 <= not w12433 and not w12434;
w12436 <= not w12375 and w12435;
w12437 <= w12435 and not w12436;
w12438 <= not w12375 and not w12436;
w12439 <= not w12437 and not w12438;
w12440 <= not w12134 and not w12137;
w12441 <= w12439 and w12440;
w12442 <= not w12439 and not w12440;
w12443 <= not w12441 and not w12442;
w12444 <= b(13) and w8105;
w12445 <= b(11) and w8458;
w12446 <= b(12) and w8100;
w12447 <= not w12445 and not w12446;
w12448 <= not w12444 and w12447;
w12449 <= w751 and w8108;
w12450 <= w12448 and not w12449;
w12451 <= a(50) and not w12450;
w12452 <= a(50) and not w12451;
w12453 <= not w12450 and not w12451;
w12454 <= not w12452 and not w12453;
w12455 <= w12443 and not w12454;
w12456 <= not w12443 and w12454;
w12457 <= not w12364 and not w12456;
w12458 <= not w12455 and w12457;
w12459 <= not w12364 and not w12458;
w12460 <= not w12455 and not w12458;
w12461 <= not w12456 and w12460;
w12462 <= not w12459 and not w12461;
w12463 <= b(16) and w7189;
w12464 <= b(14) and w7530;
w12465 <= b(15) and w7184;
w12466 <= not w12464 and not w12465;
w12467 <= not w12463 and w12466;
w12468 <= w980 and w7192;
w12469 <= w12467 and not w12468;
w12470 <= a(47) and not w12469;
w12471 <= a(47) and not w12470;
w12472 <= not w12469 and not w12470;
w12473 <= not w12471 and not w12472;
w12474 <= not w12462 and not w12473;
w12475 <= not w12462 and not w12474;
w12476 <= not w12473 and not w12474;
w12477 <= not w12475 and not w12476;
w12478 <= not w12146 and not w12149;
w12479 <= w12477 and w12478;
w12480 <= not w12477 and not w12478;
w12481 <= not w12479 and not w12480;
w12482 <= b(19) and w6338;
w12483 <= b(17) and w6645;
w12484 <= b(18) and w6333;
w12485 <= not w12483 and not w12484;
w12486 <= not w12482 and w12485;
w12487 <= w1451 and w6341;
w12488 <= w12486 and not w12487;
w12489 <= a(44) and not w12488;
w12490 <= a(44) and not w12489;
w12491 <= not w12488 and not w12489;
w12492 <= not w12490 and not w12491;
w12493 <= w12481 and not w12492;
w12494 <= not w12481 and w12492;
w12495 <= not w12363 and not w12494;
w12496 <= not w12493 and w12495;
w12497 <= not w12363 and not w12496;
w12498 <= not w12493 and not w12496;
w12499 <= not w12494 and w12498;
w12500 <= not w12497 and not w12499;
w12501 <= b(22) and w5520;
w12502 <= b(20) and w5802;
w12503 <= b(21) and w5515;
w12504 <= not w12502 and not w12503;
w12505 <= not w12501 and w12504;
w12506 <= w1888 and w5523;
w12507 <= w12505 and not w12506;
w12508 <= a(41) and not w12507;
w12509 <= a(41) and not w12508;
w12510 <= not w12507 and not w12508;
w12511 <= not w12509 and not w12510;
w12512 <= not w12500 and not w12511;
w12513 <= not w12500 and not w12512;
w12514 <= not w12511 and not w12512;
w12515 <= not w12513 and not w12514;
w12516 <= not w12160 and not w12163;
w12517 <= w12515 and w12516;
w12518 <= not w12515 and not w12516;
w12519 <= not w12517 and not w12518;
w12520 <= b(25) and w4778;
w12521 <= b(23) and w5020;
w12522 <= b(24) and w4773;
w12523 <= not w12521 and not w12522;
w12524 <= not w12520 and w12523;
w12525 <= w2228 and w4781;
w12526 <= w12524 and not w12525;
w12527 <= a(38) and not w12526;
w12528 <= a(38) and not w12527;
w12529 <= not w12526 and not w12527;
w12530 <= not w12528 and not w12529;
w12531 <= w12519 and not w12530;
w12532 <= w12519 and not w12531;
w12533 <= not w12530 and not w12531;
w12534 <= not w12532 and not w12533;
w12535 <= not w12177 and not w12183;
w12536 <= w12534 and w12535;
w12537 <= not w12534 and not w12535;
w12538 <= not w12536 and not w12537;
w12539 <= b(28) and w4030;
w12540 <= b(26) and w4275;
w12541 <= b(27) and w4025;
w12542 <= not w12540 and not w12541;
w12543 <= not w12539 and w12542;
w12544 <= w2932 and w4033;
w12545 <= w12543 and not w12544;
w12546 <= a(35) and not w12545;
w12547 <= a(35) and not w12546;
w12548 <= not w12545 and not w12546;
w12549 <= not w12547 and not w12548;
w12550 <= w12538 and not w12549;
w12551 <= w12538 and not w12550;
w12552 <= not w12549 and not w12550;
w12553 <= not w12551 and not w12552;
w12554 <= not w12196 and not w12202;
w12555 <= w12553 and w12554;
w12556 <= not w12553 and not w12554;
w12557 <= not w12555 and not w12556;
w12558 <= b(31) and w3381;
w12559 <= b(29) and w3586;
w12560 <= b(30) and w3376;
w12561 <= not w12559 and not w12560;
w12562 <= not w12558 and w12561;
w12563 <= w3384 and w3539;
w12564 <= w12562 and not w12563;
w12565 <= a(32) and not w12564;
w12566 <= a(32) and not w12565;
w12567 <= not w12564 and not w12565;
w12568 <= not w12566 and not w12567;
w12569 <= w12557 and not w12568;
w12570 <= w12557 and not w12569;
w12571 <= not w12568 and not w12569;
w12572 <= not w12570 and not w12571;
w12573 <= not w12362 and w12572;
w12574 <= w12362 and not w12572;
w12575 <= not w12573 and not w12574;
w12576 <= b(34) and w2793;
w12577 <= b(32) and w2986;
w12578 <= b(33) and w2788;
w12579 <= not w12577 and not w12578;
w12580 <= not w12576 and w12579;
w12581 <= w2796 and w4209;
w12582 <= w12580 and not w12581;
w12583 <= a(29) and not w12582;
w12584 <= a(29) and not w12583;
w12585 <= not w12582 and not w12583;
w12586 <= not w12584 and not w12585;
w12587 <= not w12575 and not w12586;
w12588 <= w12575 and w12586;
w12589 <= not w12587 and not w12588;
w12590 <= w12361 and not w12589;
w12591 <= not w12361 and w12589;
w12592 <= not w12590 and not w12591;
w12593 <= b(37) and w2282;
w12594 <= b(35) and w2428;
w12595 <= b(36) and w2277;
w12596 <= not w12594 and not w12595;
w12597 <= not w12593 and w12596;
w12598 <= w2285 and w4924;
w12599 <= w12597 and not w12598;
w12600 <= a(26) and not w12599;
w12601 <= a(26) and not w12600;
w12602 <= not w12599 and not w12600;
w12603 <= not w12601 and not w12602;
w12604 <= w12592 and not w12603;
w12605 <= w12592 and not w12604;
w12606 <= not w12603 and not w12604;
w12607 <= not w12605 and not w12606;
w12608 <= not w12239 and not w12243;
w12609 <= w12607 and w12608;
w12610 <= not w12607 and not w12608;
w12611 <= not w12609 and not w12610;
w12612 <= b(40) and w1791;
w12613 <= b(38) and w1941;
w12614 <= b(39) and w1786;
w12615 <= not w12613 and not w12614;
w12616 <= not w12612 and w12615;
w12617 <= w1794 and w5698;
w12618 <= w12616 and not w12617;
w12619 <= a(23) and not w12618;
w12620 <= a(23) and not w12619;
w12621 <= not w12618 and not w12619;
w12622 <= not w12620 and not w12621;
w12623 <= w12611 and not w12622;
w12624 <= w12611 and not w12623;
w12625 <= not w12622 and not w12623;
w12626 <= not w12624 and not w12625;
w12627 <= not w12256 and not w12262;
w12628 <= w12626 and w12627;
w12629 <= not w12626 and not w12627;
w12630 <= not w12628 and not w12629;
w12631 <= b(43) and w1370;
w12632 <= b(41) and w1506;
w12633 <= b(42) and w1365;
w12634 <= not w12632 and not w12633;
w12635 <= not w12631 and w12634;
w12636 <= w1373 and w6258;
w12637 <= w12635 and not w12636;
w12638 <= a(20) and not w12637;
w12639 <= a(20) and not w12638;
w12640 <= not w12637 and not w12638;
w12641 <= not w12639 and not w12640;
w12642 <= w12630 and not w12641;
w12643 <= not w12630 and w12641;
w12644 <= not w12359 and not w12643;
w12645 <= not w12642 and w12644;
w12646 <= not w12359 and not w12645;
w12647 <= not w12642 and not w12645;
w12648 <= not w12643 and w12647;
w12649 <= not w12646 and not w12648;
w12650 <= b(46) and w1045;
w12651 <= b(44) and w1134;
w12652 <= b(45) and w1040;
w12653 <= not w12651 and not w12652;
w12654 <= not w12650 and w12653;
w12655 <= w1048 and w7420;
w12656 <= w12654 and not w12655;
w12657 <= a(17) and not w12656;
w12658 <= a(17) and not w12657;
w12659 <= not w12656 and not w12657;
w12660 <= not w12658 and not w12659;
w12661 <= w12649 and w12660;
w12662 <= not w12649 and not w12660;
w12663 <= not w12661 and not w12662;
w12664 <= not w12358 and w12663;
w12665 <= w12358 and not w12663;
w12666 <= not w12664 and not w12665;
w12667 <= w12357 and not w12666;
w12668 <= not w12357 and w12666;
w12669 <= not w12667 and not w12668;
w12670 <= not w12346 and w12669;
w12671 <= w12346 and not w12669;
w12672 <= not w12670 and not w12671;
w12673 <= w12345 and not w12672;
w12674 <= not w12345 and w12672;
w12675 <= not w12673 and not w12674;
w12676 <= not w12334 and w12675;
w12677 <= w12334 and not w12675;
w12678 <= not w12676 and not w12677;
w12679 <= not w12333 and w12678;
w12680 <= w12678 and not w12679;
w12681 <= not w12333 and not w12679;
w12682 <= not w12680 and not w12681;
w12683 <= not w12305 and not w12308;
w12684 <= w12682 and w12683;
w12685 <= not w12682 and not w12683;
w12686 <= not w12684 and not w12685;
w12687 <= b(58) and w105;
w12688 <= b(56) and w146;
w12689 <= b(57) and w100;
w12690 <= not w12688 and not w12689;
w12691 <= not w12687 and w12690;
w12692 <= w108 and w11179;
w12693 <= w12691 and not w12692;
w12694 <= a(5) and not w12693;
w12695 <= a(5) and not w12694;
w12696 <= not w12693 and not w12694;
w12697 <= not w12695 and not w12696;
w12698 <= not w12686 and w12697;
w12699 <= w12686 and not w12697;
w12700 <= not w12698 and not w12699;
w12701 <= b(61) and w9;
w12702 <= b(59) and w27;
w12703 <= b(60) and w4;
w12704 <= not w12702 and not w12703;
w12705 <= not w12701 and w12704;
w12706 <= not w11950 and not w11952;
w12707 <= not b(60) and not b(61);
w12708 <= b(60) and b(61);
w12709 <= not w12707 and not w12708;
w12710 <= not w12706 and w12709;
w12711 <= w12706 and not w12709;
w12712 <= not w12710 and not w12711;
w12713 <= w12 and w12712;
w12714 <= w12705 and not w12713;
w12715 <= a(2) and not w12714;
w12716 <= a(2) and not w12715;
w12717 <= not w12714 and not w12715;
w12718 <= not w12716 and not w12717;
w12719 <= w12700 and not w12718;
w12720 <= w12700 and not w12719;
w12721 <= not w12718 and not w12719;
w12722 <= not w12720 and not w12721;
w12723 <= not w12311 and not w12314;
w12724 <= w12722 and w12723;
w12725 <= not w12722 and not w12723;
w12726 <= not w12724 and not w12725;
w12727 <= not w12317 and not w12320;
w12728 <= w12726 and not w12727;
w12729 <= not w12726 and w12727;
w12730 <= not w12728 and not w12729;
w12731 <= not w12725 and not w12728;
w12732 <= not w12699 and not w12719;
w12733 <= not w12674 and not w12676;
w12734 <= not w12668 and not w12670;
w12735 <= b(50) and w694;
w12736 <= b(48) and w799;
w12737 <= b(49) and w689;
w12738 <= not w12736 and not w12737;
w12739 <= not w12735 and w12738;
w12740 <= w697 and w8692;
w12741 <= w12739 and not w12740;
w12742 <= a(14) and not w12741;
w12743 <= a(14) and not w12742;
w12744 <= not w12741 and not w12742;
w12745 <= not w12743 and not w12744;
w12746 <= not w12662 and not w12664;
w12747 <= not w12623 and not w12629;
w12748 <= not w12362 and not w12572;
w12749 <= not w12569 and not w12748;
w12750 <= not w12512 and not w12518;
w12751 <= not w12474 and not w12480;
w12752 <= b(17) and w7189;
w12753 <= b(15) and w7530;
w12754 <= b(16) and w7184;
w12755 <= not w12753 and not w12754;
w12756 <= not w12752 and w12755;
w12757 <= w1099 and w7192;
w12758 <= w12756 and not w12757;
w12759 <= a(47) and not w12758;
w12760 <= a(47) and not w12759;
w12761 <= not w12758 and not w12759;
w12762 <= not w12760 and not w12761;
w12763 <= b(14) and w8105;
w12764 <= b(12) and w8458;
w12765 <= b(13) and w8100;
w12766 <= not w12764 and not w12765;
w12767 <= not w12763 and w12766;
w12768 <= w777 and w8108;
w12769 <= w12767 and not w12768;
w12770 <= a(50) and not w12769;
w12771 <= a(50) and not w12770;
w12772 <= not w12769 and not w12770;
w12773 <= not w12771 and not w12772;
w12774 <= not w12436 and not w12442;
w12775 <= b(11) and w9082;
w12776 <= b(9) and w9475;
w12777 <= b(10) and w9077;
w12778 <= not w12776 and not w12777;
w12779 <= not w12775 and w12778;
w12780 <= w561 and w9085;
w12781 <= w12779 and not w12780;
w12782 <= a(53) and not w12781;
w12783 <= a(53) and not w12782;
w12784 <= not w12781 and not w12782;
w12785 <= not w12783 and not w12784;
w12786 <= not w12431 and not w12433;
w12787 <= not w12425 and not w12427;
w12788 <= b(2) and w12411;
w12789 <= w12097 and not w12410;
w12790 <= w12405 and w12789;
w12791 <= b(0) and w12790;
w12792 <= b(1) and w12406;
w12793 <= not w12791 and not w12792;
w12794 <= not w12788 and w12793;
w12795 <= w39 and w12414;
w12796 <= w12794 and not w12795;
w12797 <= a(62) and not w12796;
w12798 <= a(62) and not w12797;
w12799 <= not w12796 and not w12797;
w12800 <= not w12798 and not w12799;
w12801 <= not w12421 and w12800;
w12802 <= w12421 and not w12800;
w12803 <= not w12801 and not w12802;
w12804 <= b(5) and w11274;
w12805 <= b(3) and w11639;
w12806 <= b(4) and w11269;
w12807 <= not w12805 and not w12806;
w12808 <= not w12804 and w12807;
w12809 <= w137 and w11277;
w12810 <= w12808 and not w12809;
w12811 <= a(59) and not w12810;
w12812 <= a(59) and not w12811;
w12813 <= not w12810 and not w12811;
w12814 <= not w12812 and not w12813;
w12815 <= w12803 and not w12814;
w12816 <= not w12803 and w12814;
w12817 <= not w12787 and not w12816;
w12818 <= not w12815 and w12817;
w12819 <= not w12787 and not w12818;
w12820 <= not w12815 and not w12818;
w12821 <= not w12816 and w12820;
w12822 <= not w12819 and not w12821;
w12823 <= b(8) and w10169;
w12824 <= b(6) and w10539;
w12825 <= b(7) and w10164;
w12826 <= not w12824 and not w12825;
w12827 <= not w12823 and w12826;
w12828 <= w328 and w10172;
w12829 <= w12827 and not w12828;
w12830 <= a(56) and not w12829;
w12831 <= a(56) and not w12830;
w12832 <= not w12829 and not w12830;
w12833 <= not w12831 and not w12832;
w12834 <= w12822 and w12833;
w12835 <= not w12822 and not w12833;
w12836 <= not w12834 and not w12835;
w12837 <= not w12786 and w12836;
w12838 <= w12786 and not w12836;
w12839 <= not w12837 and not w12838;
w12840 <= w12785 and not w12839;
w12841 <= not w12785 and w12839;
w12842 <= not w12840 and not w12841;
w12843 <= not w12774 and w12842;
w12844 <= w12774 and not w12842;
w12845 <= not w12843 and not w12844;
w12846 <= not w12773 and w12845;
w12847 <= w12845 and not w12846;
w12848 <= not w12773 and not w12846;
w12849 <= not w12847 and not w12848;
w12850 <= not w12460 and not w12849;
w12851 <= w12460 and w12849;
w12852 <= not w12850 and not w12851;
w12853 <= not w12762 and w12852;
w12854 <= not w12762 and not w12853;
w12855 <= w12852 and not w12853;
w12856 <= not w12854 and not w12855;
w12857 <= not w12751 and not w12856;
w12858 <= not w12751 and not w12857;
w12859 <= not w12856 and not w12857;
w12860 <= not w12858 and not w12859;
w12861 <= b(20) and w6338;
w12862 <= b(18) and w6645;
w12863 <= b(19) and w6333;
w12864 <= not w12862 and not w12863;
w12865 <= not w12861 and w12864;
w12866 <= w1589 and w6341;
w12867 <= w12865 and not w12866;
w12868 <= a(44) and not w12867;
w12869 <= a(44) and not w12868;
w12870 <= not w12867 and not w12868;
w12871 <= not w12869 and not w12870;
w12872 <= not w12860 and not w12871;
w12873 <= not w12860 and not w12872;
w12874 <= not w12871 and not w12872;
w12875 <= not w12873 and not w12874;
w12876 <= not w12498 and w12875;
w12877 <= w12498 and not w12875;
w12878 <= not w12876 and not w12877;
w12879 <= b(23) and w5520;
w12880 <= b(21) and w5802;
w12881 <= b(22) and w5515;
w12882 <= not w12880 and not w12881;
w12883 <= not w12879 and w12882;
w12884 <= w2043 and w5523;
w12885 <= w12883 and not w12884;
w12886 <= a(41) and not w12885;
w12887 <= a(41) and not w12886;
w12888 <= not w12885 and not w12886;
w12889 <= not w12887 and not w12888;
w12890 <= not w12878 and not w12889;
w12891 <= w12878 and w12889;
w12892 <= not w12890 and not w12891;
w12893 <= w12750 and not w12892;
w12894 <= not w12750 and w12892;
w12895 <= not w12893 and not w12894;
w12896 <= b(26) and w4778;
w12897 <= b(24) and w5020;
w12898 <= b(25) and w4773;
w12899 <= not w12897 and not w12898;
w12900 <= not w12896 and w12899;
w12901 <= w2556 and w4781;
w12902 <= w12900 and not w12901;
w12903 <= a(38) and not w12902;
w12904 <= a(38) and not w12903;
w12905 <= not w12902 and not w12903;
w12906 <= not w12904 and not w12905;
w12907 <= w12895 and not w12906;
w12908 <= w12895 and not w12907;
w12909 <= not w12906 and not w12907;
w12910 <= not w12908 and not w12909;
w12911 <= not w12531 and not w12537;
w12912 <= w12910 and w12911;
w12913 <= not w12910 and not w12911;
w12914 <= not w12912 and not w12913;
w12915 <= b(29) and w4030;
w12916 <= b(27) and w4275;
w12917 <= b(28) and w4025;
w12918 <= not w12916 and not w12917;
w12919 <= not w12915 and w12918;
w12920 <= w3126 and w4033;
w12921 <= w12919 and not w12920;
w12922 <= a(35) and not w12921;
w12923 <= a(35) and not w12922;
w12924 <= not w12921 and not w12922;
w12925 <= not w12923 and not w12924;
w12926 <= w12914 and not w12925;
w12927 <= w12914 and not w12926;
w12928 <= not w12925 and not w12926;
w12929 <= not w12927 and not w12928;
w12930 <= not w12550 and not w12556;
w12931 <= w12929 and w12930;
w12932 <= not w12929 and not w12930;
w12933 <= not w12931 and not w12932;
w12934 <= b(32) and w3381;
w12935 <= b(30) and w3586;
w12936 <= b(31) and w3376;
w12937 <= not w12935 and not w12936;
w12938 <= not w12934 and w12937;
w12939 <= w3384 and w3756;
w12940 <= w12938 and not w12939;
w12941 <= a(32) and not w12940;
w12942 <= a(32) and not w12941;
w12943 <= not w12940 and not w12941;
w12944 <= not w12942 and not w12943;
w12945 <= w12933 and not w12944;
w12946 <= not w12933 and w12944;
w12947 <= not w12749 and not w12946;
w12948 <= not w12945 and w12947;
w12949 <= not w12749 and not w12948;
w12950 <= not w12945 and not w12948;
w12951 <= not w12946 and w12950;
w12952 <= not w12949 and not w12951;
w12953 <= b(35) and w2793;
w12954 <= b(33) and w2986;
w12955 <= b(34) and w2788;
w12956 <= not w12954 and not w12955;
w12957 <= not w12953 and w12956;
w12958 <= w2796 and w4439;
w12959 <= w12957 and not w12958;
w12960 <= a(29) and not w12959;
w12961 <= a(29) and not w12960;
w12962 <= not w12959 and not w12960;
w12963 <= not w12961 and not w12962;
w12964 <= not w12952 and not w12963;
w12965 <= not w12952 and not w12964;
w12966 <= not w12963 and not w12964;
w12967 <= not w12965 and not w12966;
w12968 <= not w12587 and not w12591;
w12969 <= w12967 and w12968;
w12970 <= not w12967 and not w12968;
w12971 <= not w12969 and not w12970;
w12972 <= b(38) and w2282;
w12973 <= b(36) and w2428;
w12974 <= b(37) and w2277;
w12975 <= not w12973 and not w12974;
w12976 <= not w12972 and w12975;
w12977 <= w2285 and w4948;
w12978 <= w12976 and not w12977;
w12979 <= a(26) and not w12978;
w12980 <= a(26) and not w12979;
w12981 <= not w12978 and not w12979;
w12982 <= not w12980 and not w12981;
w12983 <= w12971 and not w12982;
w12984 <= w12971 and not w12983;
w12985 <= not w12982 and not w12983;
w12986 <= not w12984 and not w12985;
w12987 <= not w12604 and not w12610;
w12988 <= w12986 and w12987;
w12989 <= not w12986 and not w12987;
w12990 <= not w12988 and not w12989;
w12991 <= b(41) and w1791;
w12992 <= b(39) and w1941;
w12993 <= b(40) and w1786;
w12994 <= not w12992 and not w12993;
w12995 <= not w12991 and w12994;
w12996 <= w1794 and w5962;
w12997 <= w12995 and not w12996;
w12998 <= a(23) and not w12997;
w12999 <= a(23) and not w12998;
w13000 <= not w12997 and not w12998;
w13001 <= not w12999 and not w13000;
w13002 <= w12990 and not w13001;
w13003 <= not w12990 and w13001;
w13004 <= not w12747 and not w13003;
w13005 <= not w13002 and w13004;
w13006 <= not w12747 and not w13005;
w13007 <= not w13002 and not w13005;
w13008 <= not w13003 and w13007;
w13009 <= not w13006 and not w13008;
w13010 <= b(44) and w1370;
w13011 <= b(42) and w1506;
w13012 <= b(43) and w1365;
w13013 <= not w13011 and not w13012;
w13014 <= not w13010 and w13013;
w13015 <= w1373 and w6815;
w13016 <= w13014 and not w13015;
w13017 <= a(20) and not w13016;
w13018 <= a(20) and not w13017;
w13019 <= not w13016 and not w13017;
w13020 <= not w13018 and not w13019;
w13021 <= not w13009 and not w13020;
w13022 <= not w13009 and not w13021;
w13023 <= not w13020 and not w13021;
w13024 <= not w13022 and not w13023;
w13025 <= not w12647 and w13024;
w13026 <= w12647 and not w13024;
w13027 <= not w13025 and not w13026;
w13028 <= b(47) and w1045;
w13029 <= b(45) and w1134;
w13030 <= b(46) and w1040;
w13031 <= not w13029 and not w13030;
w13032 <= not w13028 and w13031;
w13033 <= w1048 and w7446;
w13034 <= w13032 and not w13033;
w13035 <= a(17) and not w13034;
w13036 <= a(17) and not w13035;
w13037 <= not w13034 and not w13035;
w13038 <= not w13036 and not w13037;
w13039 <= not w13027 and not w13038;
w13040 <= w13027 and w13038;
w13041 <= not w13039 and not w13040;
w13042 <= not w12746 and w13041;
w13043 <= w12746 and not w13041;
w13044 <= not w13042 and not w13043;
w13045 <= not w12745 and w13044;
w13046 <= w13044 and not w13045;
w13047 <= not w12745 and not w13045;
w13048 <= not w13046 and not w13047;
w13049 <= not w12734 and w13048;
w13050 <= w12734 and not w13048;
w13051 <= not w13049 and not w13050;
w13052 <= b(53) and w443;
w13053 <= b(51) and w510;
w13054 <= b(52) and w438;
w13055 <= not w13053 and not w13054;
w13056 <= not w13052 and w13055;
w13057 <= w446 and w9715;
w13058 <= w13056 and not w13057;
w13059 <= a(11) and not w13058;
w13060 <= a(11) and not w13059;
w13061 <= not w13058 and not w13059;
w13062 <= not w13060 and not w13061;
w13063 <= not w13051 and not w13062;
w13064 <= w13051 and w13062;
w13065 <= not w13063 and not w13064;
w13066 <= not w12733 and w13065;
w13067 <= w12733 and not w13065;
w13068 <= not w13066 and not w13067;
w13069 <= b(56) and w254;
w13070 <= b(54) and w284;
w13071 <= b(55) and w249;
w13072 <= not w13070 and not w13071;
w13073 <= not w13069 and w13072;
w13074 <= w257 and w10451;
w13075 <= w13073 and not w13074;
w13076 <= a(8) and not w13075;
w13077 <= a(8) and not w13076;
w13078 <= not w13075 and not w13076;
w13079 <= not w13077 and not w13078;
w13080 <= not w13068 and w13079;
w13081 <= w13068 and not w13079;
w13082 <= not w13080 and not w13081;
w13083 <= b(59) and w105;
w13084 <= b(57) and w146;
w13085 <= b(58) and w100;
w13086 <= not w13084 and not w13085;
w13087 <= not w13083 and w13086;
w13088 <= w108 and w11922;
w13089 <= w13087 and not w13088;
w13090 <= a(5) and not w13089;
w13091 <= a(5) and not w13090;
w13092 <= not w13089 and not w13090;
w13093 <= not w13091 and not w13092;
w13094 <= w13082 and not w13093;
w13095 <= w13082 and not w13094;
w13096 <= not w13093 and not w13094;
w13097 <= not w13095 and not w13096;
w13098 <= not w12679 and not w12685;
w13099 <= w13097 and w13098;
w13100 <= not w13097 and not w13098;
w13101 <= not w13099 and not w13100;
w13102 <= b(62) and w9;
w13103 <= b(60) and w27;
w13104 <= b(61) and w4;
w13105 <= not w13103 and not w13104;
w13106 <= not w13102 and w13105;
w13107 <= not w12708 and not w12710;
w13108 <= not b(61) and not b(62);
w13109 <= b(61) and b(62);
w13110 <= not w13108 and not w13109;
w13111 <= not w13107 and w13110;
w13112 <= w13107 and not w13110;
w13113 <= not w13111 and not w13112;
w13114 <= w12 and w13113;
w13115 <= w13106 and not w13114;
w13116 <= a(2) and not w13115;
w13117 <= a(2) and not w13116;
w13118 <= not w13115 and not w13116;
w13119 <= not w13117 and not w13118;
w13120 <= not w13101 and w13119;
w13121 <= w13101 and not w13119;
w13122 <= not w13120 and not w13121;
w13123 <= not w12732 and w13122;
w13124 <= w12732 and not w13122;
w13125 <= not w13123 and not w13124;
w13126 <= not w12731 and w13125;
w13127 <= w12731 and not w13125;
w13128 <= not w13126 and not w13127;
w13129 <= not w12734 and not w13048;
w13130 <= not w13045 and not w13129;
w13131 <= b(51) and w694;
w13132 <= b(49) and w799;
w13133 <= b(50) and w689;
w13134 <= not w13132 and not w13133;
w13135 <= not w13131 and w13134;
w13136 <= w697 and w8719;
w13137 <= w13135 and not w13136;
w13138 <= a(14) and not w13137;
w13139 <= a(14) and not w13138;
w13140 <= not w13137 and not w13138;
w13141 <= not w13139 and not w13140;
w13142 <= not w13039 and not w13042;
w13143 <= b(48) and w1045;
w13144 <= b(46) and w1134;
w13145 <= b(47) and w1040;
w13146 <= not w13144 and not w13145;
w13147 <= not w13143 and w13146;
w13148 <= w1048 and w7752;
w13149 <= w13147 and not w13148;
w13150 <= a(17) and not w13149;
w13151 <= a(17) and not w13150;
w13152 <= not w13149 and not w13150;
w13153 <= not w13151 and not w13152;
w13154 <= not w12647 and not w13024;
w13155 <= not w13021 and not w13154;
w13156 <= b(45) and w1370;
w13157 <= b(43) and w1506;
w13158 <= b(44) and w1365;
w13159 <= not w13157 and not w13158;
w13160 <= not w13156 and w13159;
w13161 <= w1373 and w7104;
w13162 <= w13160 and not w13161;
w13163 <= a(20) and not w13162;
w13164 <= a(20) and not w13163;
w13165 <= not w13162 and not w13163;
w13166 <= not w13164 and not w13165;
w13167 <= b(42) and w1791;
w13168 <= b(40) and w1941;
w13169 <= b(41) and w1786;
w13170 <= not w13168 and not w13169;
w13171 <= not w13167 and w13170;
w13172 <= w1794 and w6232;
w13173 <= w13171 and not w13172;
w13174 <= a(23) and not w13173;
w13175 <= a(23) and not w13174;
w13176 <= not w13173 and not w13174;
w13177 <= not w13175 and not w13176;
w13178 <= not w12983 and not w12989;
w13179 <= not w12964 and not w12970;
w13180 <= b(33) and w3381;
w13181 <= b(31) and w3586;
w13182 <= b(32) and w3376;
w13183 <= not w13181 and not w13182;
w13184 <= not w13180 and w13183;
w13185 <= w3384 and w3966;
w13186 <= w13184 and not w13185;
w13187 <= a(32) and not w13186;
w13188 <= a(32) and not w13187;
w13189 <= not w13186 and not w13187;
w13190 <= not w13188 and not w13189;
w13191 <= not w12498 and not w12875;
w13192 <= not w12872 and not w13191;
w13193 <= b(21) and w6338;
w13194 <= b(19) and w6645;
w13195 <= b(20) and w6333;
w13196 <= not w13194 and not w13195;
w13197 <= not w13193 and w13196;
w13198 <= w1727 and w6341;
w13199 <= w13197 and not w13198;
w13200 <= a(44) and not w13199;
w13201 <= a(44) and not w13200;
w13202 <= not w13199 and not w13200;
w13203 <= not w13201 and not w13202;
w13204 <= not w12853 and not w12857;
w13205 <= b(15) and w8105;
w13206 <= b(13) and w8458;
w13207 <= b(14) and w8100;
w13208 <= not w13206 and not w13207;
w13209 <= not w13205 and w13208;
w13210 <= w874 and w8108;
w13211 <= w13209 and not w13210;
w13212 <= a(50) and not w13211;
w13213 <= a(50) and not w13212;
w13214 <= not w13211 and not w13212;
w13215 <= not w13213 and not w13214;
w13216 <= not w12841 and not w12843;
w13217 <= not w12835 and not w12837;
w13218 <= b(9) and w10169;
w13219 <= b(7) and w10539;
w13220 <= b(8) and w10164;
w13221 <= not w13219 and not w13220;
w13222 <= not w13218 and w13221;
w13223 <= w394 and w10172;
w13224 <= w13222 and not w13223;
w13225 <= a(56) and not w13224;
w13226 <= a(56) and not w13225;
w13227 <= not w13224 and not w13225;
w13228 <= not w13226 and not w13227;
w13229 <= a(62) and not a(63);
w13230 <= not a(62) and a(63);
w13231 <= not w13229 and not w13230;
w13232 <= b(0) and not w13231;
w13233 <= w12802 and w13232;
w13234 <= w12802 and not w13233;
w13235 <= w13232 and not w13233;
w13236 <= not w13234 and not w13235;
w13237 <= b(3) and w12411;
w13238 <= b(1) and w12790;
w13239 <= b(2) and w12406;
w13240 <= not w13238 and not w13239;
w13241 <= not w13237 and w13240;
w13242 <= w61 and w12414;
w13243 <= w13241 and not w13242;
w13244 <= a(62) and not w13243;
w13245 <= a(62) and not w13244;
w13246 <= not w13243 and not w13244;
w13247 <= not w13245 and not w13246;
w13248 <= not w13236 and not w13247;
w13249 <= not w13236 and not w13248;
w13250 <= not w13247 and not w13248;
w13251 <= not w13249 and not w13250;
w13252 <= b(6) and w11274;
w13253 <= b(4) and w11639;
w13254 <= b(5) and w11269;
w13255 <= not w13253 and not w13254;
w13256 <= not w13252 and w13255;
w13257 <= w202 and w11277;
w13258 <= w13256 and not w13257;
w13259 <= a(59) and not w13258;
w13260 <= a(59) and not w13259;
w13261 <= not w13258 and not w13259;
w13262 <= not w13260 and not w13261;
w13263 <= w13251 and w13262;
w13264 <= not w13251 and not w13262;
w13265 <= not w13263 and not w13264;
w13266 <= not w12820 and w13265;
w13267 <= w12820 and not w13265;
w13268 <= not w13266 and not w13267;
w13269 <= not w13228 and w13268;
w13270 <= w13268 and not w13269;
w13271 <= not w13228 and not w13269;
w13272 <= not w13270 and not w13271;
w13273 <= not w13217 and w13272;
w13274 <= w13217 and not w13272;
w13275 <= not w13273 and not w13274;
w13276 <= b(12) and w9082;
w13277 <= b(10) and w9475;
w13278 <= b(11) and w9077;
w13279 <= not w13277 and not w13278;
w13280 <= not w13276 and w13279;
w13281 <= w585 and w9085;
w13282 <= w13280 and not w13281;
w13283 <= a(53) and not w13282;
w13284 <= a(53) and not w13283;
w13285 <= not w13282 and not w13283;
w13286 <= not w13284 and not w13285;
w13287 <= w13275 and w13286;
w13288 <= not w13275 and not w13286;
w13289 <= not w13287 and not w13288;
w13290 <= not w13216 and w13289;
w13291 <= w13216 and not w13289;
w13292 <= not w13290 and not w13291;
w13293 <= not w13215 and w13292;
w13294 <= w13292 and not w13293;
w13295 <= not w13215 and not w13293;
w13296 <= not w13294 and not w13295;
w13297 <= not w12846 and not w12850;
w13298 <= w13296 and w13297;
w13299 <= not w13296 and not w13297;
w13300 <= not w13298 and not w13299;
w13301 <= b(18) and w7189;
w13302 <= b(16) and w7530;
w13303 <= b(17) and w7184;
w13304 <= not w13302 and not w13303;
w13305 <= not w13301 and w13304;
w13306 <= w1309 and w7192;
w13307 <= w13305 and not w13306;
w13308 <= a(47) and not w13307;
w13309 <= a(47) and not w13308;
w13310 <= not w13307 and not w13308;
w13311 <= not w13309 and not w13310;
w13312 <= not w13300 and w13311;
w13313 <= w13300 and not w13311;
w13314 <= not w13312 and not w13313;
w13315 <= not w13204 and w13314;
w13316 <= w13204 and not w13314;
w13317 <= not w13315 and not w13316;
w13318 <= not w13203 and w13317;
w13319 <= w13203 and not w13317;
w13320 <= not w13318 and not w13319;
w13321 <= not w13192 and w13320;
w13322 <= w13192 and not w13320;
w13323 <= not w13321 and not w13322;
w13324 <= b(24) and w5520;
w13325 <= b(22) and w5802;
w13326 <= b(23) and w5515;
w13327 <= not w13325 and not w13326;
w13328 <= not w13324 and w13327;
w13329 <= w2201 and w5523;
w13330 <= w13328 and not w13329;
w13331 <= a(41) and not w13330;
w13332 <= a(41) and not w13331;
w13333 <= not w13330 and not w13331;
w13334 <= not w13332 and not w13333;
w13335 <= w13323 and not w13334;
w13336 <= w13323 and not w13335;
w13337 <= not w13334 and not w13335;
w13338 <= not w13336 and not w13337;
w13339 <= not w12890 and not w12894;
w13340 <= w13338 and w13339;
w13341 <= not w13338 and not w13339;
w13342 <= not w13340 and not w13341;
w13343 <= b(27) and w4778;
w13344 <= b(25) and w5020;
w13345 <= b(26) and w4773;
w13346 <= not w13344 and not w13345;
w13347 <= not w13343 and w13346;
w13348 <= w2733 and w4781;
w13349 <= w13347 and not w13348;
w13350 <= a(38) and not w13349;
w13351 <= a(38) and not w13350;
w13352 <= not w13349 and not w13350;
w13353 <= not w13351 and not w13352;
w13354 <= w13342 and not w13353;
w13355 <= w13342 and not w13354;
w13356 <= not w13353 and not w13354;
w13357 <= not w13355 and not w13356;
w13358 <= not w12907 and not w12913;
w13359 <= w13357 and w13358;
w13360 <= not w13357 and not w13358;
w13361 <= not w13359 and not w13360;
w13362 <= b(30) and w4030;
w13363 <= b(28) and w4275;
w13364 <= b(29) and w4025;
w13365 <= not w13363 and not w13364;
w13366 <= not w13362 and w13365;
w13367 <= w3320 and w4033;
w13368 <= w13366 and not w13367;
w13369 <= a(35) and not w13368;
w13370 <= a(35) and not w13369;
w13371 <= not w13368 and not w13369;
w13372 <= not w13370 and not w13371;
w13373 <= not w13361 and w13372;
w13374 <= w13361 and not w13372;
w13375 <= not w13373 and not w13374;
w13376 <= not w12926 and not w12932;
w13377 <= w13375 and not w13376;
w13378 <= not w13375 and w13376;
w13379 <= not w13377 and not w13378;
w13380 <= not w13190 and w13379;
w13381 <= w13379 and not w13380;
w13382 <= not w13190 and not w13380;
w13383 <= not w13381 and not w13382;
w13384 <= not w12950 and w13383;
w13385 <= w12950 and not w13383;
w13386 <= not w13384 and not w13385;
w13387 <= b(36) and w2793;
w13388 <= b(34) and w2986;
w13389 <= b(35) and w2788;
w13390 <= not w13388 and not w13389;
w13391 <= not w13387 and w13390;
w13392 <= w2796 and w4665;
w13393 <= w13391 and not w13392;
w13394 <= a(29) and not w13393;
w13395 <= a(29) and not w13394;
w13396 <= not w13393 and not w13394;
w13397 <= not w13395 and not w13396;
w13398 <= not w13386 and not w13397;
w13399 <= w13386 and w13397;
w13400 <= not w13398 and not w13399;
w13401 <= w13179 and not w13400;
w13402 <= not w13179 and w13400;
w13403 <= not w13401 and not w13402;
w13404 <= b(39) and w2282;
w13405 <= b(37) and w2428;
w13406 <= b(38) and w2277;
w13407 <= not w13405 and not w13406;
w13408 <= not w13404 and w13407;
w13409 <= w2285 and w5194;
w13410 <= w13408 and not w13409;
w13411 <= a(26) and not w13410;
w13412 <= a(26) and not w13411;
w13413 <= not w13410 and not w13411;
w13414 <= not w13412 and not w13413;
w13415 <= not w13403 and w13414;
w13416 <= w13403 and not w13414;
w13417 <= not w13415 and not w13416;
w13418 <= not w13178 and w13417;
w13419 <= w13178 and not w13417;
w13420 <= not w13418 and not w13419;
w13421 <= not w13177 and w13420;
w13422 <= not w13177 and not w13421;
w13423 <= w13420 and not w13421;
w13424 <= not w13422 and not w13423;
w13425 <= not w13007 and not w13424;
w13426 <= w13007 and not w13423;
w13427 <= not w13422 and w13426;
w13428 <= not w13425 and not w13427;
w13429 <= not w13166 and w13428;
w13430 <= not w13166 and not w13429;
w13431 <= w13428 and not w13429;
w13432 <= not w13430 and not w13431;
w13433 <= not w13155 and not w13432;
w13434 <= w13155 and not w13431;
w13435 <= not w13430 and w13434;
w13436 <= not w13433 and not w13435;
w13437 <= not w13153 and w13436;
w13438 <= not w13153 and not w13437;
w13439 <= w13436 and not w13437;
w13440 <= not w13438 and not w13439;
w13441 <= not w13142 and not w13440;
w13442 <= w13142 and not w13439;
w13443 <= not w13438 and w13442;
w13444 <= not w13441 and not w13443;
w13445 <= not w13141 and w13444;
w13446 <= w13141 and not w13444;
w13447 <= not w13445 and not w13446;
w13448 <= not w13130 and w13447;
w13449 <= w13130 and not w13447;
w13450 <= not w13448 and not w13449;
w13451 <= b(54) and w443;
w13452 <= b(52) and w510;
w13453 <= b(53) and w438;
w13454 <= not w13452 and not w13453;
w13455 <= not w13451 and w13454;
w13456 <= w446 and w9741;
w13457 <= w13455 and not w13456;
w13458 <= a(11) and not w13457;
w13459 <= a(11) and not w13458;
w13460 <= not w13457 and not w13458;
w13461 <= not w13459 and not w13460;
w13462 <= w13450 and not w13461;
w13463 <= w13450 and not w13462;
w13464 <= not w13461 and not w13462;
w13465 <= not w13463 and not w13464;
w13466 <= not w13063 and not w13066;
w13467 <= w13465 and w13466;
w13468 <= not w13465 and not w13466;
w13469 <= not w13467 and not w13468;
w13470 <= b(57) and w254;
w13471 <= b(55) and w284;
w13472 <= b(56) and w249;
w13473 <= not w13471 and not w13472;
w13474 <= not w13470 and w13473;
w13475 <= w257 and w11153;
w13476 <= w13474 and not w13475;
w13477 <= a(8) and not w13476;
w13478 <= a(8) and not w13477;
w13479 <= not w13476 and not w13477;
w13480 <= not w13478 and not w13479;
w13481 <= w13469 and not w13480;
w13482 <= w13469 and not w13481;
w13483 <= not w13480 and not w13481;
w13484 <= not w13482 and not w13483;
w13485 <= b(60) and w105;
w13486 <= b(58) and w146;
w13487 <= b(59) and w100;
w13488 <= not w13486 and not w13487;
w13489 <= not w13485 and w13488;
w13490 <= w108 and w11954;
w13491 <= w13489 and not w13490;
w13492 <= a(5) and not w13491;
w13493 <= a(5) and not w13492;
w13494 <= not w13491 and not w13492;
w13495 <= not w13493 and not w13494;
w13496 <= not w13484 and w13495;
w13497 <= w13484 and not w13495;
w13498 <= not w13496 and not w13497;
w13499 <= not w13081 and not w13094;
w13500 <= w13498 and w13499;
w13501 <= not w13498 and not w13499;
w13502 <= not w13500 and not w13501;
w13503 <= b(63) and w9;
w13504 <= b(61) and w27;
w13505 <= b(62) and w4;
w13506 <= not w13504 and not w13505;
w13507 <= not w13503 and w13506;
w13508 <= not w13109 and not w13111;
w13509 <= b(62) and not b(63);
w13510 <= not b(62) and b(63);
w13511 <= not w13509 and not w13510;
w13512 <= not w13508 and not w13511;
w13513 <= w13508 and w13511;
w13514 <= not w13512 and not w13513;
w13515 <= w12 and w13514;
w13516 <= w13507 and not w13515;
w13517 <= a(2) and not w13516;
w13518 <= a(2) and not w13517;
w13519 <= not w13516 and not w13517;
w13520 <= not w13518 and not w13519;
w13521 <= w13502 and not w13520;
w13522 <= w13502 and not w13521;
w13523 <= not w13520 and not w13521;
w13524 <= not w13522 and not w13523;
w13525 <= not w13100 and not w13121;
w13526 <= not w13524 and not w13525;
w13527 <= not w13524 and not w13526;
w13528 <= not w13525 and not w13526;
w13529 <= not w13527 and not w13528;
w13530 <= not w13123 and not w13126;
w13531 <= not w13529 and not w13530;
w13532 <= w13529 and w13530;
w13533 <= not w13531 and not w13532;
w13534 <= not w13526 and not w13531;
w13535 <= not w13501 and not w13521;
w13536 <= b(62) and w27;
w13537 <= b(63) and w4;
w13538 <= not w13536 and not w13537;
w13539 <= not b(62) and not w13512;
w13540 <= b(63) and not w13539;
w13541 <= b(63) and not w13540;
w13542 <= not w13508 and w13509;
w13543 <= not w13541 and not w13542;
w13544 <= w12 and not w13543;
w13545 <= w13538 and not w13544;
w13546 <= a(2) and not w13545;
w13547 <= a(2) and not w13546;
w13548 <= not w13545 and not w13546;
w13549 <= not w13547 and not w13548;
w13550 <= not w13484 and not w13495;
w13551 <= not w13481 and not w13550;
w13552 <= not w13462 and not w13468;
w13553 <= b(55) and w443;
w13554 <= b(53) and w510;
w13555 <= b(54) and w438;
w13556 <= not w13554 and not w13555;
w13557 <= not w13553 and w13556;
w13558 <= w446 and w10427;
w13559 <= w13557 and not w13558;
w13560 <= a(11) and not w13559;
w13561 <= a(11) and not w13560;
w13562 <= not w13559 and not w13560;
w13563 <= not w13561 and not w13562;
w13564 <= not w13445 and not w13448;
w13565 <= b(52) and w694;
w13566 <= b(50) and w799;
w13567 <= b(51) and w689;
w13568 <= not w13566 and not w13567;
w13569 <= not w13565 and w13568;
w13570 <= w697 and w9371;
w13571 <= w13569 and not w13570;
w13572 <= a(14) and not w13571;
w13573 <= a(14) and not w13572;
w13574 <= not w13571 and not w13572;
w13575 <= not w13573 and not w13574;
w13576 <= not w13437 and not w13441;
w13577 <= b(49) and w1045;
w13578 <= b(47) and w1134;
w13579 <= b(48) and w1040;
w13580 <= not w13578 and not w13579;
w13581 <= not w13577 and w13580;
w13582 <= w1048 and w8368;
w13583 <= w13581 and not w13582;
w13584 <= a(17) and not w13583;
w13585 <= a(17) and not w13584;
w13586 <= not w13583 and not w13584;
w13587 <= not w13585 and not w13586;
w13588 <= not w13429 and not w13433;
w13589 <= b(46) and w1370;
w13590 <= b(44) and w1506;
w13591 <= b(45) and w1365;
w13592 <= not w13590 and not w13591;
w13593 <= not w13589 and w13592;
w13594 <= w1373 and w7420;
w13595 <= w13593 and not w13594;
w13596 <= a(20) and not w13595;
w13597 <= a(20) and not w13596;
w13598 <= not w13595 and not w13596;
w13599 <= not w13597 and not w13598;
w13600 <= not w13421 and not w13425;
w13601 <= b(34) and w3381;
w13602 <= b(32) and w3586;
w13603 <= b(33) and w3376;
w13604 <= not w13602 and not w13603;
w13605 <= not w13601 and w13604;
w13606 <= w3384 and w4209;
w13607 <= w13605 and not w13606;
w13608 <= a(32) and not w13607;
w13609 <= a(32) and not w13608;
w13610 <= not w13607 and not w13608;
w13611 <= not w13609 and not w13610;
w13612 <= b(22) and w6338;
w13613 <= b(20) and w6645;
w13614 <= b(21) and w6333;
w13615 <= not w13613 and not w13614;
w13616 <= not w13612 and w13615;
w13617 <= w1888 and w6341;
w13618 <= w13616 and not w13617;
w13619 <= a(44) and not w13618;
w13620 <= a(44) and not w13619;
w13621 <= not w13618 and not w13619;
w13622 <= not w13620 and not w13621;
w13623 <= b(16) and w8105;
w13624 <= b(14) and w8458;
w13625 <= b(15) and w8100;
w13626 <= not w13624 and not w13625;
w13627 <= not w13623 and w13626;
w13628 <= w980 and w8108;
w13629 <= w13627 and not w13628;
w13630 <= a(50) and not w13629;
w13631 <= a(50) and not w13630;
w13632 <= not w13629 and not w13630;
w13633 <= not w13631 and not w13632;
w13634 <= b(10) and w10169;
w13635 <= b(8) and w10539;
w13636 <= b(9) and w10164;
w13637 <= not w13635 and not w13636;
w13638 <= not w13634 and w13637;
w13639 <= w481 and w10172;
w13640 <= w13638 and not w13639;
w13641 <= a(56) and not w13640;
w13642 <= a(56) and not w13641;
w13643 <= not w13640 and not w13641;
w13644 <= not w13642 and not w13643;
w13645 <= not w13264 and not w13266;
w13646 <= a(63) and w13231;
w13647 <= b(0) and w13646;
w13648 <= b(1) and not w13231;
w13649 <= not w13647 and not w13648;
w13650 <= b(4) and w12411;
w13651 <= b(2) and w12790;
w13652 <= b(3) and w12406;
w13653 <= not w13651 and not w13652;
w13654 <= not w13650 and w13653;
w13655 <= w89 and w12414;
w13656 <= w13654 and not w13655;
w13657 <= a(62) and not w13656;
w13658 <= a(62) and not w13657;
w13659 <= not w13656 and not w13657;
w13660 <= not w13658 and not w13659;
w13661 <= not w13649 and not w13660;
w13662 <= not w13649 and not w13661;
w13663 <= not w13660 and not w13661;
w13664 <= not w13662 and not w13663;
w13665 <= not w13233 and not w13248;
w13666 <= w13664 and w13665;
w13667 <= not w13664 and not w13665;
w13668 <= not w13666 and not w13667;
w13669 <= b(7) and w11274;
w13670 <= b(5) and w11639;
w13671 <= b(6) and w11269;
w13672 <= not w13670 and not w13671;
w13673 <= not w13669 and w13672;
w13674 <= w227 and w11277;
w13675 <= w13673 and not w13674;
w13676 <= a(59) and not w13675;
w13677 <= a(59) and not w13676;
w13678 <= not w13675 and not w13676;
w13679 <= not w13677 and not w13678;
w13680 <= not w13668 and w13679;
w13681 <= w13668 and not w13679;
w13682 <= not w13680 and not w13681;
w13683 <= not w13645 and w13682;
w13684 <= w13645 and not w13682;
w13685 <= not w13683 and not w13684;
w13686 <= not w13644 and w13685;
w13687 <= w13685 and not w13686;
w13688 <= not w13644 and not w13686;
w13689 <= not w13687 and not w13688;
w13690 <= not w13217 and not w13272;
w13691 <= not w13269 and not w13690;
w13692 <= w13689 and w13691;
w13693 <= not w13689 and not w13691;
w13694 <= not w13692 and not w13693;
w13695 <= b(13) and w9082;
w13696 <= b(11) and w9475;
w13697 <= b(12) and w9077;
w13698 <= not w13696 and not w13697;
w13699 <= not w13695 and w13698;
w13700 <= w751 and w9085;
w13701 <= w13699 and not w13700;
w13702 <= a(53) and not w13701;
w13703 <= a(53) and not w13702;
w13704 <= not w13701 and not w13702;
w13705 <= not w13703 and not w13704;
w13706 <= not w13694 and w13705;
w13707 <= w13694 and not w13705;
w13708 <= not w13706 and not w13707;
w13709 <= not w13288 and not w13290;
w13710 <= w13708 and not w13709;
w13711 <= not w13708 and w13709;
w13712 <= not w13710 and not w13711;
w13713 <= not w13633 and w13712;
w13714 <= w13712 and not w13713;
w13715 <= not w13633 and not w13713;
w13716 <= not w13714 and not w13715;
w13717 <= not w13293 and not w13299;
w13718 <= w13716 and w13717;
w13719 <= not w13716 and not w13717;
w13720 <= not w13718 and not w13719;
w13721 <= b(19) and w7189;
w13722 <= b(17) and w7530;
w13723 <= b(18) and w7184;
w13724 <= not w13722 and not w13723;
w13725 <= not w13721 and w13724;
w13726 <= w1451 and w7192;
w13727 <= w13725 and not w13726;
w13728 <= a(47) and not w13727;
w13729 <= a(47) and not w13728;
w13730 <= not w13727 and not w13728;
w13731 <= not w13729 and not w13730;
w13732 <= not w13720 and w13731;
w13733 <= w13720 and not w13731;
w13734 <= not w13732 and not w13733;
w13735 <= not w13313 and not w13315;
w13736 <= w13734 and not w13735;
w13737 <= not w13734 and w13735;
w13738 <= not w13736 and not w13737;
w13739 <= not w13622 and w13738;
w13740 <= w13738 and not w13739;
w13741 <= not w13622 and not w13739;
w13742 <= not w13740 and not w13741;
w13743 <= not w13318 and not w13321;
w13744 <= w13742 and w13743;
w13745 <= not w13742 and not w13743;
w13746 <= not w13744 and not w13745;
w13747 <= b(25) and w5520;
w13748 <= b(23) and w5802;
w13749 <= b(24) and w5515;
w13750 <= not w13748 and not w13749;
w13751 <= not w13747 and w13750;
w13752 <= w2228 and w5523;
w13753 <= w13751 and not w13752;
w13754 <= a(41) and not w13753;
w13755 <= a(41) and not w13754;
w13756 <= not w13753 and not w13754;
w13757 <= not w13755 and not w13756;
w13758 <= w13746 and not w13757;
w13759 <= w13746 and not w13758;
w13760 <= not w13757 and not w13758;
w13761 <= not w13759 and not w13760;
w13762 <= not w13335 and not w13341;
w13763 <= w13761 and w13762;
w13764 <= not w13761 and not w13762;
w13765 <= not w13763 and not w13764;
w13766 <= b(28) and w4778;
w13767 <= b(26) and w5020;
w13768 <= b(27) and w4773;
w13769 <= not w13767 and not w13768;
w13770 <= not w13766 and w13769;
w13771 <= w2932 and w4781;
w13772 <= w13770 and not w13771;
w13773 <= a(38) and not w13772;
w13774 <= a(38) and not w13773;
w13775 <= not w13772 and not w13773;
w13776 <= not w13774 and not w13775;
w13777 <= w13765 and not w13776;
w13778 <= w13765 and not w13777;
w13779 <= not w13776 and not w13777;
w13780 <= not w13778 and not w13779;
w13781 <= not w13354 and not w13360;
w13782 <= w13780 and w13781;
w13783 <= not w13780 and not w13781;
w13784 <= not w13782 and not w13783;
w13785 <= b(31) and w4030;
w13786 <= b(29) and w4275;
w13787 <= b(30) and w4025;
w13788 <= not w13786 and not w13787;
w13789 <= not w13785 and w13788;
w13790 <= w3539 and w4033;
w13791 <= w13789 and not w13790;
w13792 <= a(35) and not w13791;
w13793 <= a(35) and not w13792;
w13794 <= not w13791 and not w13792;
w13795 <= not w13793 and not w13794;
w13796 <= not w13784 and w13795;
w13797 <= w13784 and not w13795;
w13798 <= not w13796 and not w13797;
w13799 <= not w13374 and not w13377;
w13800 <= w13798 and not w13799;
w13801 <= not w13798 and w13799;
w13802 <= not w13800 and not w13801;
w13803 <= not w13611 and w13802;
w13804 <= w13802 and not w13803;
w13805 <= not w13611 and not w13803;
w13806 <= not w13804 and not w13805;
w13807 <= not w12950 and not w13383;
w13808 <= not w13380 and not w13807;
w13809 <= w13806 and w13808;
w13810 <= not w13806 and not w13808;
w13811 <= not w13809 and not w13810;
w13812 <= b(37) and w2793;
w13813 <= b(35) and w2986;
w13814 <= b(36) and w2788;
w13815 <= not w13813 and not w13814;
w13816 <= not w13812 and w13815;
w13817 <= w2796 and w4924;
w13818 <= w13816 and not w13817;
w13819 <= a(29) and not w13818;
w13820 <= a(29) and not w13819;
w13821 <= not w13818 and not w13819;
w13822 <= not w13820 and not w13821;
w13823 <= w13811 and not w13822;
w13824 <= w13811 and not w13823;
w13825 <= not w13822 and not w13823;
w13826 <= not w13824 and not w13825;
w13827 <= not w13398 and not w13402;
w13828 <= w13826 and w13827;
w13829 <= not w13826 and not w13827;
w13830 <= not w13828 and not w13829;
w13831 <= b(40) and w2282;
w13832 <= b(38) and w2428;
w13833 <= b(39) and w2277;
w13834 <= not w13832 and not w13833;
w13835 <= not w13831 and w13834;
w13836 <= w2285 and w5698;
w13837 <= w13835 and not w13836;
w13838 <= a(26) and not w13837;
w13839 <= a(26) and not w13838;
w13840 <= not w13837 and not w13838;
w13841 <= not w13839 and not w13840;
w13842 <= w13830 and not w13841;
w13843 <= w13830 and not w13842;
w13844 <= not w13841 and not w13842;
w13845 <= not w13843 and not w13844;
w13846 <= not w13416 and not w13418;
w13847 <= not w13845 and not w13846;
w13848 <= not w13845 and not w13847;
w13849 <= not w13846 and not w13847;
w13850 <= not w13848 and not w13849;
w13851 <= b(43) and w1791;
w13852 <= b(41) and w1941;
w13853 <= b(42) and w1786;
w13854 <= not w13852 and not w13853;
w13855 <= not w13851 and w13854;
w13856 <= w1794 and w6258;
w13857 <= w13855 and not w13856;
w13858 <= a(23) and not w13857;
w13859 <= a(23) and not w13858;
w13860 <= not w13857 and not w13858;
w13861 <= not w13859 and not w13860;
w13862 <= not w13850 and w13861;
w13863 <= w13850 and not w13861;
w13864 <= not w13862 and not w13863;
w13865 <= not w13600 and not w13864;
w13866 <= w13600 and w13864;
w13867 <= not w13865 and not w13866;
w13868 <= not w13599 and w13867;
w13869 <= not w13599 and not w13868;
w13870 <= w13867 and not w13868;
w13871 <= not w13869 and not w13870;
w13872 <= not w13588 and not w13871;
w13873 <= w13588 and not w13870;
w13874 <= not w13869 and w13873;
w13875 <= not w13872 and not w13874;
w13876 <= not w13587 and w13875;
w13877 <= not w13587 and not w13876;
w13878 <= w13875 and not w13876;
w13879 <= not w13877 and not w13878;
w13880 <= not w13576 and not w13879;
w13881 <= w13576 and not w13878;
w13882 <= not w13877 and w13881;
w13883 <= not w13880 and not w13882;
w13884 <= not w13575 and w13883;
w13885 <= w13575 and not w13883;
w13886 <= not w13884 and not w13885;
w13887 <= not w13564 and w13886;
w13888 <= w13564 and not w13886;
w13889 <= not w13887 and not w13888;
w13890 <= not w13563 and w13889;
w13891 <= w13563 and not w13889;
w13892 <= not w13890 and not w13891;
w13893 <= not w13552 and w13892;
w13894 <= w13552 and not w13892;
w13895 <= not w13893 and not w13894;
w13896 <= b(58) and w254;
w13897 <= b(56) and w284;
w13898 <= b(57) and w249;
w13899 <= not w13897 and not w13898;
w13900 <= not w13896 and w13899;
w13901 <= w257 and w11179;
w13902 <= w13900 and not w13901;
w13903 <= a(8) and not w13902;
w13904 <= a(8) and not w13903;
w13905 <= not w13902 and not w13903;
w13906 <= not w13904 and not w13905;
w13907 <= w13895 and not w13906;
w13908 <= w13895 and not w13907;
w13909 <= not w13906 and not w13907;
w13910 <= not w13908 and not w13909;
w13911 <= b(61) and w105;
w13912 <= b(59) and w146;
w13913 <= b(60) and w100;
w13914 <= not w13912 and not w13913;
w13915 <= not w13911 and w13914;
w13916 <= w108 and w12712;
w13917 <= w13915 and not w13916;
w13918 <= a(5) and not w13917;
w13919 <= a(5) and not w13918;
w13920 <= not w13917 and not w13918;
w13921 <= not w13919 and not w13920;
w13922 <= not w13910 and w13921;
w13923 <= w13910 and not w13921;
w13924 <= not w13922 and not w13923;
w13925 <= not w13551 and not w13924;
w13926 <= w13551 and w13924;
w13927 <= not w13925 and not w13926;
w13928 <= not w13549 and w13927;
w13929 <= w13549 and not w13927;
w13930 <= not w13928 and not w13929;
w13931 <= not w13535 and w13930;
w13932 <= w13535 and not w13930;
w13933 <= not w13931 and not w13932;
w13934 <= not w13534 and w13933;
w13935 <= w13534 and not w13933;
w13936 <= not w13934 and not w13935;
w13937 <= b(53) and w694;
w13938 <= b(51) and w799;
w13939 <= b(52) and w689;
w13940 <= not w13938 and not w13939;
w13941 <= not w13937 and w13940;
w13942 <= w697 and w9715;
w13943 <= w13941 and not w13942;
w13944 <= a(14) and not w13943;
w13945 <= a(14) and not w13944;
w13946 <= not w13943 and not w13944;
w13947 <= not w13945 and not w13946;
w13948 <= not w13876 and not w13880;
w13949 <= not w13868 and not w13872;
w13950 <= b(47) and w1370;
w13951 <= b(45) and w1506;
w13952 <= b(46) and w1365;
w13953 <= not w13951 and not w13952;
w13954 <= not w13950 and w13953;
w13955 <= w1373 and w7446;
w13956 <= w13954 and not w13955;
w13957 <= a(20) and not w13956;
w13958 <= a(20) and not w13957;
w13959 <= not w13956 and not w13957;
w13960 <= not w13958 and not w13959;
w13961 <= not w13842 and not w13847;
w13962 <= not w13797 and not w13800;
w13963 <= not w13739 and not w13745;
w13964 <= not w13733 and not w13736;
w13965 <= not w13713 and not w13719;
w13966 <= not w13707 and not w13710;
w13967 <= b(14) and w9082;
w13968 <= b(12) and w9475;
w13969 <= b(13) and w9077;
w13970 <= not w13968 and not w13969;
w13971 <= not w13967 and w13970;
w13972 <= w777 and w9085;
w13973 <= w13971 and not w13972;
w13974 <= a(53) and not w13973;
w13975 <= a(53) and not w13974;
w13976 <= not w13973 and not w13974;
w13977 <= not w13975 and not w13976;
w13978 <= not w13686 and not w13693;
w13979 <= not w13681 and not w13683;
w13980 <= b(1) and w13646;
w13981 <= b(2) and not w13231;
w13982 <= not w13980 and not w13981;
w13983 <= b(5) and w12411;
w13984 <= b(3) and w12790;
w13985 <= b(4) and w12406;
w13986 <= not w13984 and not w13985;
w13987 <= not w13983 and w13986;
w13988 <= w137 and w12414;
w13989 <= w13987 and not w13988;
w13990 <= a(62) and not w13989;
w13991 <= a(62) and not w13990;
w13992 <= not w13989 and not w13990;
w13993 <= not w13991 and not w13992;
w13994 <= not w13982 and not w13993;
w13995 <= not w13982 and not w13994;
w13996 <= not w13993 and not w13994;
w13997 <= not w13995 and not w13996;
w13998 <= not w13661 and not w13667;
w13999 <= w13997 and w13998;
w14000 <= not w13997 and not w13998;
w14001 <= not w13999 and not w14000;
w14002 <= b(8) and w11274;
w14003 <= b(6) and w11639;
w14004 <= b(7) and w11269;
w14005 <= not w14003 and not w14004;
w14006 <= not w14002 and w14005;
w14007 <= w328 and w11277;
w14008 <= w14006 and not w14007;
w14009 <= a(59) and not w14008;
w14010 <= a(59) and not w14009;
w14011 <= not w14008 and not w14009;
w14012 <= not w14010 and not w14011;
w14013 <= w14001 and not w14012;
w14014 <= not w14001 and w14012;
w14015 <= not w13979 and not w14014;
w14016 <= not w14013 and w14015;
w14017 <= not w13979 and not w14016;
w14018 <= not w14013 and not w14016;
w14019 <= not w14014 and w14018;
w14020 <= not w14017 and not w14019;
w14021 <= b(11) and w10169;
w14022 <= b(9) and w10539;
w14023 <= b(10) and w10164;
w14024 <= not w14022 and not w14023;
w14025 <= not w14021 and w14024;
w14026 <= w561 and w10172;
w14027 <= w14025 and not w14026;
w14028 <= a(56) and not w14027;
w14029 <= a(56) and not w14028;
w14030 <= not w14027 and not w14028;
w14031 <= not w14029 and not w14030;
w14032 <= w14020 and w14031;
w14033 <= not w14020 and not w14031;
w14034 <= not w14032 and not w14033;
w14035 <= not w13978 and w14034;
w14036 <= w13978 and not w14034;
w14037 <= not w14035 and not w14036;
w14038 <= not w13977 and w14037;
w14039 <= w14037 and not w14038;
w14040 <= not w13977 and not w14038;
w14041 <= not w14039 and not w14040;
w14042 <= not w13966 and w14041;
w14043 <= w13966 and not w14041;
w14044 <= not w14042 and not w14043;
w14045 <= b(17) and w8105;
w14046 <= b(15) and w8458;
w14047 <= b(16) and w8100;
w14048 <= not w14046 and not w14047;
w14049 <= not w14045 and w14048;
w14050 <= w1099 and w8108;
w14051 <= w14049 and not w14050;
w14052 <= a(50) and not w14051;
w14053 <= a(50) and not w14052;
w14054 <= not w14051 and not w14052;
w14055 <= not w14053 and not w14054;
w14056 <= not w14044 and not w14055;
w14057 <= w14044 and w14055;
w14058 <= not w14056 and not w14057;
w14059 <= w13965 and not w14058;
w14060 <= not w13965 and w14058;
w14061 <= not w14059 and not w14060;
w14062 <= b(20) and w7189;
w14063 <= b(18) and w7530;
w14064 <= b(19) and w7184;
w14065 <= not w14063 and not w14064;
w14066 <= not w14062 and w14065;
w14067 <= w1589 and w7192;
w14068 <= w14066 and not w14067;
w14069 <= a(47) and not w14068;
w14070 <= a(47) and not w14069;
w14071 <= not w14068 and not w14069;
w14072 <= not w14070 and not w14071;
w14073 <= w14061 and not w14072;
w14074 <= w14061 and not w14073;
w14075 <= not w14072 and not w14073;
w14076 <= not w14074 and not w14075;
w14077 <= not w13964 and w14076;
w14078 <= w13964 and not w14076;
w14079 <= not w14077 and not w14078;
w14080 <= b(23) and w6338;
w14081 <= b(21) and w6645;
w14082 <= b(22) and w6333;
w14083 <= not w14081 and not w14082;
w14084 <= not w14080 and w14083;
w14085 <= w2043 and w6341;
w14086 <= w14084 and not w14085;
w14087 <= a(44) and not w14086;
w14088 <= a(44) and not w14087;
w14089 <= not w14086 and not w14087;
w14090 <= not w14088 and not w14089;
w14091 <= not w14079 and not w14090;
w14092 <= w14079 and w14090;
w14093 <= not w14091 and not w14092;
w14094 <= w13963 and not w14093;
w14095 <= not w13963 and w14093;
w14096 <= not w14094 and not w14095;
w14097 <= b(26) and w5520;
w14098 <= b(24) and w5802;
w14099 <= b(25) and w5515;
w14100 <= not w14098 and not w14099;
w14101 <= not w14097 and w14100;
w14102 <= w2556 and w5523;
w14103 <= w14101 and not w14102;
w14104 <= a(41) and not w14103;
w14105 <= a(41) and not w14104;
w14106 <= not w14103 and not w14104;
w14107 <= not w14105 and not w14106;
w14108 <= w14096 and not w14107;
w14109 <= w14096 and not w14108;
w14110 <= not w14107 and not w14108;
w14111 <= not w14109 and not w14110;
w14112 <= not w13758 and not w13764;
w14113 <= w14111 and w14112;
w14114 <= not w14111 and not w14112;
w14115 <= not w14113 and not w14114;
w14116 <= b(29) and w4778;
w14117 <= b(27) and w5020;
w14118 <= b(28) and w4773;
w14119 <= not w14117 and not w14118;
w14120 <= not w14116 and w14119;
w14121 <= w3126 and w4781;
w14122 <= w14120 and not w14121;
w14123 <= a(38) and not w14122;
w14124 <= a(38) and not w14123;
w14125 <= not w14122 and not w14123;
w14126 <= not w14124 and not w14125;
w14127 <= w14115 and not w14126;
w14128 <= w14115 and not w14127;
w14129 <= not w14126 and not w14127;
w14130 <= not w14128 and not w14129;
w14131 <= not w13777 and not w13783;
w14132 <= w14130 and w14131;
w14133 <= not w14130 and not w14131;
w14134 <= not w14132 and not w14133;
w14135 <= b(32) and w4030;
w14136 <= b(30) and w4275;
w14137 <= b(31) and w4025;
w14138 <= not w14136 and not w14137;
w14139 <= not w14135 and w14138;
w14140 <= w3756 and w4033;
w14141 <= w14139 and not w14140;
w14142 <= a(35) and not w14141;
w14143 <= a(35) and not w14142;
w14144 <= not w14141 and not w14142;
w14145 <= not w14143 and not w14144;
w14146 <= w14134 and not w14145;
w14147 <= not w14134 and w14145;
w14148 <= not w13962 and not w14147;
w14149 <= not w14146 and w14148;
w14150 <= not w13962 and not w14149;
w14151 <= not w14146 and not w14149;
w14152 <= not w14147 and w14151;
w14153 <= not w14150 and not w14152;
w14154 <= b(35) and w3381;
w14155 <= b(33) and w3586;
w14156 <= b(34) and w3376;
w14157 <= not w14155 and not w14156;
w14158 <= not w14154 and w14157;
w14159 <= w3384 and w4439;
w14160 <= w14158 and not w14159;
w14161 <= a(32) and not w14160;
w14162 <= a(32) and not w14161;
w14163 <= not w14160 and not w14161;
w14164 <= not w14162 and not w14163;
w14165 <= not w14153 and not w14164;
w14166 <= not w14153 and not w14165;
w14167 <= not w14164 and not w14165;
w14168 <= not w14166 and not w14167;
w14169 <= not w13803 and not w13810;
w14170 <= w14168 and w14169;
w14171 <= not w14168 and not w14169;
w14172 <= not w14170 and not w14171;
w14173 <= b(38) and w2793;
w14174 <= b(36) and w2986;
w14175 <= b(37) and w2788;
w14176 <= not w14174 and not w14175;
w14177 <= not w14173 and w14176;
w14178 <= w2796 and w4948;
w14179 <= w14177 and not w14178;
w14180 <= a(29) and not w14179;
w14181 <= a(29) and not w14180;
w14182 <= not w14179 and not w14180;
w14183 <= not w14181 and not w14182;
w14184 <= w14172 and not w14183;
w14185 <= w14172 and not w14184;
w14186 <= not w14183 and not w14184;
w14187 <= not w14185 and not w14186;
w14188 <= not w13823 and not w13829;
w14189 <= w14187 and w14188;
w14190 <= not w14187 and not w14188;
w14191 <= not w14189 and not w14190;
w14192 <= b(41) and w2282;
w14193 <= b(39) and w2428;
w14194 <= b(40) and w2277;
w14195 <= not w14193 and not w14194;
w14196 <= not w14192 and w14195;
w14197 <= w2285 and w5962;
w14198 <= w14196 and not w14197;
w14199 <= a(26) and not w14198;
w14200 <= a(26) and not w14199;
w14201 <= not w14198 and not w14199;
w14202 <= not w14200 and not w14201;
w14203 <= w14191 and not w14202;
w14204 <= not w14191 and w14202;
w14205 <= not w13961 and not w14204;
w14206 <= not w14203 and w14205;
w14207 <= not w13961 and not w14206;
w14208 <= not w14203 and not w14206;
w14209 <= not w14204 and w14208;
w14210 <= not w14207 and not w14209;
w14211 <= b(44) and w1791;
w14212 <= b(42) and w1941;
w14213 <= b(43) and w1786;
w14214 <= not w14212 and not w14213;
w14215 <= not w14211 and w14214;
w14216 <= w1794 and w6815;
w14217 <= w14215 and not w14216;
w14218 <= a(23) and not w14217;
w14219 <= a(23) and not w14218;
w14220 <= not w14217 and not w14218;
w14221 <= not w14219 and not w14220;
w14222 <= not w14210 and not w14221;
w14223 <= not w14210 and not w14222;
w14224 <= not w14221 and not w14222;
w14225 <= not w14223 and not w14224;
w14226 <= not w13850 and not w13861;
w14227 <= not w13865 and not w14226;
w14228 <= not w14225 and not w14227;
w14229 <= w14225 and w14227;
w14230 <= not w14228 and not w14229;
w14231 <= not w13960 and w14230;
w14232 <= not w13960 and not w14231;
w14233 <= w14230 and not w14231;
w14234 <= not w14232 and not w14233;
w14235 <= not w13949 and not w14234;
w14236 <= not w13949 and not w14235;
w14237 <= not w14234 and not w14235;
w14238 <= not w14236 and not w14237;
w14239 <= b(50) and w1045;
w14240 <= b(48) and w1134;
w14241 <= b(49) and w1040;
w14242 <= not w14240 and not w14241;
w14243 <= not w14239 and w14242;
w14244 <= w1048 and w8692;
w14245 <= w14243 and not w14244;
w14246 <= a(17) and not w14245;
w14247 <= a(17) and not w14246;
w14248 <= not w14245 and not w14246;
w14249 <= not w14247 and not w14248;
w14250 <= w14238 and w14249;
w14251 <= not w14238 and not w14249;
w14252 <= not w14250 and not w14251;
w14253 <= not w13948 and w14252;
w14254 <= w13948 and not w14252;
w14255 <= not w14253 and not w14254;
w14256 <= not w13947 and w14255;
w14257 <= w14255 and not w14256;
w14258 <= not w13947 and not w14256;
w14259 <= not w14257 and not w14258;
w14260 <= not w13884 and not w13887;
w14261 <= w14259 and w14260;
w14262 <= not w14259 and not w14260;
w14263 <= not w14261 and not w14262;
w14264 <= b(56) and w443;
w14265 <= b(54) and w510;
w14266 <= b(55) and w438;
w14267 <= not w14265 and not w14266;
w14268 <= not w14264 and w14267;
w14269 <= w446 and w10451;
w14270 <= w14268 and not w14269;
w14271 <= a(11) and not w14270;
w14272 <= a(11) and not w14271;
w14273 <= not w14270 and not w14271;
w14274 <= not w14272 and not w14273;
w14275 <= not w14263 and w14274;
w14276 <= w14263 and not w14274;
w14277 <= not w14275 and not w14276;
w14278 <= b(59) and w254;
w14279 <= b(57) and w284;
w14280 <= b(58) and w249;
w14281 <= not w14279 and not w14280;
w14282 <= not w14278 and w14281;
w14283 <= w257 and w11922;
w14284 <= w14282 and not w14283;
w14285 <= a(8) and not w14284;
w14286 <= a(8) and not w14285;
w14287 <= not w14284 and not w14285;
w14288 <= not w14286 and not w14287;
w14289 <= w14277 and not w14288;
w14290 <= w14277 and not w14289;
w14291 <= not w14288 and not w14289;
w14292 <= not w14290 and not w14291;
w14293 <= not w13890 and not w13893;
w14294 <= w14292 and w14293;
w14295 <= not w14292 and not w14293;
w14296 <= not w14294 and not w14295;
w14297 <= b(62) and w105;
w14298 <= b(60) and w146;
w14299 <= b(61) and w100;
w14300 <= not w14298 and not w14299;
w14301 <= not w14297 and w14300;
w14302 <= w108 and w13113;
w14303 <= w14301 and not w14302;
w14304 <= a(5) and not w14303;
w14305 <= a(5) and not w14304;
w14306 <= not w14303 and not w14304;
w14307 <= not w14305 and not w14306;
w14308 <= w14296 and not w14307;
w14309 <= w14296 and not w14308;
w14310 <= not w14307 and not w14308;
w14311 <= not w14309 and not w14310;
w14312 <= not w13910 and not w13921;
w14313 <= not w13907 and not w14312;
w14314 <= w12 and w13540;
w14315 <= not a(2) and not w14314;
w14316 <= b(63) and w27;
w14317 <= not w14314 and not w14316;
w14318 <= a(2) and not w14317;
w14319 <= not w14315 and not w14318;
w14320 <= not w14313 and w14319;
w14321 <= w14313 and not w14319;
w14322 <= not w14320 and not w14321;
w14323 <= not w14311 and w14322;
w14324 <= not w14311 and not w14323;
w14325 <= w14322 and not w14323;
w14326 <= not w14324 and not w14325;
w14327 <= not w13925 and not w13928;
w14328 <= w14326 and w14327;
w14329 <= not w14326 and not w14327;
w14330 <= not w14328 and not w14329;
w14331 <= not w13931 and not w13934;
w14332 <= w14330 and not w14331;
w14333 <= not w14330 and w14331;
w14334 <= not w14332 and not w14333;
w14335 <= not w14295 and not w14308;
w14336 <= b(63) and w105;
w14337 <= b(61) and w146;
w14338 <= b(62) and w100;
w14339 <= not w14337 and not w14338;
w14340 <= not w14336 and w14339;
w14341 <= w108 and w13514;
w14342 <= w14340 and not w14341;
w14343 <= a(5) and not w14342;
w14344 <= a(5) and not w14343;
w14345 <= not w14342 and not w14343;
w14346 <= not w14344 and not w14345;
w14347 <= not w14335 and not w14346;
w14348 <= not w14335 and not w14347;
w14349 <= not w14346 and not w14347;
w14350 <= not w14348 and not w14349;
w14351 <= b(57) and w443;
w14352 <= b(55) and w510;
w14353 <= b(56) and w438;
w14354 <= not w14352 and not w14353;
w14355 <= not w14351 and w14354;
w14356 <= w446 and w11153;
w14357 <= w14355 and not w14356;
w14358 <= a(11) and not w14357;
w14359 <= a(11) and not w14358;
w14360 <= not w14357 and not w14358;
w14361 <= not w14359 and not w14360;
w14362 <= not w14256 and not w14262;
w14363 <= w14361 and w14362;
w14364 <= not w14361 and not w14362;
w14365 <= not w14363 and not w14364;
w14366 <= b(51) and w1045;
w14367 <= b(49) and w1134;
w14368 <= b(50) and w1040;
w14369 <= not w14367 and not w14368;
w14370 <= not w14366 and w14369;
w14371 <= w1048 and w8719;
w14372 <= w14370 and not w14371;
w14373 <= a(17) and not w14372;
w14374 <= a(17) and not w14373;
w14375 <= not w14372 and not w14373;
w14376 <= not w14374 and not w14375;
w14377 <= not w14231 and not w14235;
w14378 <= w14376 and w14377;
w14379 <= not w14376 and not w14377;
w14380 <= not w14378 and not w14379;
w14381 <= b(48) and w1370;
w14382 <= b(46) and w1506;
w14383 <= b(47) and w1365;
w14384 <= not w14382 and not w14383;
w14385 <= not w14381 and w14384;
w14386 <= w1373 and w7752;
w14387 <= w14385 and not w14386;
w14388 <= a(20) and not w14387;
w14389 <= a(20) and not w14388;
w14390 <= not w14387 and not w14388;
w14391 <= not w14389 and not w14390;
w14392 <= not w14222 and not w14228;
w14393 <= w14391 and w14392;
w14394 <= not w14391 and not w14392;
w14395 <= not w14393 and not w14394;
w14396 <= b(45) and w1791;
w14397 <= b(43) and w1941;
w14398 <= b(44) and w1786;
w14399 <= not w14397 and not w14398;
w14400 <= not w14396 and w14399;
w14401 <= w1794 and w7104;
w14402 <= w14400 and not w14401;
w14403 <= a(23) and not w14402;
w14404 <= a(23) and not w14403;
w14405 <= not w14402 and not w14403;
w14406 <= not w14404 and not w14405;
w14407 <= not w14208 and w14406;
w14408 <= w14208 and not w14406;
w14409 <= not w14407 and not w14408;
w14410 <= b(42) and w2282;
w14411 <= b(40) and w2428;
w14412 <= b(41) and w2277;
w14413 <= not w14411 and not w14412;
w14414 <= not w14410 and w14413;
w14415 <= w2285 and w6232;
w14416 <= w14414 and not w14415;
w14417 <= a(26) and not w14416;
w14418 <= a(26) and not w14417;
w14419 <= not w14416 and not w14417;
w14420 <= not w14418 and not w14419;
w14421 <= not w14184 and not w14190;
w14422 <= w14420 and w14421;
w14423 <= not w14420 and not w14421;
w14424 <= not w14422 and not w14423;
w14425 <= not w14165 and not w14171;
w14426 <= b(39) and w2793;
w14427 <= b(37) and w2986;
w14428 <= b(38) and w2788;
w14429 <= not w14427 and not w14428;
w14430 <= not w14426 and w14429;
w14431 <= not w2796 and w14430;
w14432 <= not w5194 and w14430;
w14433 <= not w14431 and not w14432;
w14434 <= a(29) and not w14433;
w14435 <= not a(29) and w14433;
w14436 <= not w14434 and not w14435;
w14437 <= not w14425 and not w14436;
w14438 <= w14425 and w14436;
w14439 <= not w14437 and not w14438;
w14440 <= b(33) and w4030;
w14441 <= b(31) and w4275;
w14442 <= b(32) and w4025;
w14443 <= not w14441 and not w14442;
w14444 <= not w14440 and w14443;
w14445 <= w3966 and w4033;
w14446 <= w14444 and not w14445;
w14447 <= a(35) and not w14446;
w14448 <= a(35) and not w14447;
w14449 <= not w14446 and not w14447;
w14450 <= not w14448 and not w14449;
w14451 <= b(24) and w6338;
w14452 <= b(22) and w6645;
w14453 <= b(23) and w6333;
w14454 <= not w14452 and not w14453;
w14455 <= not w14451 and w14454;
w14456 <= w2201 and w6341;
w14457 <= w14455 and not w14456;
w14458 <= a(44) and not w14457;
w14459 <= a(44) and not w14458;
w14460 <= not w14457 and not w14458;
w14461 <= not w14459 and not w14460;
w14462 <= b(15) and w9082;
w14463 <= b(13) and w9475;
w14464 <= b(14) and w9077;
w14465 <= not w14463 and not w14464;
w14466 <= not w14462 and w14465;
w14467 <= w874 and w9085;
w14468 <= w14466 and not w14467;
w14469 <= a(53) and not w14468;
w14470 <= a(53) and not w14469;
w14471 <= not w14468 and not w14469;
w14472 <= not w14470 and not w14471;
w14473 <= not w14033 and not w14035;
w14474 <= not w13994 and not w14000;
w14475 <= b(2) and w13646;
w14476 <= b(3) and not w13231;
w14477 <= not w14475 and not w14476;
w14478 <= a(2) and not w14477;
w14479 <= not a(2) and w14477;
w14480 <= not w14478 and not w14479;
w14481 <= b(6) and w12411;
w14482 <= b(4) and w12790;
w14483 <= b(5) and w12406;
w14484 <= not w14482 and not w14483;
w14485 <= not w14481 and w14484;
w14486 <= not w12414 and w14485;
w14487 <= not w202 and w14485;
w14488 <= not w14486 and not w14487;
w14489 <= a(62) and not w14488;
w14490 <= not a(62) and w14488;
w14491 <= not w14489 and not w14490;
w14492 <= w14480 and not w14491;
w14493 <= not w14480 and w14491;
w14494 <= not w14492 and not w14493;
w14495 <= not w14474 and w14494;
w14496 <= w14474 and not w14494;
w14497 <= not w14495 and not w14496;
w14498 <= b(9) and w11274;
w14499 <= b(7) and w11639;
w14500 <= b(8) and w11269;
w14501 <= not w14499 and not w14500;
w14502 <= not w14498 and w14501;
w14503 <= w394 and w11277;
w14504 <= w14502 and not w14503;
w14505 <= a(59) and not w14504;
w14506 <= a(59) and not w14505;
w14507 <= not w14504 and not w14505;
w14508 <= not w14506 and not w14507;
w14509 <= w14497 and not w14508;
w14510 <= w14497 and not w14509;
w14511 <= not w14508 and not w14509;
w14512 <= not w14510 and not w14511;
w14513 <= not w14018 and w14512;
w14514 <= w14018 and not w14512;
w14515 <= not w14513 and not w14514;
w14516 <= b(12) and w10169;
w14517 <= b(10) and w10539;
w14518 <= b(11) and w10164;
w14519 <= not w14517 and not w14518;
w14520 <= not w14516 and w14519;
w14521 <= w585 and w10172;
w14522 <= w14520 and not w14521;
w14523 <= a(56) and not w14522;
w14524 <= a(56) and not w14523;
w14525 <= not w14522 and not w14523;
w14526 <= not w14524 and not w14525;
w14527 <= w14515 and w14526;
w14528 <= not w14515 and not w14526;
w14529 <= not w14527 and not w14528;
w14530 <= not w14473 and w14529;
w14531 <= w14473 and not w14529;
w14532 <= not w14530 and not w14531;
w14533 <= not w14472 and w14532;
w14534 <= w14532 and not w14533;
w14535 <= not w14472 and not w14533;
w14536 <= not w14534 and not w14535;
w14537 <= not w13966 and not w14041;
w14538 <= not w14038 and not w14537;
w14539 <= w14536 and w14538;
w14540 <= not w14536 and not w14538;
w14541 <= not w14539 and not w14540;
w14542 <= b(18) and w8105;
w14543 <= b(16) and w8458;
w14544 <= b(17) and w8100;
w14545 <= not w14543 and not w14544;
w14546 <= not w14542 and w14545;
w14547 <= w1309 and w8108;
w14548 <= w14546 and not w14547;
w14549 <= a(50) and not w14548;
w14550 <= a(50) and not w14549;
w14551 <= not w14548 and not w14549;
w14552 <= not w14550 and not w14551;
w14553 <= w14541 and not w14552;
w14554 <= w14541 and not w14553;
w14555 <= not w14552 and not w14553;
w14556 <= not w14554 and not w14555;
w14557 <= not w14056 and not w14060;
w14558 <= w14556 and w14557;
w14559 <= not w14556 and not w14557;
w14560 <= not w14558 and not w14559;
w14561 <= b(21) and w7189;
w14562 <= b(19) and w7530;
w14563 <= b(20) and w7184;
w14564 <= not w14562 and not w14563;
w14565 <= not w14561 and w14564;
w14566 <= w1727 and w7192;
w14567 <= w14565 and not w14566;
w14568 <= a(47) and not w14567;
w14569 <= a(47) and not w14568;
w14570 <= not w14567 and not w14568;
w14571 <= not w14569 and not w14570;
w14572 <= not w14560 and w14571;
w14573 <= w14560 and not w14571;
w14574 <= not w14572 and not w14573;
w14575 <= not w13964 and not w14076;
w14576 <= not w14073 and not w14575;
w14577 <= w14574 and not w14576;
w14578 <= not w14574 and w14576;
w14579 <= not w14577 and not w14578;
w14580 <= not w14461 and w14579;
w14581 <= w14579 and not w14580;
w14582 <= not w14461 and not w14580;
w14583 <= not w14581 and not w14582;
w14584 <= not w14091 and not w14095;
w14585 <= w14583 and w14584;
w14586 <= not w14583 and not w14584;
w14587 <= not w14585 and not w14586;
w14588 <= b(27) and w5520;
w14589 <= b(25) and w5802;
w14590 <= b(26) and w5515;
w14591 <= not w14589 and not w14590;
w14592 <= not w14588 and w14591;
w14593 <= w2733 and w5523;
w14594 <= w14592 and not w14593;
w14595 <= a(41) and not w14594;
w14596 <= a(41) and not w14595;
w14597 <= not w14594 and not w14595;
w14598 <= not w14596 and not w14597;
w14599 <= w14587 and not w14598;
w14600 <= w14587 and not w14599;
w14601 <= not w14598 and not w14599;
w14602 <= not w14600 and not w14601;
w14603 <= not w14108 and not w14114;
w14604 <= w14602 and w14603;
w14605 <= not w14602 and not w14603;
w14606 <= not w14604 and not w14605;
w14607 <= b(30) and w4778;
w14608 <= b(28) and w5020;
w14609 <= b(29) and w4773;
w14610 <= not w14608 and not w14609;
w14611 <= not w14607 and w14610;
w14612 <= w3320 and w4781;
w14613 <= w14611 and not w14612;
w14614 <= a(38) and not w14613;
w14615 <= a(38) and not w14614;
w14616 <= not w14613 and not w14614;
w14617 <= not w14615 and not w14616;
w14618 <= not w14606 and w14617;
w14619 <= w14606 and not w14617;
w14620 <= not w14618 and not w14619;
w14621 <= not w14127 and not w14133;
w14622 <= w14620 and not w14621;
w14623 <= not w14620 and w14621;
w14624 <= not w14622 and not w14623;
w14625 <= not w14450 and w14624;
w14626 <= w14624 and not w14625;
w14627 <= not w14450 and not w14625;
w14628 <= not w14626 and not w14627;
w14629 <= b(36) and w3381;
w14630 <= b(34) and w3586;
w14631 <= b(35) and w3376;
w14632 <= not w14630 and not w14631;
w14633 <= not w14629 and w14632;
w14634 <= not w3384 and w14633;
w14635 <= not w4665 and w14633;
w14636 <= not w14634 and not w14635;
w14637 <= a(32) and not w14636;
w14638 <= not a(32) and w14636;
w14639 <= not w14637 and not w14638;
w14640 <= not w14151 and not w14639;
w14641 <= not w14151 and not w14640;
w14642 <= not w14639 and not w14640;
w14643 <= not w14641 and not w14642;
w14644 <= not w14628 and not w14643;
w14645 <= not w14628 and not w14644;
w14646 <= not w14643 and not w14644;
w14647 <= not w14645 and not w14646;
w14648 <= w14439 and not w14647;
w14649 <= w14439 and not w14648;
w14650 <= not w14647 and not w14648;
w14651 <= not w14649 and not w14650;
w14652 <= w14424 and not w14651;
w14653 <= not w14424 and w14651;
w14654 <= not w14409 and not w14653;
w14655 <= not w14652 and w14654;
w14656 <= not w14409 and not w14655;
w14657 <= not w14653 and not w14655;
w14658 <= not w14652 and w14657;
w14659 <= not w14656 and not w14658;
w14660 <= w14395 and not w14659;
w14661 <= not w14395 and w14659;
w14662 <= w14380 and not w14661;
w14663 <= not w14660 and w14662;
w14664 <= w14380 and not w14663;
w14665 <= not w14661 and not w14663;
w14666 <= not w14660 and w14665;
w14667 <= not w14664 and not w14666;
w14668 <= not w14251 and not w14253;
w14669 <= b(54) and w694;
w14670 <= b(52) and w799;
w14671 <= b(53) and w689;
w14672 <= not w14670 and not w14671;
w14673 <= not w14669 and w14672;
w14674 <= not w697 and w14673;
w14675 <= not w9741 and w14673;
w14676 <= not w14674 and not w14675;
w14677 <= a(14) and not w14676;
w14678 <= not a(14) and w14676;
w14679 <= not w14677 and not w14678;
w14680 <= not w14668 and not w14679;
w14681 <= not w14668 and not w14680;
w14682 <= not w14679 and not w14680;
w14683 <= not w14681 and not w14682;
w14684 <= not w14667 and not w14683;
w14685 <= not w14667 and not w14684;
w14686 <= not w14683 and not w14684;
w14687 <= not w14685 and not w14686;
w14688 <= w14365 and not w14687;
w14689 <= w14365 and not w14688;
w14690 <= not w14687 and not w14688;
w14691 <= not w14689 and not w14690;
w14692 <= b(60) and w254;
w14693 <= b(58) and w284;
w14694 <= b(59) and w249;
w14695 <= not w14693 and not w14694;
w14696 <= not w14692 and w14695;
w14697 <= w257 and w11954;
w14698 <= w14696 and not w14697;
w14699 <= a(8) and not w14698;
w14700 <= a(8) and not w14699;
w14701 <= not w14698 and not w14699;
w14702 <= not w14700 and not w14701;
w14703 <= not w14276 and not w14289;
w14704 <= not w14702 and not w14703;
w14705 <= not w14702 and not w14704;
w14706 <= not w14703 and not w14704;
w14707 <= not w14705 and not w14706;
w14708 <= not w14691 and not w14707;
w14709 <= not w14691 and not w14708;
w14710 <= not w14707 and not w14708;
w14711 <= not w14709 and not w14710;
w14712 <= not w14350 and not w14711;
w14713 <= not w14350 and not w14712;
w14714 <= not w14711 and not w14712;
w14715 <= not w14713 and not w14714;
w14716 <= not w14320 and not w14323;
w14717 <= w14715 and w14716;
w14718 <= not w14715 and not w14716;
w14719 <= not w14717 and not w14718;
w14720 <= not w14329 and not w14332;
w14721 <= w14719 and not w14720;
w14722 <= not w14719 and w14720;
w14723 <= not w14721 and not w14722;
w14724 <= not w14718 and not w14721;
w14725 <= not w14347 and not w14712;
w14726 <= b(55) and w694;
w14727 <= b(53) and w799;
w14728 <= b(54) and w689;
w14729 <= not w14727 and not w14728;
w14730 <= not w14726 and w14729;
w14731 <= w697 and w10427;
w14732 <= w14730 and not w14731;
w14733 <= a(14) and not w14732;
w14734 <= a(14) and not w14733;
w14735 <= not w14732 and not w14733;
w14736 <= not w14734 and not w14735;
w14737 <= not w14379 and not w14663;
w14738 <= w14736 and w14737;
w14739 <= not w14736 and not w14737;
w14740 <= not w14738 and not w14739;
w14741 <= b(49) and w1370;
w14742 <= b(47) and w1506;
w14743 <= b(48) and w1365;
w14744 <= not w14742 and not w14743;
w14745 <= not w14741 and w14744;
w14746 <= w1373 and w8368;
w14747 <= w14745 and not w14746;
w14748 <= a(20) and not w14747;
w14749 <= a(20) and not w14748;
w14750 <= not w14747 and not w14748;
w14751 <= not w14749 and not w14750;
w14752 <= not w14208 and not w14406;
w14753 <= not w14655 and not w14752;
w14754 <= w14751 and w14753;
w14755 <= not w14751 and not w14753;
w14756 <= not w14754 and not w14755;
w14757 <= b(43) and w2282;
w14758 <= b(41) and w2428;
w14759 <= b(42) and w2277;
w14760 <= not w14758 and not w14759;
w14761 <= not w14757 and w14760;
w14762 <= w2285 and w6258;
w14763 <= w14761 and not w14762;
w14764 <= a(26) and not w14763;
w14765 <= a(26) and not w14764;
w14766 <= not w14763 and not w14764;
w14767 <= not w14765 and not w14766;
w14768 <= not w14437 and not w14648;
w14769 <= w14767 and w14768;
w14770 <= not w14767 and not w14768;
w14771 <= not w14769 and not w14770;
w14772 <= not w14622 and not w14625;
w14773 <= b(37) and w3381;
w14774 <= b(35) and w3586;
w14775 <= b(36) and w3376;
w14776 <= not w14774 and not w14775;
w14777 <= not w14773 and w14776;
w14778 <= not w3384 and w14777;
w14779 <= not w4924 and w14777;
w14780 <= not w14778 and not w14779;
w14781 <= a(32) and not w14780;
w14782 <= not a(32) and w14780;
w14783 <= not w14781 and not w14782;
w14784 <= not w14772 and not w14783;
w14785 <= w14772 and w14783;
w14786 <= not w14784 and not w14785;
w14787 <= b(34) and w4030;
w14788 <= b(32) and w4275;
w14789 <= b(33) and w4025;
w14790 <= not w14788 and not w14789;
w14791 <= not w14787 and w14790;
w14792 <= w4033 and w4209;
w14793 <= w14791 and not w14792;
w14794 <= a(35) and not w14793;
w14795 <= a(35) and not w14794;
w14796 <= not w14793 and not w14794;
w14797 <= not w14795 and not w14796;
w14798 <= not w14605 and not w14619;
w14799 <= b(16) and w9082;
w14800 <= b(14) and w9475;
w14801 <= b(15) and w9077;
w14802 <= not w14800 and not w14801;
w14803 <= not w14799 and w14802;
w14804 <= w980 and w9085;
w14805 <= w14803 and not w14804;
w14806 <= a(53) and not w14805;
w14807 <= a(53) and not w14806;
w14808 <= not w14805 and not w14806;
w14809 <= not w14807 and not w14808;
w14810 <= b(7) and w12411;
w14811 <= b(5) and w12790;
w14812 <= b(6) and w12406;
w14813 <= not w14811 and not w14812;
w14814 <= not w14810 and w14813;
w14815 <= w227 and w12414;
w14816 <= w14814 and not w14815;
w14817 <= a(62) and not w14816;
w14818 <= a(62) and not w14817;
w14819 <= not w14816 and not w14817;
w14820 <= not w14818 and not w14819;
w14821 <= b(3) and w13646;
w14822 <= b(4) and not w13231;
w14823 <= not w14821 and not w14822;
w14824 <= a(2) and not w14823;
w14825 <= a(2) and not w14824;
w14826 <= not w14823 and not w14824;
w14827 <= not w14825 and not w14826;
w14828 <= not w14820 and not w14827;
w14829 <= not w14820 and not w14828;
w14830 <= not w14827 and not w14828;
w14831 <= not w14829 and not w14830;
w14832 <= not w14478 and not w14492;
w14833 <= w14831 and w14832;
w14834 <= not w14831 and not w14832;
w14835 <= not w14833 and not w14834;
w14836 <= b(10) and w11274;
w14837 <= b(8) and w11639;
w14838 <= b(9) and w11269;
w14839 <= not w14837 and not w14838;
w14840 <= not w14836 and w14839;
w14841 <= w481 and w11277;
w14842 <= w14840 and not w14841;
w14843 <= a(59) and not w14842;
w14844 <= a(59) and not w14843;
w14845 <= not w14842 and not w14843;
w14846 <= not w14844 and not w14845;
w14847 <= w14835 and not w14846;
w14848 <= w14835 and not w14847;
w14849 <= not w14846 and not w14847;
w14850 <= not w14848 and not w14849;
w14851 <= not w14495 and not w14509;
w14852 <= w14850 and w14851;
w14853 <= not w14850 and not w14851;
w14854 <= not w14852 and not w14853;
w14855 <= b(13) and w10169;
w14856 <= b(11) and w10539;
w14857 <= b(12) and w10164;
w14858 <= not w14856 and not w14857;
w14859 <= not w14855 and w14858;
w14860 <= w751 and w10172;
w14861 <= w14859 and not w14860;
w14862 <= a(56) and not w14861;
w14863 <= a(56) and not w14862;
w14864 <= not w14861 and not w14862;
w14865 <= not w14863 and not w14864;
w14866 <= not w14854 and w14865;
w14867 <= w14854 and not w14865;
w14868 <= not w14866 and not w14867;
w14869 <= not w14018 and not w14512;
w14870 <= not w14528 and not w14869;
w14871 <= w14868 and not w14870;
w14872 <= not w14868 and w14870;
w14873 <= not w14871 and not w14872;
w14874 <= not w14809 and w14873;
w14875 <= w14873 and not w14874;
w14876 <= not w14809 and not w14874;
w14877 <= not w14875 and not w14876;
w14878 <= not w14530 and not w14533;
w14879 <= w14877 and w14878;
w14880 <= not w14877 and not w14878;
w14881 <= not w14879 and not w14880;
w14882 <= b(19) and w8105;
w14883 <= b(17) and w8458;
w14884 <= b(18) and w8100;
w14885 <= not w14883 and not w14884;
w14886 <= not w14882 and w14885;
w14887 <= w1451 and w8108;
w14888 <= w14886 and not w14887;
w14889 <= a(50) and not w14888;
w14890 <= a(50) and not w14889;
w14891 <= not w14888 and not w14889;
w14892 <= not w14890 and not w14891;
w14893 <= w14881 and not w14892;
w14894 <= w14881 and not w14893;
w14895 <= not w14892 and not w14893;
w14896 <= not w14894 and not w14895;
w14897 <= not w14540 and not w14553;
w14898 <= w14896 and w14897;
w14899 <= not w14896 and not w14897;
w14900 <= not w14898 and not w14899;
w14901 <= b(22) and w7189;
w14902 <= b(20) and w7530;
w14903 <= b(21) and w7184;
w14904 <= not w14902 and not w14903;
w14905 <= not w14901 and w14904;
w14906 <= w1888 and w7192;
w14907 <= w14905 and not w14906;
w14908 <= a(47) and not w14907;
w14909 <= a(47) and not w14908;
w14910 <= not w14907 and not w14908;
w14911 <= not w14909 and not w14910;
w14912 <= w14900 and not w14911;
w14913 <= w14900 and not w14912;
w14914 <= not w14911 and not w14912;
w14915 <= not w14913 and not w14914;
w14916 <= not w14559 and not w14573;
w14917 <= not w14915 and not w14916;
w14918 <= not w14915 and not w14917;
w14919 <= not w14916 and not w14917;
w14920 <= not w14918 and not w14919;
w14921 <= b(25) and w6338;
w14922 <= b(23) and w6645;
w14923 <= b(24) and w6333;
w14924 <= not w14922 and not w14923;
w14925 <= not w14921 and w14924;
w14926 <= w2228 and w6341;
w14927 <= w14925 and not w14926;
w14928 <= a(44) and not w14927;
w14929 <= a(44) and not w14928;
w14930 <= not w14927 and not w14928;
w14931 <= not w14929 and not w14930;
w14932 <= not w14920 and not w14931;
w14933 <= not w14920 and not w14932;
w14934 <= not w14931 and not w14932;
w14935 <= not w14933 and not w14934;
w14936 <= not w14577 and not w14580;
w14937 <= w14935 and w14936;
w14938 <= not w14935 and not w14936;
w14939 <= not w14937 and not w14938;
w14940 <= b(28) and w5520;
w14941 <= b(26) and w5802;
w14942 <= b(27) and w5515;
w14943 <= not w14941 and not w14942;
w14944 <= not w14940 and w14943;
w14945 <= w2932 and w5523;
w14946 <= w14944 and not w14945;
w14947 <= a(41) and not w14946;
w14948 <= a(41) and not w14947;
w14949 <= not w14946 and not w14947;
w14950 <= not w14948 and not w14949;
w14951 <= w14939 and not w14950;
w14952 <= w14939 and not w14951;
w14953 <= not w14950 and not w14951;
w14954 <= not w14952 and not w14953;
w14955 <= not w14586 and not w14599;
w14956 <= w14954 and w14955;
w14957 <= not w14954 and not w14955;
w14958 <= not w14956 and not w14957;
w14959 <= b(31) and w4778;
w14960 <= b(29) and w5020;
w14961 <= b(30) and w4773;
w14962 <= not w14960 and not w14961;
w14963 <= not w14959 and w14962;
w14964 <= w3539 and w4781;
w14965 <= w14963 and not w14964;
w14966 <= a(38) and not w14965;
w14967 <= a(38) and not w14966;
w14968 <= not w14965 and not w14966;
w14969 <= not w14967 and not w14968;
w14970 <= not w14958 and w14969;
w14971 <= w14958 and not w14969;
w14972 <= not w14970 and not w14971;
w14973 <= not w14798 and w14972;
w14974 <= not w14798 and not w14973;
w14975 <= w14972 and not w14973;
w14976 <= not w14974 and not w14975;
w14977 <= not w14797 and not w14976;
w14978 <= not w14797 and not w14977;
w14979 <= not w14976 and not w14977;
w14980 <= not w14978 and not w14979;
w14981 <= not w14786 and w14980;
w14982 <= w14786 and not w14980;
w14983 <= not w14981 and not w14982;
w14984 <= not w14640 and not w14644;
w14985 <= b(40) and w2793;
w14986 <= b(38) and w2986;
w14987 <= b(39) and w2788;
w14988 <= not w14986 and not w14987;
w14989 <= not w14985 and w14988;
w14990 <= not w2796 and w14989;
w14991 <= not w5698 and w14989;
w14992 <= not w14990 and not w14991;
w14993 <= a(29) and not w14992;
w14994 <= not a(29) and w14992;
w14995 <= not w14993 and not w14994;
w14996 <= not w14984 and not w14995;
w14997 <= not w14984 and not w14996;
w14998 <= not w14995 and not w14996;
w14999 <= not w14997 and not w14998;
w15000 <= w14983 and not w14999;
w15001 <= w14983 and not w15000;
w15002 <= not w14999 and not w15000;
w15003 <= not w15001 and not w15002;
w15004 <= w14771 and not w15003;
w15005 <= w14771 and not w15004;
w15006 <= not w15003 and not w15004;
w15007 <= not w15005 and not w15006;
w15008 <= b(46) and w1791;
w15009 <= b(44) and w1941;
w15010 <= b(45) and w1786;
w15011 <= not w15009 and not w15010;
w15012 <= not w15008 and w15011;
w15013 <= w1794 and w7420;
w15014 <= w15012 and not w15013;
w15015 <= a(23) and not w15014;
w15016 <= a(23) and not w15015;
w15017 <= not w15014 and not w15015;
w15018 <= not w15016 and not w15017;
w15019 <= not w14423 and not w14652;
w15020 <= not w15018 and not w15019;
w15021 <= not w15018 and not w15020;
w15022 <= not w15019 and not w15020;
w15023 <= not w15021 and not w15022;
w15024 <= not w15007 and w15023;
w15025 <= w15007 and not w15023;
w15026 <= not w15024 and not w15025;
w15027 <= w14756 and not w15026;
w15028 <= w14756 and not w15027;
w15029 <= not w15026 and not w15027;
w15030 <= not w15028 and not w15029;
w15031 <= b(52) and w1045;
w15032 <= b(50) and w1134;
w15033 <= b(51) and w1040;
w15034 <= not w15032 and not w15033;
w15035 <= not w15031 and w15034;
w15036 <= w1048 and w9371;
w15037 <= w15035 and not w15036;
w15038 <= a(17) and not w15037;
w15039 <= a(17) and not w15038;
w15040 <= not w15037 and not w15038;
w15041 <= not w15039 and not w15040;
w15042 <= not w14394 and not w14660;
w15043 <= not w15041 and not w15042;
w15044 <= not w15041 and not w15043;
w15045 <= not w15042 and not w15043;
w15046 <= not w15044 and not w15045;
w15047 <= not w15030 and w15046;
w15048 <= w15030 and not w15046;
w15049 <= not w15047 and not w15048;
w15050 <= w14740 and not w15049;
w15051 <= w14740 and not w15050;
w15052 <= not w15049 and not w15050;
w15053 <= not w15051 and not w15052;
w15054 <= not w14680 and not w14684;
w15055 <= b(58) and w443;
w15056 <= b(56) and w510;
w15057 <= b(57) and w438;
w15058 <= not w15056 and not w15057;
w15059 <= not w15055 and w15058;
w15060 <= not w446 and w15059;
w15061 <= not w11179 and w15059;
w15062 <= not w15060 and not w15061;
w15063 <= a(11) and not w15062;
w15064 <= not a(11) and w15062;
w15065 <= not w15063 and not w15064;
w15066 <= not w15054 and not w15065;
w15067 <= not w15054 and not w15066;
w15068 <= not w15065 and not w15066;
w15069 <= not w15067 and not w15068;
w15070 <= not w15053 and not w15069;
w15071 <= not w15053 and not w15070;
w15072 <= not w15069 and not w15070;
w15073 <= not w15071 and not w15072;
w15074 <= not w14364 and not w14688;
w15075 <= b(61) and w254;
w15076 <= b(59) and w284;
w15077 <= b(60) and w249;
w15078 <= not w15076 and not w15077;
w15079 <= not w15075 and w15078;
w15080 <= not w257 and w15079;
w15081 <= not w12712 and w15079;
w15082 <= not w15080 and not w15081;
w15083 <= a(8) and not w15082;
w15084 <= not a(8) and w15082;
w15085 <= not w15083 and not w15084;
w15086 <= not w15074 and not w15085;
w15087 <= not w15074 and not w15086;
w15088 <= not w15085 and not w15086;
w15089 <= not w15087 and not w15088;
w15090 <= not w15073 and not w15089;
w15091 <= not w15073 and not w15090;
w15092 <= not w15089 and not w15090;
w15093 <= not w15091 and not w15092;
w15094 <= not w14704 and not w14708;
w15095 <= b(62) and w146;
w15096 <= b(63) and w100;
w15097 <= not w15095 and not w15096;
w15098 <= not w108 and w15097;
w15099 <= w13543 and w15097;
w15100 <= not w15098 and not w15099;
w15101 <= a(5) and not w15100;
w15102 <= not a(5) and w15100;
w15103 <= not w15101 and not w15102;
w15104 <= not w15094 and not w15103;
w15105 <= not w15094 and not w15104;
w15106 <= not w15103 and not w15104;
w15107 <= not w15105 and not w15106;
w15108 <= not w15093 and not w15107;
w15109 <= w15093 and not w15106;
w15110 <= not w15105 and w15109;
w15111 <= not w15108 and not w15110;
w15112 <= not w14725 and w15111;
w15113 <= not w14725 and not w15112;
w15114 <= w15111 and not w15112;
w15115 <= not w15113 and not w15114;
w15116 <= not w14724 and not w15115;
w15117 <= w14724 and not w15114;
w15118 <= not w15113 and w15117;
w15119 <= not w15116 and not w15118;
w15120 <= not w15112 and not w15116;
w15121 <= not w15104 and not w15108;
w15122 <= not w15086 and not w15090;
w15123 <= b(63) and w146;
w15124 <= w108 and w13540;
w15125 <= not w15123 and not w15124;
w15126 <= a(5) and not w15125;
w15127 <= a(5) and not w15126;
w15128 <= not w15125 and not w15126;
w15129 <= not w15127 and not w15128;
w15130 <= not w15122 and not w15129;
w15131 <= not w15122 and not w15130;
w15132 <= not w15129 and not w15130;
w15133 <= not w15131 and not w15132;
w15134 <= b(59) and w443;
w15135 <= b(57) and w510;
w15136 <= b(58) and w438;
w15137 <= not w15135 and not w15136;
w15138 <= not w15134 and w15137;
w15139 <= w446 and w11922;
w15140 <= w15138 and not w15139;
w15141 <= a(11) and not w15140;
w15142 <= a(11) and not w15141;
w15143 <= not w15140 and not w15141;
w15144 <= not w15142 and not w15143;
w15145 <= not w14739 and not w15050;
w15146 <= w15144 and w15145;
w15147 <= not w15144 and not w15145;
w15148 <= not w15146 and not w15147;
w15149 <= b(56) and w694;
w15150 <= b(54) and w799;
w15151 <= b(55) and w689;
w15152 <= not w15150 and not w15151;
w15153 <= not w15149 and w15152;
w15154 <= w697 and w10451;
w15155 <= w15153 and not w15154;
w15156 <= a(14) and not w15155;
w15157 <= a(14) and not w15156;
w15158 <= not w15155 and not w15156;
w15159 <= not w15157 and not w15158;
w15160 <= not w15030 and not w15046;
w15161 <= not w15043 and not w15160;
w15162 <= not w15159 and not w15161;
w15163 <= not w15159 and not w15162;
w15164 <= not w15161 and not w15162;
w15165 <= not w15163 and not w15164;
w15166 <= not w14755 and not w15027;
w15167 <= b(53) and w1045;
w15168 <= b(51) and w1134;
w15169 <= b(52) and w1040;
w15170 <= not w15168 and not w15169;
w15171 <= not w15167 and w15170;
w15172 <= not w1048 and w15171;
w15173 <= not w9715 and w15171;
w15174 <= not w15172 and not w15173;
w15175 <= a(17) and not w15174;
w15176 <= not a(17) and w15174;
w15177 <= not w15175 and not w15176;
w15178 <= not w15166 and not w15177;
w15179 <= w15166 and w15177;
w15180 <= not w15178 and not w15179;
w15181 <= b(50) and w1370;
w15182 <= b(48) and w1506;
w15183 <= b(49) and w1365;
w15184 <= not w15182 and not w15183;
w15185 <= not w15181 and w15184;
w15186 <= w1373 and w8692;
w15187 <= w15185 and not w15186;
w15188 <= a(20) and not w15187;
w15189 <= a(20) and not w15188;
w15190 <= not w15187 and not w15188;
w15191 <= not w15189 and not w15190;
w15192 <= not w15007 and not w15023;
w15193 <= not w15020 and not w15192;
w15194 <= not w15191 and not w15193;
w15195 <= not w15191 and not w15194;
w15196 <= not w15193 and not w15194;
w15197 <= not w15195 and not w15196;
w15198 <= b(47) and w1791;
w15199 <= b(45) and w1941;
w15200 <= b(46) and w1786;
w15201 <= not w15199 and not w15200;
w15202 <= not w15198 and w15201;
w15203 <= w1794 and w7446;
w15204 <= w15202 and not w15203;
w15205 <= a(23) and not w15204;
w15206 <= a(23) and not w15205;
w15207 <= not w15204 and not w15205;
w15208 <= not w15206 and not w15207;
w15209 <= not w14770 and not w15004;
w15210 <= w15208 and w15209;
w15211 <= not w15208 and not w15209;
w15212 <= not w15210 and not w15211;
w15213 <= b(41) and w2793;
w15214 <= b(39) and w2986;
w15215 <= b(40) and w2788;
w15216 <= not w15214 and not w15215;
w15217 <= not w15213 and w15216;
w15218 <= w2796 and w5962;
w15219 <= w15217 and not w15218;
w15220 <= a(29) and not w15219;
w15221 <= a(29) and not w15220;
w15222 <= not w15219 and not w15220;
w15223 <= not w15221 and not w15222;
w15224 <= not w14784 and not w14982;
w15225 <= w15223 and w15224;
w15226 <= not w15223 and not w15224;
w15227 <= not w15225 and not w15226;
w15228 <= b(35) and w4030;
w15229 <= b(33) and w4275;
w15230 <= b(34) and w4025;
w15231 <= not w15229 and not w15230;
w15232 <= not w15228 and w15231;
w15233 <= w4033 and w4439;
w15234 <= w15232 and not w15233;
w15235 <= a(35) and not w15234;
w15236 <= a(35) and not w15235;
w15237 <= not w15234 and not w15235;
w15238 <= not w15236 and not w15237;
w15239 <= b(23) and w7189;
w15240 <= b(21) and w7530;
w15241 <= b(22) and w7184;
w15242 <= not w15240 and not w15241;
w15243 <= not w15239 and w15242;
w15244 <= w2043 and w7192;
w15245 <= w15243 and not w15244;
w15246 <= a(47) and not w15245;
w15247 <= a(47) and not w15246;
w15248 <= not w15245 and not w15246;
w15249 <= not w15247 and not w15248;
w15250 <= b(14) and w10169;
w15251 <= b(12) and w10539;
w15252 <= b(13) and w10164;
w15253 <= not w15251 and not w15252;
w15254 <= not w15250 and w15253;
w15255 <= w777 and w10172;
w15256 <= w15254 and not w15255;
w15257 <= a(56) and not w15256;
w15258 <= a(56) and not w15257;
w15259 <= not w15256 and not w15257;
w15260 <= not w15258 and not w15259;
w15261 <= b(8) and w12411;
w15262 <= b(6) and w12790;
w15263 <= b(7) and w12406;
w15264 <= not w15262 and not w15263;
w15265 <= not w15261 and w15264;
w15266 <= w328 and w12414;
w15267 <= w15265 and not w15266;
w15268 <= a(62) and not w15267;
w15269 <= a(62) and not w15268;
w15270 <= not w15267 and not w15268;
w15271 <= not w15269 and not w15270;
w15272 <= b(4) and w13646;
w15273 <= b(5) and not w13231;
w15274 <= not w15272 and not w15273;
w15275 <= a(2) and not w15274;
w15276 <= a(2) and not w15275;
w15277 <= not w15274 and not w15275;
w15278 <= not w15276 and not w15277;
w15279 <= not w15271 and not w15278;
w15280 <= not w15271 and not w15279;
w15281 <= not w15278 and not w15279;
w15282 <= not w15280 and not w15281;
w15283 <= not w14824 and not w14828;
w15284 <= w15282 and w15283;
w15285 <= not w15282 and not w15283;
w15286 <= not w15284 and not w15285;
w15287 <= b(11) and w11274;
w15288 <= b(9) and w11639;
w15289 <= b(10) and w11269;
w15290 <= not w15288 and not w15289;
w15291 <= not w15287 and w15290;
w15292 <= w561 and w11277;
w15293 <= w15291 and not w15292;
w15294 <= a(59) and not w15293;
w15295 <= a(59) and not w15294;
w15296 <= not w15293 and not w15294;
w15297 <= not w15295 and not w15296;
w15298 <= not w15286 and w15297;
w15299 <= w15286 and not w15297;
w15300 <= not w15298 and not w15299;
w15301 <= not w14834 and not w14847;
w15302 <= w15300 and not w15301;
w15303 <= not w15300 and w15301;
w15304 <= not w15302 and not w15303;
w15305 <= not w15260 and w15304;
w15306 <= w15304 and not w15305;
w15307 <= not w15260 and not w15305;
w15308 <= not w15306 and not w15307;
w15309 <= not w14853 and not w14867;
w15310 <= not w15308 and not w15309;
w15311 <= not w15308 and not w15310;
w15312 <= not w15309 and not w15310;
w15313 <= not w15311 and not w15312;
w15314 <= b(17) and w9082;
w15315 <= b(15) and w9475;
w15316 <= b(16) and w9077;
w15317 <= not w15315 and not w15316;
w15318 <= not w15314 and w15317;
w15319 <= w1099 and w9085;
w15320 <= w15318 and not w15319;
w15321 <= a(53) and not w15320;
w15322 <= a(53) and not w15321;
w15323 <= not w15320 and not w15321;
w15324 <= not w15322 and not w15323;
w15325 <= not w15313 and not w15324;
w15326 <= not w15313 and not w15325;
w15327 <= not w15324 and not w15325;
w15328 <= not w15326 and not w15327;
w15329 <= not w14871 and not w14874;
w15330 <= w15328 and w15329;
w15331 <= not w15328 and not w15329;
w15332 <= not w15330 and not w15331;
w15333 <= b(20) and w8105;
w15334 <= b(18) and w8458;
w15335 <= b(19) and w8100;
w15336 <= not w15334 and not w15335;
w15337 <= not w15333 and w15336;
w15338 <= w1589 and w8108;
w15339 <= w15337 and not w15338;
w15340 <= a(50) and not w15339;
w15341 <= a(50) and not w15340;
w15342 <= not w15339 and not w15340;
w15343 <= not w15341 and not w15342;
w15344 <= not w15332 and w15343;
w15345 <= w15332 and not w15343;
w15346 <= not w15344 and not w15345;
w15347 <= not w14880 and not w14893;
w15348 <= w15346 and not w15347;
w15349 <= not w15346 and w15347;
w15350 <= not w15348 and not w15349;
w15351 <= not w15249 and w15350;
w15352 <= w15350 and not w15351;
w15353 <= not w15249 and not w15351;
w15354 <= not w15352 and not w15353;
w15355 <= not w14899 and not w14912;
w15356 <= w15354 and w15355;
w15357 <= not w15354 and not w15355;
w15358 <= not w15356 and not w15357;
w15359 <= b(26) and w6338;
w15360 <= b(24) and w6645;
w15361 <= b(25) and w6333;
w15362 <= not w15360 and not w15361;
w15363 <= not w15359 and w15362;
w15364 <= w2556 and w6341;
w15365 <= w15363 and not w15364;
w15366 <= a(44) and not w15365;
w15367 <= a(44) and not w15366;
w15368 <= not w15365 and not w15366;
w15369 <= not w15367 and not w15368;
w15370 <= w15358 and not w15369;
w15371 <= w15358 and not w15370;
w15372 <= not w15369 and not w15370;
w15373 <= not w15371 and not w15372;
w15374 <= not w14917 and not w14932;
w15375 <= w15373 and w15374;
w15376 <= not w15373 and not w15374;
w15377 <= not w15375 and not w15376;
w15378 <= b(29) and w5520;
w15379 <= b(27) and w5802;
w15380 <= b(28) and w5515;
w15381 <= not w15379 and not w15380;
w15382 <= not w15378 and w15381;
w15383 <= w3126 and w5523;
w15384 <= w15382 and not w15383;
w15385 <= a(41) and not w15384;
w15386 <= a(41) and not w15385;
w15387 <= not w15384 and not w15385;
w15388 <= not w15386 and not w15387;
w15389 <= w15377 and not w15388;
w15390 <= w15377 and not w15389;
w15391 <= not w15388 and not w15389;
w15392 <= not w15390 and not w15391;
w15393 <= not w14938 and not w14951;
w15394 <= w15392 and w15393;
w15395 <= not w15392 and not w15393;
w15396 <= not w15394 and not w15395;
w15397 <= b(32) and w4778;
w15398 <= b(30) and w5020;
w15399 <= b(31) and w4773;
w15400 <= not w15398 and not w15399;
w15401 <= not w15397 and w15400;
w15402 <= w3756 and w4781;
w15403 <= w15401 and not w15402;
w15404 <= a(38) and not w15403;
w15405 <= a(38) and not w15404;
w15406 <= not w15403 and not w15404;
w15407 <= not w15405 and not w15406;
w15408 <= not w15396 and w15407;
w15409 <= w15396 and not w15407;
w15410 <= not w15408 and not w15409;
w15411 <= not w14957 and not w14971;
w15412 <= w15410 and not w15411;
w15413 <= not w15410 and w15411;
w15414 <= not w15412 and not w15413;
w15415 <= not w15238 and w15414;
w15416 <= w15414 and not w15415;
w15417 <= not w15238 and not w15415;
w15418 <= not w15416 and not w15417;
w15419 <= not w14973 and not w14977;
w15420 <= b(38) and w3381;
w15421 <= b(36) and w3586;
w15422 <= b(37) and w3376;
w15423 <= not w15421 and not w15422;
w15424 <= not w15420 and w15423;
w15425 <= not w3384 and w15424;
w15426 <= not w4948 and w15424;
w15427 <= not w15425 and not w15426;
w15428 <= a(32) and not w15427;
w15429 <= not a(32) and w15427;
w15430 <= not w15428 and not w15429;
w15431 <= not w15419 and not w15430;
w15432 <= w15419 and w15430;
w15433 <= not w15431 and not w15432;
w15434 <= not w15418 and w15433;
w15435 <= not w15418 and not w15434;
w15436 <= w15433 and not w15434;
w15437 <= not w15435 and not w15436;
w15438 <= w15227 and not w15437;
w15439 <= w15227 and not w15438;
w15440 <= not w15437 and not w15438;
w15441 <= not w15439 and not w15440;
w15442 <= not w14996 and not w15000;
w15443 <= b(44) and w2282;
w15444 <= b(42) and w2428;
w15445 <= b(43) and w2277;
w15446 <= not w15444 and not w15445;
w15447 <= not w15443 and w15446;
w15448 <= not w2285 and w15447;
w15449 <= not w6815 and w15447;
w15450 <= not w15448 and not w15449;
w15451 <= a(26) and not w15450;
w15452 <= not a(26) and w15450;
w15453 <= not w15451 and not w15452;
w15454 <= not w15442 and not w15453;
w15455 <= not w15442 and not w15454;
w15456 <= not w15453 and not w15454;
w15457 <= not w15455 and not w15456;
w15458 <= not w15441 and not w15457;
w15459 <= not w15441 and not w15458;
w15460 <= not w15457 and not w15458;
w15461 <= not w15459 and not w15460;
w15462 <= w15212 and not w15461;
w15463 <= w15212 and not w15462;
w15464 <= not w15461 and not w15462;
w15465 <= not w15463 and not w15464;
w15466 <= not w15197 and w15465;
w15467 <= w15197 and not w15465;
w15468 <= not w15466 and not w15467;
w15469 <= w15180 and not w15468;
w15470 <= w15180 and not w15469;
w15471 <= not w15468 and not w15469;
w15472 <= not w15470 and not w15471;
w15473 <= not w15165 and w15472;
w15474 <= w15165 and not w15472;
w15475 <= not w15473 and not w15474;
w15476 <= w15148 and not w15475;
w15477 <= w15148 and not w15476;
w15478 <= not w15475 and not w15476;
w15479 <= not w15477 and not w15478;
w15480 <= not w15066 and not w15070;
w15481 <= b(62) and w254;
w15482 <= b(60) and w284;
w15483 <= b(61) and w249;
w15484 <= not w15482 and not w15483;
w15485 <= not w15481 and w15484;
w15486 <= not w257 and w15485;
w15487 <= not w13113 and w15485;
w15488 <= not w15486 and not w15487;
w15489 <= a(8) and not w15488;
w15490 <= not a(8) and w15488;
w15491 <= not w15489 and not w15490;
w15492 <= not w15480 and not w15491;
w15493 <= not w15480 and not w15492;
w15494 <= not w15491 and not w15492;
w15495 <= not w15493 and not w15494;
w15496 <= not w15479 and not w15495;
w15497 <= w15479 and not w15494;
w15498 <= not w15493 and w15497;
w15499 <= not w15496 and not w15498;
w15500 <= not w15133 and w15499;
w15501 <= w15133 and not w15499;
w15502 <= not w15500 and not w15501;
w15503 <= not w15121 and w15502;
w15504 <= not w15121 and not w15503;
w15505 <= w15502 and not w15503;
w15506 <= not w15504 and not w15505;
w15507 <= not w15120 and not w15506;
w15508 <= w15120 and not w15505;
w15509 <= not w15504 and w15508;
w15510 <= not w15507 and not w15509;
w15511 <= not w15503 and not w15507;
w15512 <= not w15130 and not w15500;
w15513 <= not w15492 and not w15496;
w15514 <= b(63) and w254;
w15515 <= b(61) and w284;
w15516 <= b(62) and w249;
w15517 <= not w15515 and not w15516;
w15518 <= not w15514 and w15517;
w15519 <= w257 and w13514;
w15520 <= w15518 and not w15519;
w15521 <= a(8) and not w15520;
w15522 <= a(8) and not w15521;
w15523 <= not w15520 and not w15521;
w15524 <= not w15522 and not w15523;
w15525 <= not w15513 and not w15524;
w15526 <= not w15513 and not w15525;
w15527 <= not w15524 and not w15525;
w15528 <= not w15526 and not w15527;
w15529 <= b(60) and w443;
w15530 <= b(58) and w510;
w15531 <= b(59) and w438;
w15532 <= not w15530 and not w15531;
w15533 <= not w15529 and w15532;
w15534 <= w446 and w11954;
w15535 <= w15533 and not w15534;
w15536 <= a(11) and not w15535;
w15537 <= a(11) and not w15536;
w15538 <= not w15535 and not w15536;
w15539 <= not w15537 and not w15538;
w15540 <= not w15147 and not w15476;
w15541 <= w15539 and w15540;
w15542 <= not w15539 and not w15540;
w15543 <= not w15541 and not w15542;
w15544 <= not w15178 and not w15469;
w15545 <= b(54) and w1045;
w15546 <= b(52) and w1134;
w15547 <= b(53) and w1040;
w15548 <= not w15546 and not w15547;
w15549 <= not w15545 and w15548;
w15550 <= w1048 and w9741;
w15551 <= w15549 and not w15550;
w15552 <= a(17) and not w15551;
w15553 <= a(17) and not w15552;
w15554 <= not w15551 and not w15552;
w15555 <= not w15553 and not w15554;
w15556 <= not w15544 and not w15555;
w15557 <= not w15544 and not w15556;
w15558 <= not w15555 and not w15556;
w15559 <= not w15557 and not w15558;
w15560 <= b(48) and w1791;
w15561 <= b(46) and w1941;
w15562 <= b(47) and w1786;
w15563 <= not w15561 and not w15562;
w15564 <= not w15560 and w15563;
w15565 <= w1794 and w7752;
w15566 <= w15564 and not w15565;
w15567 <= a(23) and not w15566;
w15568 <= a(23) and not w15567;
w15569 <= not w15566 and not w15567;
w15570 <= not w15568 and not w15569;
w15571 <= not w15211 and not w15462;
w15572 <= w15570 and w15571;
w15573 <= not w15570 and not w15571;
w15574 <= not w15572 and not w15573;
w15575 <= not w15454 and not w15458;
w15576 <= b(45) and w2282;
w15577 <= b(43) and w2428;
w15578 <= b(44) and w2277;
w15579 <= not w15577 and not w15578;
w15580 <= not w15576 and w15579;
w15581 <= w2285 and w7104;
w15582 <= w15580 and not w15581;
w15583 <= a(26) and not w15582;
w15584 <= a(26) and not w15583;
w15585 <= not w15582 and not w15583;
w15586 <= not w15584 and not w15585;
w15587 <= not w15575 and not w15586;
w15588 <= not w15575 and not w15587;
w15589 <= not w15586 and not w15587;
w15590 <= not w15588 and not w15589;
w15591 <= b(42) and w2793;
w15592 <= b(40) and w2986;
w15593 <= b(41) and w2788;
w15594 <= not w15592 and not w15593;
w15595 <= not w15591 and w15594;
w15596 <= w2796 and w6232;
w15597 <= w15595 and not w15596;
w15598 <= a(29) and not w15597;
w15599 <= a(29) and not w15598;
w15600 <= not w15597 and not w15598;
w15601 <= not w15599 and not w15600;
w15602 <= not w15226 and not w15438;
w15603 <= w15601 and w15602;
w15604 <= not w15601 and not w15602;
w15605 <= not w15603 and not w15604;
w15606 <= not w15412 and not w15415;
w15607 <= not w15395 and not w15409;
w15608 <= not w15376 and not w15389;
w15609 <= not w15348 and not w15351;
w15610 <= not w15331 and not w15345;
w15611 <= not w15285 and not w15299;
w15612 <= b(12) and w11274;
w15613 <= b(10) and w11639;
w15614 <= b(11) and w11269;
w15615 <= not w15613 and not w15614;
w15616 <= not w15612 and w15615;
w15617 <= w585 and w11277;
w15618 <= w15616 and not w15617;
w15619 <= a(59) and not w15618;
w15620 <= a(59) and not w15619;
w15621 <= not w15618 and not w15619;
w15622 <= not w15620 and not w15621;
w15623 <= not w15275 and not w15279;
w15624 <= b(5) and w13646;
w15625 <= b(6) and not w13231;
w15626 <= not w15624 and not w15625;
w15627 <= a(2) and not a(5);
w15628 <= not a(2) and a(5);
w15629 <= not w15627 and not w15628;
w15630 <= not w15626 and not w15629;
w15631 <= w15626 and w15629;
w15632 <= not w15630 and not w15631;
w15633 <= w15623 and not w15632;
w15634 <= not w15623 and w15632;
w15635 <= not w15633 and not w15634;
w15636 <= b(9) and w12411;
w15637 <= b(7) and w12790;
w15638 <= b(8) and w12406;
w15639 <= not w15637 and not w15638;
w15640 <= not w15636 and w15639;
w15641 <= w394 and w12414;
w15642 <= w15640 and not w15641;
w15643 <= a(62) and not w15642;
w15644 <= a(62) and not w15643;
w15645 <= not w15642 and not w15643;
w15646 <= not w15644 and not w15645;
w15647 <= not w15635 and w15646;
w15648 <= w15635 and not w15646;
w15649 <= not w15647 and not w15648;
w15650 <= not w15622 and w15649;
w15651 <= not w15622 and not w15650;
w15652 <= w15649 and not w15650;
w15653 <= not w15651 and not w15652;
w15654 <= not w15611 and not w15653;
w15655 <= not w15611 and not w15654;
w15656 <= not w15653 and not w15654;
w15657 <= not w15655 and not w15656;
w15658 <= b(15) and w10169;
w15659 <= b(13) and w10539;
w15660 <= b(14) and w10164;
w15661 <= not w15659 and not w15660;
w15662 <= not w15658 and w15661;
w15663 <= w874 and w10172;
w15664 <= w15662 and not w15663;
w15665 <= a(56) and not w15664;
w15666 <= a(56) and not w15665;
w15667 <= not w15664 and not w15665;
w15668 <= not w15666 and not w15667;
w15669 <= not w15657 and not w15668;
w15670 <= not w15657 and not w15669;
w15671 <= not w15668 and not w15669;
w15672 <= not w15670 and not w15671;
w15673 <= not w15302 and not w15305;
w15674 <= w15672 and w15673;
w15675 <= not w15672 and not w15673;
w15676 <= not w15674 and not w15675;
w15677 <= b(18) and w9082;
w15678 <= b(16) and w9475;
w15679 <= b(17) and w9077;
w15680 <= not w15678 and not w15679;
w15681 <= not w15677 and w15680;
w15682 <= w1309 and w9085;
w15683 <= w15681 and not w15682;
w15684 <= a(53) and not w15683;
w15685 <= a(53) and not w15684;
w15686 <= not w15683 and not w15684;
w15687 <= not w15685 and not w15686;
w15688 <= w15676 and not w15687;
w15689 <= w15676 and not w15688;
w15690 <= not w15687 and not w15688;
w15691 <= not w15689 and not w15690;
w15692 <= not w15310 and not w15325;
w15693 <= w15691 and w15692;
w15694 <= not w15691 and not w15692;
w15695 <= not w15693 and not w15694;
w15696 <= b(21) and w8105;
w15697 <= b(19) and w8458;
w15698 <= b(20) and w8100;
w15699 <= not w15697 and not w15698;
w15700 <= not w15696 and w15699;
w15701 <= w1727 and w8108;
w15702 <= w15700 and not w15701;
w15703 <= a(50) and not w15702;
w15704 <= a(50) and not w15703;
w15705 <= not w15702 and not w15703;
w15706 <= not w15704 and not w15705;
w15707 <= w15695 and not w15706;
w15708 <= w15695 and not w15707;
w15709 <= not w15706 and not w15707;
w15710 <= not w15708 and not w15709;
w15711 <= not w15610 and w15710;
w15712 <= w15610 and not w15710;
w15713 <= not w15711 and not w15712;
w15714 <= b(24) and w7189;
w15715 <= b(22) and w7530;
w15716 <= b(23) and w7184;
w15717 <= not w15715 and not w15716;
w15718 <= not w15714 and w15717;
w15719 <= w2201 and w7192;
w15720 <= w15718 and not w15719;
w15721 <= a(47) and not w15720;
w15722 <= a(47) and not w15721;
w15723 <= not w15720 and not w15721;
w15724 <= not w15722 and not w15723;
w15725 <= not w15713 and not w15724;
w15726 <= w15713 and w15724;
w15727 <= not w15725 and not w15726;
w15728 <= w15609 and not w15727;
w15729 <= not w15609 and w15727;
w15730 <= not w15728 and not w15729;
w15731 <= b(27) and w6338;
w15732 <= b(25) and w6645;
w15733 <= b(26) and w6333;
w15734 <= not w15732 and not w15733;
w15735 <= not w15731 and w15734;
w15736 <= w2733 and w6341;
w15737 <= w15735 and not w15736;
w15738 <= a(44) and not w15737;
w15739 <= a(44) and not w15738;
w15740 <= not w15737 and not w15738;
w15741 <= not w15739 and not w15740;
w15742 <= w15730 and not w15741;
w15743 <= w15730 and not w15742;
w15744 <= not w15741 and not w15742;
w15745 <= not w15743 and not w15744;
w15746 <= not w15357 and not w15370;
w15747 <= w15745 and w15746;
w15748 <= not w15745 and not w15746;
w15749 <= not w15747 and not w15748;
w15750 <= b(30) and w5520;
w15751 <= b(28) and w5802;
w15752 <= b(29) and w5515;
w15753 <= not w15751 and not w15752;
w15754 <= not w15750 and w15753;
w15755 <= w3320 and w5523;
w15756 <= w15754 and not w15755;
w15757 <= a(41) and not w15756;
w15758 <= a(41) and not w15757;
w15759 <= not w15756 and not w15757;
w15760 <= not w15758 and not w15759;
w15761 <= w15749 and not w15760;
w15762 <= not w15749 and w15760;
w15763 <= not w15608 and not w15762;
w15764 <= not w15761 and w15763;
w15765 <= not w15608 and not w15764;
w15766 <= not w15761 and not w15764;
w15767 <= not w15762 and w15766;
w15768 <= not w15765 and not w15767;
w15769 <= b(33) and w4778;
w15770 <= b(31) and w5020;
w15771 <= b(32) and w4773;
w15772 <= not w15770 and not w15771;
w15773 <= not w15769 and w15772;
w15774 <= w3966 and w4781;
w15775 <= w15773 and not w15774;
w15776 <= a(38) and not w15775;
w15777 <= a(38) and not w15776;
w15778 <= not w15775 and not w15776;
w15779 <= not w15777 and not w15778;
w15780 <= not w15768 and not w15779;
w15781 <= not w15768 and not w15780;
w15782 <= not w15779 and not w15780;
w15783 <= not w15781 and not w15782;
w15784 <= not w15607 and w15783;
w15785 <= w15607 and not w15783;
w15786 <= not w15784 and not w15785;
w15787 <= b(36) and w4030;
w15788 <= b(34) and w4275;
w15789 <= b(35) and w4025;
w15790 <= not w15788 and not w15789;
w15791 <= not w15787 and w15790;
w15792 <= w4033 and w4665;
w15793 <= w15791 and not w15792;
w15794 <= a(35) and not w15793;
w15795 <= a(35) and not w15794;
w15796 <= not w15793 and not w15794;
w15797 <= not w15795 and not w15796;
w15798 <= not w15786 and not w15797;
w15799 <= w15786 and w15797;
w15800 <= not w15798 and not w15799;
w15801 <= w15606 and not w15800;
w15802 <= not w15606 and w15800;
w15803 <= not w15801 and not w15802;
w15804 <= b(39) and w3381;
w15805 <= b(37) and w3586;
w15806 <= b(38) and w3376;
w15807 <= not w15805 and not w15806;
w15808 <= not w15804 and w15807;
w15809 <= w3384 and w5194;
w15810 <= w15808 and not w15809;
w15811 <= a(32) and not w15810;
w15812 <= a(32) and not w15811;
w15813 <= not w15810 and not w15811;
w15814 <= not w15812 and not w15813;
w15815 <= not w15431 and not w15434;
w15816 <= w15814 and w15815;
w15817 <= not w15814 and not w15815;
w15818 <= not w15816 and not w15817;
w15819 <= w15803 and w15818;
w15820 <= not w15803 and not w15818;
w15821 <= not w15819 and not w15820;
w15822 <= w15605 and w15821;
w15823 <= not w15605 and not w15821;
w15824 <= not w15822 and not w15823;
w15825 <= not w15590 and not w15824;
w15826 <= w15590 and w15824;
w15827 <= not w15825 and not w15826;
w15828 <= w15574 and not w15827;
w15829 <= w15574 and not w15828;
w15830 <= not w15827 and not w15828;
w15831 <= not w15829 and not w15830;
w15832 <= b(51) and w1370;
w15833 <= b(49) and w1506;
w15834 <= b(50) and w1365;
w15835 <= not w15833 and not w15834;
w15836 <= not w15832 and w15835;
w15837 <= w1373 and w8719;
w15838 <= w15836 and not w15837;
w15839 <= a(20) and not w15838;
w15840 <= a(20) and not w15839;
w15841 <= not w15838 and not w15839;
w15842 <= not w15840 and not w15841;
w15843 <= not w15197 and not w15465;
w15844 <= not w15194 and not w15843;
w15845 <= not w15842 and not w15844;
w15846 <= w15842 and w15844;
w15847 <= not w15845 and not w15846;
w15848 <= not w15831 and w15847;
w15849 <= not w15831 and not w15848;
w15850 <= w15847 and not w15848;
w15851 <= not w15849 and not w15850;
w15852 <= not w15559 and not w15851;
w15853 <= not w15559 and not w15852;
w15854 <= not w15851 and not w15852;
w15855 <= not w15853 and not w15854;
w15856 <= b(57) and w694;
w15857 <= b(55) and w799;
w15858 <= b(56) and w689;
w15859 <= not w15857 and not w15858;
w15860 <= not w15856 and w15859;
w15861 <= w697 and w11153;
w15862 <= w15860 and not w15861;
w15863 <= a(14) and not w15862;
w15864 <= a(14) and not w15863;
w15865 <= not w15862 and not w15863;
w15866 <= not w15864 and not w15865;
w15867 <= not w15165 and not w15472;
w15868 <= not w15162 and not w15867;
w15869 <= not w15866 and not w15868;
w15870 <= w15866 and w15868;
w15871 <= not w15869 and not w15870;
w15872 <= not w15855 and w15871;
w15873 <= not w15855 and not w15872;
w15874 <= w15871 and not w15872;
w15875 <= not w15873 and not w15874;
w15876 <= w15543 and not w15875;
w15877 <= w15543 and not w15876;
w15878 <= not w15875 and not w15876;
w15879 <= not w15877 and not w15878;
w15880 <= not w15528 and w15879;
w15881 <= w15528 and not w15879;
w15882 <= not w15880 and not w15881;
w15883 <= not w15512 and not w15882;
w15884 <= w15512 and w15882;
w15885 <= not w15883 and not w15884;
w15886 <= not w15511 and w15885;
w15887 <= w15511 and not w15885;
w15888 <= not w15886 and not w15887;
w15889 <= not w15542 and not w15876;
w15890 <= b(62) and w284;
w15891 <= b(63) and w249;
w15892 <= not w15890 and not w15891;
w15893 <= not w257 and w15892;
w15894 <= w13543 and w15892;
w15895 <= not w15893 and not w15894;
w15896 <= a(8) and not w15895;
w15897 <= not a(8) and w15895;
w15898 <= not w15896 and not w15897;
w15899 <= not w15889 and not w15898;
w15900 <= w15889 and w15898;
w15901 <= not w15899 and not w15900;
w15902 <= b(61) and w443;
w15903 <= b(59) and w510;
w15904 <= b(60) and w438;
w15905 <= not w15903 and not w15904;
w15906 <= not w15902 and w15905;
w15907 <= w446 and w12712;
w15908 <= w15906 and not w15907;
w15909 <= a(11) and not w15908;
w15910 <= a(11) and not w15909;
w15911 <= not w15908 and not w15909;
w15912 <= not w15910 and not w15911;
w15913 <= not w15869 and not w15872;
w15914 <= w15912 and w15913;
w15915 <= not w15912 and not w15913;
w15916 <= not w15914 and not w15915;
w15917 <= not w15556 and not w15852;
w15918 <= b(58) and w694;
w15919 <= b(56) and w799;
w15920 <= b(57) and w689;
w15921 <= not w15919 and not w15920;
w15922 <= not w15918 and w15921;
w15923 <= not w697 and w15922;
w15924 <= not w11179 and w15922;
w15925 <= not w15923 and not w15924;
w15926 <= a(14) and not w15925;
w15927 <= not a(14) and w15925;
w15928 <= not w15926 and not w15927;
w15929 <= not w15917 and not w15928;
w15930 <= w15917 and w15928;
w15931 <= not w15929 and not w15930;
w15932 <= b(55) and w1045;
w15933 <= b(53) and w1134;
w15934 <= b(54) and w1040;
w15935 <= not w15933 and not w15934;
w15936 <= not w15932 and w15935;
w15937 <= w1048 and w10427;
w15938 <= w15936 and not w15937;
w15939 <= a(17) and not w15938;
w15940 <= a(17) and not w15939;
w15941 <= not w15938 and not w15939;
w15942 <= not w15940 and not w15941;
w15943 <= not w15845 and not w15848;
w15944 <= w15942 and w15943;
w15945 <= not w15942 and not w15943;
w15946 <= not w15944 and not w15945;
w15947 <= b(52) and w1370;
w15948 <= b(50) and w1506;
w15949 <= b(51) and w1365;
w15950 <= not w15948 and not w15949;
w15951 <= not w15947 and w15950;
w15952 <= w1373 and w9371;
w15953 <= w15951 and not w15952;
w15954 <= a(20) and not w15953;
w15955 <= a(20) and not w15954;
w15956 <= not w15953 and not w15954;
w15957 <= not w15955 and not w15956;
w15958 <= not w15573 and not w15828;
w15959 <= w15957 and w15958;
w15960 <= not w15957 and not w15958;
w15961 <= not w15959 and not w15960;
w15962 <= b(49) and w1791;
w15963 <= b(47) and w1941;
w15964 <= b(48) and w1786;
w15965 <= not w15963 and not w15964;
w15966 <= not w15962 and w15965;
w15967 <= w1794 and w8368;
w15968 <= w15966 and not w15967;
w15969 <= a(23) and not w15968;
w15970 <= a(23) and not w15969;
w15971 <= not w15968 and not w15969;
w15972 <= not w15970 and not w15971;
w15973 <= not w15590 and w15824;
w15974 <= not w15587 and not w15973;
w15975 <= not w15972 and not w15974;
w15976 <= not w15972 and not w15975;
w15977 <= not w15974 and not w15975;
w15978 <= not w15976 and not w15977;
w15979 <= not w15604 and not w15822;
w15980 <= b(46) and w2282;
w15981 <= b(44) and w2428;
w15982 <= b(45) and w2277;
w15983 <= not w15981 and not w15982;
w15984 <= not w15980 and w15983;
w15985 <= not w2285 and w15984;
w15986 <= not w7420 and w15984;
w15987 <= not w15985 and not w15986;
w15988 <= a(26) and not w15987;
w15989 <= not a(26) and w15987;
w15990 <= not w15988 and not w15989;
w15991 <= not w15979 and not w15990;
w15992 <= w15979 and w15990;
w15993 <= not w15991 and not w15992;
w15994 <= b(43) and w2793;
w15995 <= b(41) and w2986;
w15996 <= b(42) and w2788;
w15997 <= not w15995 and not w15996;
w15998 <= not w15994 and w15997;
w15999 <= w2796 and w6258;
w16000 <= w15998 and not w15999;
w16001 <= a(29) and not w16000;
w16002 <= a(29) and not w16001;
w16003 <= not w16000 and not w16001;
w16004 <= not w16002 and not w16003;
w16005 <= not w15817 and not w15819;
w16006 <= not w16004 and not w16005;
w16007 <= not w16004 and not w16006;
w16008 <= not w16005 and not w16006;
w16009 <= not w16007 and not w16008;
w16010 <= b(40) and w3381;
w16011 <= b(38) and w3586;
w16012 <= b(39) and w3376;
w16013 <= not w16011 and not w16012;
w16014 <= not w16010 and w16013;
w16015 <= w3384 and w5698;
w16016 <= w16014 and not w16015;
w16017 <= a(32) and not w16016;
w16018 <= a(32) and not w16017;
w16019 <= not w16016 and not w16017;
w16020 <= not w16018 and not w16019;
w16021 <= not w15798 and not w15802;
w16022 <= w16020 and w16021;
w16023 <= not w16020 and not w16021;
w16024 <= not w16022 and not w16023;
w16025 <= b(37) and w4030;
w16026 <= b(35) and w4275;
w16027 <= b(36) and w4025;
w16028 <= not w16026 and not w16027;
w16029 <= not w16025 and w16028;
w16030 <= w4033 and w4924;
w16031 <= w16029 and not w16030;
w16032 <= a(35) and not w16031;
w16033 <= a(35) and not w16032;
w16034 <= not w16031 and not w16032;
w16035 <= not w16033 and not w16034;
w16036 <= not w15607 and not w15783;
w16037 <= not w15780 and not w16036;
w16038 <= b(34) and w4778;
w16039 <= b(32) and w5020;
w16040 <= b(33) and w4773;
w16041 <= not w16039 and not w16040;
w16042 <= not w16038 and w16041;
w16043 <= w4209 and w4781;
w16044 <= w16042 and not w16043;
w16045 <= a(38) and not w16044;
w16046 <= a(38) and not w16045;
w16047 <= not w16044 and not w16045;
w16048 <= not w16046 and not w16047;
w16049 <= not w15634 and not w15648;
w16050 <= not a(2) and not a(5);
w16051 <= not w15630 and not w16050;
w16052 <= b(6) and w13646;
w16053 <= b(7) and not w13231;
w16054 <= not w16052 and not w16053;
w16055 <= not w16051 and w16054;
w16056 <= w16051 and not w16054;
w16057 <= not w16055 and not w16056;
w16058 <= b(10) and w12411;
w16059 <= b(8) and w12790;
w16060 <= b(9) and w12406;
w16061 <= not w16059 and not w16060;
w16062 <= not w16058 and w16061;
w16063 <= not w12414 and w16062;
w16064 <= not w481 and w16062;
w16065 <= not w16063 and not w16064;
w16066 <= a(62) and not w16065;
w16067 <= not a(62) and w16065;
w16068 <= not w16066 and not w16067;
w16069 <= w16057 and not w16068;
w16070 <= not w16057 and w16068;
w16071 <= not w16069 and not w16070;
w16072 <= not w16049 and w16071;
w16073 <= w16049 and not w16071;
w16074 <= not w16072 and not w16073;
w16075 <= b(13) and w11274;
w16076 <= b(11) and w11639;
w16077 <= b(12) and w11269;
w16078 <= not w16076 and not w16077;
w16079 <= not w16075 and w16078;
w16080 <= w751 and w11277;
w16081 <= w16079 and not w16080;
w16082 <= a(59) and not w16081;
w16083 <= a(59) and not w16082;
w16084 <= not w16081 and not w16082;
w16085 <= not w16083 and not w16084;
w16086 <= w16074 and not w16085;
w16087 <= w16074 and not w16086;
w16088 <= not w16085 and not w16086;
w16089 <= not w16087 and not w16088;
w16090 <= not w15650 and not w15654;
w16091 <= w16089 and w16090;
w16092 <= not w16089 and not w16090;
w16093 <= not w16091 and not w16092;
w16094 <= b(16) and w10169;
w16095 <= b(14) and w10539;
w16096 <= b(15) and w10164;
w16097 <= not w16095 and not w16096;
w16098 <= not w16094 and w16097;
w16099 <= w980 and w10172;
w16100 <= w16098 and not w16099;
w16101 <= a(56) and not w16100;
w16102 <= a(56) and not w16101;
w16103 <= not w16100 and not w16101;
w16104 <= not w16102 and not w16103;
w16105 <= w16093 and not w16104;
w16106 <= w16093 and not w16105;
w16107 <= not w16104 and not w16105;
w16108 <= not w16106 and not w16107;
w16109 <= not w15669 and not w15675;
w16110 <= w16108 and w16109;
w16111 <= not w16108 and not w16109;
w16112 <= not w16110 and not w16111;
w16113 <= b(19) and w9082;
w16114 <= b(17) and w9475;
w16115 <= b(18) and w9077;
w16116 <= not w16114 and not w16115;
w16117 <= not w16113 and w16116;
w16118 <= w1451 and w9085;
w16119 <= w16117 and not w16118;
w16120 <= a(53) and not w16119;
w16121 <= a(53) and not w16120;
w16122 <= not w16119 and not w16120;
w16123 <= not w16121 and not w16122;
w16124 <= w16112 and not w16123;
w16125 <= w16112 and not w16124;
w16126 <= not w16123 and not w16124;
w16127 <= not w16125 and not w16126;
w16128 <= not w15688 and not w15694;
w16129 <= w16127 and w16128;
w16130 <= not w16127 and not w16128;
w16131 <= not w16129 and not w16130;
w16132 <= b(22) and w8105;
w16133 <= b(20) and w8458;
w16134 <= b(21) and w8100;
w16135 <= not w16133 and not w16134;
w16136 <= not w16132 and w16135;
w16137 <= w1888 and w8108;
w16138 <= w16136 and not w16137;
w16139 <= a(50) and not w16138;
w16140 <= a(50) and not w16139;
w16141 <= not w16138 and not w16139;
w16142 <= not w16140 and not w16141;
w16143 <= w16131 and not w16142;
w16144 <= w16131 and not w16143;
w16145 <= not w16142 and not w16143;
w16146 <= not w16144 and not w16145;
w16147 <= not w15610 and not w15710;
w16148 <= not w15707 and not w16147;
w16149 <= w16146 and w16148;
w16150 <= not w16146 and not w16148;
w16151 <= not w16149 and not w16150;
w16152 <= b(25) and w7189;
w16153 <= b(23) and w7530;
w16154 <= b(24) and w7184;
w16155 <= not w16153 and not w16154;
w16156 <= not w16152 and w16155;
w16157 <= w2228 and w7192;
w16158 <= w16156 and not w16157;
w16159 <= a(47) and not w16158;
w16160 <= a(47) and not w16159;
w16161 <= not w16158 and not w16159;
w16162 <= not w16160 and not w16161;
w16163 <= w16151 and not w16162;
w16164 <= w16151 and not w16163;
w16165 <= not w16162 and not w16163;
w16166 <= not w16164 and not w16165;
w16167 <= not w15725 and not w15729;
w16168 <= w16166 and w16167;
w16169 <= not w16166 and not w16167;
w16170 <= not w16168 and not w16169;
w16171 <= b(28) and w6338;
w16172 <= b(26) and w6645;
w16173 <= b(27) and w6333;
w16174 <= not w16172 and not w16173;
w16175 <= not w16171 and w16174;
w16176 <= w2932 and w6341;
w16177 <= w16175 and not w16176;
w16178 <= a(44) and not w16177;
w16179 <= a(44) and not w16178;
w16180 <= not w16177 and not w16178;
w16181 <= not w16179 and not w16180;
w16182 <= w16170 and not w16181;
w16183 <= w16170 and not w16182;
w16184 <= not w16181 and not w16182;
w16185 <= not w16183 and not w16184;
w16186 <= not w15742 and not w15748;
w16187 <= w16185 and w16186;
w16188 <= not w16185 and not w16186;
w16189 <= not w16187 and not w16188;
w16190 <= b(31) and w5520;
w16191 <= b(29) and w5802;
w16192 <= b(30) and w5515;
w16193 <= not w16191 and not w16192;
w16194 <= not w16190 and w16193;
w16195 <= w3539 and w5523;
w16196 <= w16194 and not w16195;
w16197 <= a(41) and not w16196;
w16198 <= a(41) and not w16197;
w16199 <= not w16196 and not w16197;
w16200 <= not w16198 and not w16199;
w16201 <= not w16189 and w16200;
w16202 <= w16189 and not w16200;
w16203 <= not w16201 and not w16202;
w16204 <= not w15766 and w16203;
w16205 <= w15766 and not w16203;
w16206 <= not w16204 and not w16205;
w16207 <= not w16048 and w16206;
w16208 <= w16048 and not w16206;
w16209 <= not w16207 and not w16208;
w16210 <= not w16037 and w16209;
w16211 <= w16037 and not w16209;
w16212 <= not w16210 and not w16211;
w16213 <= not w16035 and w16212;
w16214 <= not w16035 and not w16213;
w16215 <= w16212 and not w16213;
w16216 <= not w16214 and not w16215;
w16217 <= w16024 and not w16216;
w16218 <= w16024 and not w16217;
w16219 <= not w16216 and not w16217;
w16220 <= not w16218 and not w16219;
w16221 <= not w16009 and w16220;
w16222 <= w16009 and not w16220;
w16223 <= not w16221 and not w16222;
w16224 <= w15993 and not w16223;
w16225 <= w15993 and not w16224;
w16226 <= not w16223 and not w16224;
w16227 <= not w16225 and not w16226;
w16228 <= not w15978 and w16227;
w16229 <= w15978 and not w16227;
w16230 <= not w16228 and not w16229;
w16231 <= w15961 and not w16230;
w16232 <= w15961 and not w16231;
w16233 <= not w16230 and not w16231;
w16234 <= not w16232 and not w16233;
w16235 <= w15946 and not w16234;
w16236 <= not w15946 and w16234;
w16237 <= w15931 and not w16236;
w16238 <= not w16235 and w16237;
w16239 <= w15931 and not w16238;
w16240 <= not w16236 and not w16238;
w16241 <= not w16235 and w16240;
w16242 <= not w16239 and not w16241;
w16243 <= w15916 and not w16242;
w16244 <= not w15916 and w16242;
w16245 <= w15901 and not w16244;
w16246 <= not w16243 and w16245;
w16247 <= w15901 and not w16246;
w16248 <= not w16244 and not w16246;
w16249 <= not w16243 and w16248;
w16250 <= not w16247 and not w16249;
w16251 <= not w15528 and not w15879;
w16252 <= not w15525 and not w16251;
w16253 <= not w16250 and not w16252;
w16254 <= not w16250 and not w16253;
w16255 <= not w16252 and not w16253;
w16256 <= not w16254 and not w16255;
w16257 <= not w15883 and not w15886;
w16258 <= not w16256 and not w16257;
w16259 <= w16256 and w16257;
w16260 <= not w16258 and not w16259;
w16261 <= not w16253 and not w16258;
w16262 <= not w15899 and not w16246;
w16263 <= not w15915 and not w16243;
w16264 <= b(63) and w284;
w16265 <= w257 and w13540;
w16266 <= not w16264 and not w16265;
w16267 <= a(8) and not w16266;
w16268 <= a(8) and not w16267;
w16269 <= not w16266 and not w16267;
w16270 <= not w16268 and not w16269;
w16271 <= not w16263 and not w16270;
w16272 <= not w16263 and not w16271;
w16273 <= not w16270 and not w16271;
w16274 <= not w16272 and not w16273;
w16275 <= b(56) and w1045;
w16276 <= b(54) and w1134;
w16277 <= b(55) and w1040;
w16278 <= not w16276 and not w16277;
w16279 <= not w16275 and w16278;
w16280 <= w1048 and w10451;
w16281 <= w16279 and not w16280;
w16282 <= a(17) and not w16281;
w16283 <= a(17) and not w16282;
w16284 <= not w16281 and not w16282;
w16285 <= not w16283 and not w16284;
w16286 <= not w15960 and not w16231;
w16287 <= w16285 and w16286;
w16288 <= not w16285 and not w16286;
w16289 <= not w16287 and not w16288;
w16290 <= b(50) and w1791;
w16291 <= b(48) and w1941;
w16292 <= b(49) and w1786;
w16293 <= not w16291 and not w16292;
w16294 <= not w16290 and w16293;
w16295 <= w1794 and w8692;
w16296 <= w16294 and not w16295;
w16297 <= a(23) and not w16296;
w16298 <= a(23) and not w16297;
w16299 <= not w16296 and not w16297;
w16300 <= not w16298 and not w16299;
w16301 <= not w15991 and not w16224;
w16302 <= w16300 and w16301;
w16303 <= not w16300 and not w16301;
w16304 <= not w16302 and not w16303;
w16305 <= b(47) and w2282;
w16306 <= b(45) and w2428;
w16307 <= b(46) and w2277;
w16308 <= not w16306 and not w16307;
w16309 <= not w16305 and w16308;
w16310 <= w2285 and w7446;
w16311 <= w16309 and not w16310;
w16312 <= a(26) and not w16311;
w16313 <= a(26) and not w16312;
w16314 <= not w16311 and not w16312;
w16315 <= not w16313 and not w16314;
w16316 <= not w16009 and not w16220;
w16317 <= not w16006 and not w16316;
w16318 <= not w16315 and not w16317;
w16319 <= not w16315 and not w16318;
w16320 <= not w16317 and not w16318;
w16321 <= not w16319 and not w16320;
w16322 <= b(41) and w3381;
w16323 <= b(39) and w3586;
w16324 <= b(40) and w3376;
w16325 <= not w16323 and not w16324;
w16326 <= not w16322 and w16325;
w16327 <= w3384 and w5962;
w16328 <= w16326 and not w16327;
w16329 <= a(32) and not w16328;
w16330 <= a(32) and not w16329;
w16331 <= not w16328 and not w16329;
w16332 <= not w16330 and not w16331;
w16333 <= not w16210 and not w16213;
w16334 <= w16332 and w16333;
w16335 <= not w16332 and not w16333;
w16336 <= not w16334 and not w16335;
w16337 <= b(35) and w4778;
w16338 <= b(33) and w5020;
w16339 <= b(34) and w4773;
w16340 <= not w16338 and not w16339;
w16341 <= not w16337 and w16340;
w16342 <= w4439 and w4781;
w16343 <= w16341 and not w16342;
w16344 <= a(38) and not w16343;
w16345 <= a(38) and not w16344;
w16346 <= not w16343 and not w16344;
w16347 <= not w16345 and not w16346;
w16348 <= b(26) and w7189;
w16349 <= b(24) and w7530;
w16350 <= b(25) and w7184;
w16351 <= not w16349 and not w16350;
w16352 <= not w16348 and w16351;
w16353 <= w2556 and w7192;
w16354 <= w16352 and not w16353;
w16355 <= a(47) and not w16354;
w16356 <= a(47) and not w16355;
w16357 <= not w16354 and not w16355;
w16358 <= not w16356 and not w16357;
w16359 <= not w16130 and not w16143;
w16360 <= b(23) and w8105;
w16361 <= b(21) and w8458;
w16362 <= b(22) and w8100;
w16363 <= not w16361 and not w16362;
w16364 <= not w16360 and w16363;
w16365 <= w2043 and w8108;
w16366 <= w16364 and not w16365;
w16367 <= a(50) and not w16366;
w16368 <= a(50) and not w16367;
w16369 <= not w16366 and not w16367;
w16370 <= not w16368 and not w16369;
w16371 <= not w16111 and not w16124;
w16372 <= not w16072 and not w16086;
w16373 <= not w16055 and not w16069;
w16374 <= b(7) and w13646;
w16375 <= b(8) and not w13231;
w16376 <= not w16374 and not w16375;
w16377 <= w16054 and not w16376;
w16378 <= not w16054 and w16376;
w16379 <= not w16373 and not w16378;
w16380 <= not w16377 and w16379;
w16381 <= not w16373 and not w16380;
w16382 <= not w16378 and not w16380;
w16383 <= not w16377 and w16382;
w16384 <= not w16381 and not w16383;
w16385 <= b(11) and w12411;
w16386 <= b(9) and w12790;
w16387 <= b(10) and w12406;
w16388 <= not w16386 and not w16387;
w16389 <= not w16385 and w16388;
w16390 <= w561 and w12414;
w16391 <= w16389 and not w16390;
w16392 <= a(62) and not w16391;
w16393 <= a(62) and not w16392;
w16394 <= not w16391 and not w16392;
w16395 <= not w16393 and not w16394;
w16396 <= not w16384 and w16395;
w16397 <= w16384 and not w16395;
w16398 <= not w16396 and not w16397;
w16399 <= b(14) and w11274;
w16400 <= b(12) and w11639;
w16401 <= b(13) and w11269;
w16402 <= not w16400 and not w16401;
w16403 <= not w16399 and w16402;
w16404 <= w777 and w11277;
w16405 <= w16403 and not w16404;
w16406 <= a(59) and not w16405;
w16407 <= a(59) and not w16406;
w16408 <= not w16405 and not w16406;
w16409 <= not w16407 and not w16408;
w16410 <= not w16398 and not w16409;
w16411 <= w16398 and w16409;
w16412 <= not w16410 and not w16411;
w16413 <= w16372 and not w16412;
w16414 <= not w16372 and w16412;
w16415 <= not w16413 and not w16414;
w16416 <= b(17) and w10169;
w16417 <= b(15) and w10539;
w16418 <= b(16) and w10164;
w16419 <= not w16417 and not w16418;
w16420 <= not w16416 and w16419;
w16421 <= w1099 and w10172;
w16422 <= w16420 and not w16421;
w16423 <= a(56) and not w16422;
w16424 <= a(56) and not w16423;
w16425 <= not w16422 and not w16423;
w16426 <= not w16424 and not w16425;
w16427 <= w16415 and not w16426;
w16428 <= w16415 and not w16427;
w16429 <= not w16426 and not w16427;
w16430 <= not w16428 and not w16429;
w16431 <= not w16092 and not w16105;
w16432 <= w16430 and w16431;
w16433 <= not w16430 and not w16431;
w16434 <= not w16432 and not w16433;
w16435 <= b(20) and w9082;
w16436 <= b(18) and w9475;
w16437 <= b(19) and w9077;
w16438 <= not w16436 and not w16437;
w16439 <= not w16435 and w16438;
w16440 <= w1589 and w9085;
w16441 <= w16439 and not w16440;
w16442 <= a(53) and not w16441;
w16443 <= a(53) and not w16442;
w16444 <= not w16441 and not w16442;
w16445 <= not w16443 and not w16444;
w16446 <= not w16434 and w16445;
w16447 <= w16434 and not w16445;
w16448 <= not w16446 and not w16447;
w16449 <= not w16371 and w16448;
w16450 <= not w16371 and not w16449;
w16451 <= w16448 and not w16449;
w16452 <= not w16450 and not w16451;
w16453 <= not w16370 and not w16452;
w16454 <= w16370 and not w16451;
w16455 <= not w16450 and w16454;
w16456 <= not w16453 and not w16455;
w16457 <= not w16359 and w16456;
w16458 <= w16359 and not w16456;
w16459 <= not w16457 and not w16458;
w16460 <= not w16358 and w16459;
w16461 <= w16459 and not w16460;
w16462 <= not w16358 and not w16460;
w16463 <= not w16461 and not w16462;
w16464 <= not w16150 and not w16163;
w16465 <= w16463 and w16464;
w16466 <= not w16463 and not w16464;
w16467 <= not w16465 and not w16466;
w16468 <= b(29) and w6338;
w16469 <= b(27) and w6645;
w16470 <= b(28) and w6333;
w16471 <= not w16469 and not w16470;
w16472 <= not w16468 and w16471;
w16473 <= w3126 and w6341;
w16474 <= w16472 and not w16473;
w16475 <= a(44) and not w16474;
w16476 <= a(44) and not w16475;
w16477 <= not w16474 and not w16475;
w16478 <= not w16476 and not w16477;
w16479 <= w16467 and not w16478;
w16480 <= w16467 and not w16479;
w16481 <= not w16478 and not w16479;
w16482 <= not w16480 and not w16481;
w16483 <= not w16169 and not w16182;
w16484 <= w16482 and w16483;
w16485 <= not w16482 and not w16483;
w16486 <= not w16484 and not w16485;
w16487 <= b(32) and w5520;
w16488 <= b(30) and w5802;
w16489 <= b(31) and w5515;
w16490 <= not w16488 and not w16489;
w16491 <= not w16487 and w16490;
w16492 <= w3756 and w5523;
w16493 <= w16491 and not w16492;
w16494 <= a(41) and not w16493;
w16495 <= a(41) and not w16494;
w16496 <= not w16493 and not w16494;
w16497 <= not w16495 and not w16496;
w16498 <= not w16486 and w16497;
w16499 <= w16486 and not w16497;
w16500 <= not w16498 and not w16499;
w16501 <= not w16188 and not w16202;
w16502 <= w16500 and not w16501;
w16503 <= not w16500 and w16501;
w16504 <= not w16502 and not w16503;
w16505 <= not w16347 and w16504;
w16506 <= w16504 and not w16505;
w16507 <= not w16347 and not w16505;
w16508 <= not w16506 and not w16507;
w16509 <= not w16204 and not w16207;
w16510 <= w16508 and w16509;
w16511 <= not w16508 and not w16509;
w16512 <= not w16510 and not w16511;
w16513 <= b(38) and w4030;
w16514 <= b(36) and w4275;
w16515 <= b(37) and w4025;
w16516 <= not w16514 and not w16515;
w16517 <= not w16513 and w16516;
w16518 <= w4033 and w4948;
w16519 <= w16517 and not w16518;
w16520 <= a(35) and not w16519;
w16521 <= a(35) and not w16520;
w16522 <= not w16519 and not w16520;
w16523 <= not w16521 and not w16522;
w16524 <= w16512 and not w16523;
w16525 <= not w16512 and w16523;
w16526 <= w16336 and not w16525;
w16527 <= not w16524 and w16526;
w16528 <= w16336 and not w16527;
w16529 <= not w16525 and not w16527;
w16530 <= not w16524 and w16529;
w16531 <= not w16528 and not w16530;
w16532 <= not w16023 and not w16217;
w16533 <= b(44) and w2793;
w16534 <= b(42) and w2986;
w16535 <= b(43) and w2788;
w16536 <= not w16534 and not w16535;
w16537 <= not w16533 and w16536;
w16538 <= not w2796 and w16537;
w16539 <= not w6815 and w16537;
w16540 <= not w16538 and not w16539;
w16541 <= a(29) and not w16540;
w16542 <= not a(29) and w16540;
w16543 <= not w16541 and not w16542;
w16544 <= not w16532 and not w16543;
w16545 <= not w16532 and not w16544;
w16546 <= not w16543 and not w16544;
w16547 <= not w16545 and not w16546;
w16548 <= not w16531 and not w16547;
w16549 <= not w16531 and not w16548;
w16550 <= not w16547 and not w16548;
w16551 <= not w16549 and not w16550;
w16552 <= not w16321 and not w16551;
w16553 <= not w16321 and not w16552;
w16554 <= not w16551 and not w16552;
w16555 <= not w16553 and not w16554;
w16556 <= not w16304 and w16555;
w16557 <= w16304 and not w16555;
w16558 <= not w16556 and not w16557;
w16559 <= not w15978 and not w16227;
w16560 <= not w15975 and not w16559;
w16561 <= b(53) and w1370;
w16562 <= b(51) and w1506;
w16563 <= b(52) and w1365;
w16564 <= not w16562 and not w16563;
w16565 <= not w16561 and w16564;
w16566 <= not w1373 and w16565;
w16567 <= not w9715 and w16565;
w16568 <= not w16566 and not w16567;
w16569 <= a(20) and not w16568;
w16570 <= not a(20) and w16568;
w16571 <= not w16569 and not w16570;
w16572 <= not w16560 and not w16571;
w16573 <= not w16560 and not w16572;
w16574 <= not w16571 and not w16572;
w16575 <= not w16573 and not w16574;
w16576 <= w16558 and not w16575;
w16577 <= w16558 and not w16576;
w16578 <= not w16575 and not w16576;
w16579 <= not w16577 and not w16578;
w16580 <= w16289 and not w16579;
w16581 <= w16289 and not w16580;
w16582 <= not w16579 and not w16580;
w16583 <= not w16581 and not w16582;
w16584 <= b(59) and w694;
w16585 <= b(57) and w799;
w16586 <= b(58) and w689;
w16587 <= not w16585 and not w16586;
w16588 <= not w16584 and w16587;
w16589 <= w697 and w11922;
w16590 <= w16588 and not w16589;
w16591 <= a(14) and not w16590;
w16592 <= a(14) and not w16591;
w16593 <= not w16590 and not w16591;
w16594 <= not w16592 and not w16593;
w16595 <= not w15945 and not w16235;
w16596 <= not w16594 and not w16595;
w16597 <= not w16594 and not w16596;
w16598 <= not w16595 and not w16596;
w16599 <= not w16597 and not w16598;
w16600 <= not w16583 and w16599;
w16601 <= w16583 and not w16599;
w16602 <= not w16600 and not w16601;
w16603 <= not w15929 and not w16238;
w16604 <= b(62) and w443;
w16605 <= b(60) and w510;
w16606 <= b(61) and w438;
w16607 <= not w16605 and not w16606;
w16608 <= not w16604 and w16607;
w16609 <= not w446 and w16608;
w16610 <= not w13113 and w16608;
w16611 <= not w16609 and not w16610;
w16612 <= a(11) and not w16611;
w16613 <= not a(11) and w16611;
w16614 <= not w16612 and not w16613;
w16615 <= not w16603 and not w16614;
w16616 <= not w16603 and not w16615;
w16617 <= not w16614 and not w16615;
w16618 <= not w16616 and not w16617;
w16619 <= not w16602 and not w16618;
w16620 <= w16602 and not w16617;
w16621 <= not w16616 and w16620;
w16622 <= not w16619 and not w16621;
w16623 <= not w16274 and w16622;
w16624 <= w16274 and not w16622;
w16625 <= not w16623 and not w16624;
w16626 <= not w16262 and w16625;
w16627 <= not w16262 and not w16626;
w16628 <= w16625 and not w16626;
w16629 <= not w16627 and not w16628;
w16630 <= not w16261 and not w16629;
w16631 <= w16261 and not w16628;
w16632 <= not w16627 and w16631;
w16633 <= not w16630 and not w16632;
w16634 <= not w16626 and not w16630;
w16635 <= not w16271 and not w16623;
w16636 <= not w16615 and not w16619;
w16637 <= b(63) and w443;
w16638 <= b(61) and w510;
w16639 <= b(62) and w438;
w16640 <= not w16638 and not w16639;
w16641 <= not w16637 and w16640;
w16642 <= w446 and w13514;
w16643 <= w16641 and not w16642;
w16644 <= a(11) and not w16643;
w16645 <= a(11) and not w16644;
w16646 <= not w16643 and not w16644;
w16647 <= not w16645 and not w16646;
w16648 <= not w16636 and not w16647;
w16649 <= not w16636 and not w16648;
w16650 <= not w16647 and not w16648;
w16651 <= not w16649 and not w16650;
w16652 <= not w16583 and not w16599;
w16653 <= not w16596 and not w16652;
w16654 <= b(60) and w694;
w16655 <= b(58) and w799;
w16656 <= b(59) and w689;
w16657 <= not w16655 and not w16656;
w16658 <= not w16654 and w16657;
w16659 <= w697 and w11954;
w16660 <= w16658 and not w16659;
w16661 <= a(14) and not w16660;
w16662 <= a(14) and not w16661;
w16663 <= not w16660 and not w16661;
w16664 <= not w16662 and not w16663;
w16665 <= not w16653 and w16664;
w16666 <= w16653 and not w16664;
w16667 <= not w16665 and not w16666;
w16668 <= b(57) and w1045;
w16669 <= b(55) and w1134;
w16670 <= b(56) and w1040;
w16671 <= not w16669 and not w16670;
w16672 <= not w16668 and w16671;
w16673 <= w1048 and w11153;
w16674 <= w16672 and not w16673;
w16675 <= a(17) and not w16674;
w16676 <= a(17) and not w16675;
w16677 <= not w16674 and not w16675;
w16678 <= not w16676 and not w16677;
w16679 <= not w16288 and not w16580;
w16680 <= w16678 and w16679;
w16681 <= not w16678 and not w16679;
w16682 <= not w16680 and not w16681;
w16683 <= not w16572 and not w16576;
w16684 <= b(54) and w1370;
w16685 <= b(52) and w1506;
w16686 <= b(53) and w1365;
w16687 <= not w16685 and not w16686;
w16688 <= not w16684 and w16687;
w16689 <= w1373 and w9741;
w16690 <= w16688 and not w16689;
w16691 <= a(20) and not w16690;
w16692 <= a(20) and not w16691;
w16693 <= not w16690 and not w16691;
w16694 <= not w16692 and not w16693;
w16695 <= not w16683 and not w16694;
w16696 <= not w16683 and not w16695;
w16697 <= not w16694 and not w16695;
w16698 <= not w16696 and not w16697;
w16699 <= b(48) and w2282;
w16700 <= b(46) and w2428;
w16701 <= b(47) and w2277;
w16702 <= not w16700 and not w16701;
w16703 <= not w16699 and w16702;
w16704 <= w2285 and w7752;
w16705 <= w16703 and not w16704;
w16706 <= a(26) and not w16705;
w16707 <= a(26) and not w16706;
w16708 <= not w16705 and not w16706;
w16709 <= not w16707 and not w16708;
w16710 <= not w16318 and not w16552;
w16711 <= w16709 and w16710;
w16712 <= not w16709 and not w16710;
w16713 <= not w16711 and not w16712;
w16714 <= not w16544 and not w16548;
w16715 <= b(45) and w2793;
w16716 <= b(43) and w2986;
w16717 <= b(44) and w2788;
w16718 <= not w16716 and not w16717;
w16719 <= not w16715 and w16718;
w16720 <= w2796 and w7104;
w16721 <= w16719 and not w16720;
w16722 <= a(29) and not w16721;
w16723 <= a(29) and not w16722;
w16724 <= not w16721 and not w16722;
w16725 <= not w16723 and not w16724;
w16726 <= not w16714 and not w16725;
w16727 <= not w16714 and not w16726;
w16728 <= not w16725 and not w16726;
w16729 <= not w16727 and not w16728;
w16730 <= not w16335 and not w16527;
w16731 <= b(42) and w3381;
w16732 <= b(40) and w3586;
w16733 <= b(41) and w3376;
w16734 <= not w16732 and not w16733;
w16735 <= not w16731 and w16734;
w16736 <= w3384 and w6232;
w16737 <= w16735 and not w16736;
w16738 <= a(32) and not w16737;
w16739 <= a(32) and not w16738;
w16740 <= not w16737 and not w16738;
w16741 <= not w16739 and not w16740;
w16742 <= not w16730 and not w16741;
w16743 <= not w16730 and not w16742;
w16744 <= not w16741 and not w16742;
w16745 <= not w16743 and not w16744;
w16746 <= not w16502 and not w16505;
w16747 <= not w16485 and not w16499;
w16748 <= not w16466 and not w16479;
w16749 <= not w16449 and not w16453;
w16750 <= b(24) and w8105;
w16751 <= b(22) and w8458;
w16752 <= b(23) and w8100;
w16753 <= not w16751 and not w16752;
w16754 <= not w16750 and w16753;
w16755 <= w2201 and w8108;
w16756 <= w16754 and not w16755;
w16757 <= a(50) and not w16756;
w16758 <= a(50) and not w16757;
w16759 <= not w16756 and not w16757;
w16760 <= not w16758 and not w16759;
w16761 <= b(18) and w10169;
w16762 <= b(16) and w10539;
w16763 <= b(17) and w10164;
w16764 <= not w16762 and not w16763;
w16765 <= not w16761 and w16764;
w16766 <= w1309 and w10172;
w16767 <= w16765 and not w16766;
w16768 <= a(56) and not w16767;
w16769 <= a(56) and not w16768;
w16770 <= not w16767 and not w16768;
w16771 <= not w16769 and not w16770;
w16772 <= not w16384 and not w16395;
w16773 <= not w16410 and not w16772;
w16774 <= b(12) and w12411;
w16775 <= b(10) and w12790;
w16776 <= b(11) and w12406;
w16777 <= not w16775 and not w16776;
w16778 <= not w16774 and w16777;
w16779 <= w585 and w12414;
w16780 <= w16778 and not w16779;
w16781 <= a(62) and not w16780;
w16782 <= a(62) and not w16781;
w16783 <= not w16780 and not w16781;
w16784 <= not w16782 and not w16783;
w16785 <= b(8) and w13646;
w16786 <= b(9) and not w13231;
w16787 <= not w16785 and not w16786;
w16788 <= a(8) and not w16376;
w16789 <= not a(8) and w16376;
w16790 <= not w16788 and not w16789;
w16791 <= not w16787 and not w16790;
w16792 <= w16787 and w16790;
w16793 <= not w16791 and not w16792;
w16794 <= not w16382 and w16793;
w16795 <= w16382 and not w16793;
w16796 <= not w16794 and not w16795;
w16797 <= w16784 and w16796;
w16798 <= not w16784 and not w16796;
w16799 <= not w16797 and not w16798;
w16800 <= b(15) and w11274;
w16801 <= b(13) and w11639;
w16802 <= b(14) and w11269;
w16803 <= not w16801 and not w16802;
w16804 <= not w16800 and w16803;
w16805 <= w874 and w11277;
w16806 <= w16804 and not w16805;
w16807 <= a(59) and not w16806;
w16808 <= a(59) and not w16807;
w16809 <= not w16806 and not w16807;
w16810 <= not w16808 and not w16809;
w16811 <= not w16799 and not w16810;
w16812 <= w16799 and w16810;
w16813 <= not w16811 and not w16812;
w16814 <= not w16773 and w16813;
w16815 <= w16773 and not w16813;
w16816 <= not w16814 and not w16815;
w16817 <= not w16771 and w16816;
w16818 <= w16816 and not w16817;
w16819 <= not w16771 and not w16817;
w16820 <= not w16818 and not w16819;
w16821 <= not w16414 and not w16427;
w16822 <= w16820 and w16821;
w16823 <= not w16820 and not w16821;
w16824 <= not w16822 and not w16823;
w16825 <= b(21) and w9082;
w16826 <= b(19) and w9475;
w16827 <= b(20) and w9077;
w16828 <= not w16826 and not w16827;
w16829 <= not w16825 and w16828;
w16830 <= w1727 and w9085;
w16831 <= w16829 and not w16830;
w16832 <= a(53) and not w16831;
w16833 <= a(53) and not w16832;
w16834 <= not w16831 and not w16832;
w16835 <= not w16833 and not w16834;
w16836 <= w16824 and not w16835;
w16837 <= w16824 and not w16836;
w16838 <= not w16835 and not w16836;
w16839 <= not w16837 and not w16838;
w16840 <= not w16433 and not w16447;
w16841 <= not w16839 and not w16840;
w16842 <= w16839 and w16840;
w16843 <= not w16841 and not w16842;
w16844 <= not w16760 and w16843;
w16845 <= not w16760 and not w16844;
w16846 <= w16843 and not w16844;
w16847 <= not w16845 and not w16846;
w16848 <= not w16749 and not w16847;
w16849 <= not w16749 and not w16848;
w16850 <= not w16847 and not w16848;
w16851 <= not w16849 and not w16850;
w16852 <= b(27) and w7189;
w16853 <= b(25) and w7530;
w16854 <= b(26) and w7184;
w16855 <= not w16853 and not w16854;
w16856 <= not w16852 and w16855;
w16857 <= w2733 and w7192;
w16858 <= w16856 and not w16857;
w16859 <= a(47) and not w16858;
w16860 <= a(47) and not w16859;
w16861 <= not w16858 and not w16859;
w16862 <= not w16860 and not w16861;
w16863 <= not w16851 and not w16862;
w16864 <= not w16851 and not w16863;
w16865 <= not w16862 and not w16863;
w16866 <= not w16864 and not w16865;
w16867 <= not w16457 and not w16460;
w16868 <= w16866 and w16867;
w16869 <= not w16866 and not w16867;
w16870 <= not w16868 and not w16869;
w16871 <= b(30) and w6338;
w16872 <= b(28) and w6645;
w16873 <= b(29) and w6333;
w16874 <= not w16872 and not w16873;
w16875 <= not w16871 and w16874;
w16876 <= w3320 and w6341;
w16877 <= w16875 and not w16876;
w16878 <= a(44) and not w16877;
w16879 <= a(44) and not w16878;
w16880 <= not w16877 and not w16878;
w16881 <= not w16879 and not w16880;
w16882 <= w16870 and not w16881;
w16883 <= not w16870 and w16881;
w16884 <= not w16748 and not w16883;
w16885 <= not w16882 and w16884;
w16886 <= not w16748 and not w16885;
w16887 <= not w16882 and not w16885;
w16888 <= not w16883 and w16887;
w16889 <= not w16886 and not w16888;
w16890 <= b(33) and w5520;
w16891 <= b(31) and w5802;
w16892 <= b(32) and w5515;
w16893 <= not w16891 and not w16892;
w16894 <= not w16890 and w16893;
w16895 <= w3966 and w5523;
w16896 <= w16894 and not w16895;
w16897 <= a(41) and not w16896;
w16898 <= a(41) and not w16897;
w16899 <= not w16896 and not w16897;
w16900 <= not w16898 and not w16899;
w16901 <= not w16889 and not w16900;
w16902 <= not w16889 and not w16901;
w16903 <= not w16900 and not w16901;
w16904 <= not w16902 and not w16903;
w16905 <= not w16747 and w16904;
w16906 <= w16747 and not w16904;
w16907 <= not w16905 and not w16906;
w16908 <= b(36) and w4778;
w16909 <= b(34) and w5020;
w16910 <= b(35) and w4773;
w16911 <= not w16909 and not w16910;
w16912 <= not w16908 and w16911;
w16913 <= w4665 and w4781;
w16914 <= w16912 and not w16913;
w16915 <= a(38) and not w16914;
w16916 <= a(38) and not w16915;
w16917 <= not w16914 and not w16915;
w16918 <= not w16916 and not w16917;
w16919 <= not w16907 and not w16918;
w16920 <= w16907 and w16918;
w16921 <= not w16919 and not w16920;
w16922 <= w16746 and not w16921;
w16923 <= not w16746 and w16921;
w16924 <= not w16922 and not w16923;
w16925 <= b(39) and w4030;
w16926 <= b(37) and w4275;
w16927 <= b(38) and w4025;
w16928 <= not w16926 and not w16927;
w16929 <= not w16925 and w16928;
w16930 <= w4033 and w5194;
w16931 <= w16929 and not w16930;
w16932 <= a(35) and not w16931;
w16933 <= a(35) and not w16932;
w16934 <= not w16931 and not w16932;
w16935 <= not w16933 and not w16934;
w16936 <= w16924 and not w16935;
w16937 <= w16924 and not w16936;
w16938 <= not w16935 and not w16936;
w16939 <= not w16937 and not w16938;
w16940 <= not w16511 and not w16524;
w16941 <= not w16939 and not w16940;
w16942 <= not w16939 and not w16941;
w16943 <= not w16940 and not w16941;
w16944 <= not w16942 and not w16943;
w16945 <= not w16745 and not w16944;
w16946 <= not w16745 and not w16945;
w16947 <= not w16944 and not w16945;
w16948 <= not w16946 and not w16947;
w16949 <= not w16729 and w16948;
w16950 <= w16729 and not w16948;
w16951 <= not w16949 and not w16950;
w16952 <= w16713 and not w16951;
w16953 <= w16713 and not w16952;
w16954 <= not w16951 and not w16952;
w16955 <= not w16953 and not w16954;
w16956 <= b(51) and w1791;
w16957 <= b(49) and w1941;
w16958 <= b(50) and w1786;
w16959 <= not w16957 and not w16958;
w16960 <= not w16956 and w16959;
w16961 <= w1794 and w8719;
w16962 <= w16960 and not w16961;
w16963 <= a(23) and not w16962;
w16964 <= a(23) and not w16963;
w16965 <= not w16962 and not w16963;
w16966 <= not w16964 and not w16965;
w16967 <= not w16303 and not w16557;
w16968 <= not w16966 and not w16967;
w16969 <= w16966 and w16967;
w16970 <= not w16968 and not w16969;
w16971 <= not w16955 and w16970;
w16972 <= not w16955 and not w16971;
w16973 <= w16970 and not w16971;
w16974 <= not w16972 and not w16973;
w16975 <= not w16698 and not w16974;
w16976 <= not w16698 and not w16975;
w16977 <= not w16974 and not w16975;
w16978 <= not w16976 and not w16977;
w16979 <= w16682 and not w16978;
w16980 <= not w16682 and w16978;
w16981 <= not w16667 and not w16980;
w16982 <= not w16979 and w16981;
w16983 <= not w16667 and not w16982;
w16984 <= not w16980 and not w16982;
w16985 <= not w16979 and w16984;
w16986 <= not w16983 and not w16985;
w16987 <= not w16651 and w16986;
w16988 <= w16651 and not w16986;
w16989 <= not w16987 and not w16988;
w16990 <= not w16635 and not w16989;
w16991 <= not w16635 and not w16990;
w16992 <= not w16989 and not w16990;
w16993 <= not w16991 and not w16992;
w16994 <= not w16634 and not w16993;
w16995 <= w16634 and not w16992;
w16996 <= not w16991 and w16995;
w16997 <= not w16994 and not w16996;
w16998 <= not w16990 and not w16994;
w16999 <= not w16651 and not w16986;
w17000 <= not w16648 and not w16999;
w17001 <= b(61) and w694;
w17002 <= b(59) and w799;
w17003 <= b(60) and w689;
w17004 <= not w17002 and not w17003;
w17005 <= not w17001 and w17004;
w17006 <= w697 and w12712;
w17007 <= w17005 and not w17006;
w17008 <= a(14) and not w17007;
w17009 <= a(14) and not w17008;
w17010 <= not w17007 and not w17008;
w17011 <= not w17009 and not w17010;
w17012 <= not w16681 and not w16979;
w17013 <= not w17011 and not w17012;
w17014 <= not w17011 and not w17013;
w17015 <= not w17012 and not w17013;
w17016 <= not w17014 and not w17015;
w17017 <= b(55) and w1370;
w17018 <= b(53) and w1506;
w17019 <= b(54) and w1365;
w17020 <= not w17018 and not w17019;
w17021 <= not w17017 and w17020;
w17022 <= w1373 and w10427;
w17023 <= w17021 and not w17022;
w17024 <= a(20) and not w17023;
w17025 <= a(20) and not w17024;
w17026 <= not w17023 and not w17024;
w17027 <= not w17025 and not w17026;
w17028 <= not w16968 and not w16971;
w17029 <= w17027 and w17028;
w17030 <= not w17027 and not w17028;
w17031 <= not w17029 and not w17030;
w17032 <= b(52) and w1791;
w17033 <= b(50) and w1941;
w17034 <= b(51) and w1786;
w17035 <= not w17033 and not w17034;
w17036 <= not w17032 and w17035;
w17037 <= w1794 and w9371;
w17038 <= w17036 and not w17037;
w17039 <= a(23) and not w17038;
w17040 <= a(23) and not w17039;
w17041 <= not w17038 and not w17039;
w17042 <= not w17040 and not w17041;
w17043 <= not w16712 and not w16952;
w17044 <= w17042 and w17043;
w17045 <= not w17042 and not w17043;
w17046 <= not w17044 and not w17045;
w17047 <= b(49) and w2282;
w17048 <= b(47) and w2428;
w17049 <= b(48) and w2277;
w17050 <= not w17048 and not w17049;
w17051 <= not w17047 and w17050;
w17052 <= w2285 and w8368;
w17053 <= w17051 and not w17052;
w17054 <= a(26) and not w17053;
w17055 <= a(26) and not w17054;
w17056 <= not w17053 and not w17054;
w17057 <= not w17055 and not w17056;
w17058 <= not w16729 and not w16948;
w17059 <= not w16726 and not w17058;
w17060 <= not w17057 and not w17059;
w17061 <= not w17057 and not w17060;
w17062 <= not w17059 and not w17060;
w17063 <= not w17061 and not w17062;
w17064 <= b(43) and w3381;
w17065 <= b(41) and w3586;
w17066 <= b(42) and w3376;
w17067 <= not w17065 and not w17066;
w17068 <= not w17064 and w17067;
w17069 <= w3384 and w6258;
w17070 <= w17068 and not w17069;
w17071 <= a(32) and not w17070;
w17072 <= a(32) and not w17071;
w17073 <= not w17070 and not w17071;
w17074 <= not w17072 and not w17073;
w17075 <= not w16936 and not w16941;
w17076 <= w17074 and w17075;
w17077 <= not w17074 and not w17075;
w17078 <= not w17076 and not w17077;
w17079 <= b(40) and w4030;
w17080 <= b(38) and w4275;
w17081 <= b(39) and w4025;
w17082 <= not w17080 and not w17081;
w17083 <= not w17079 and w17082;
w17084 <= w4033 and w5698;
w17085 <= w17083 and not w17084;
w17086 <= a(35) and not w17085;
w17087 <= a(35) and not w17086;
w17088 <= not w17085 and not w17086;
w17089 <= not w17087 and not w17088;
w17090 <= not w16919 and not w16923;
w17091 <= b(37) and w4778;
w17092 <= b(35) and w5020;
w17093 <= b(36) and w4773;
w17094 <= not w17092 and not w17093;
w17095 <= not w17091 and w17094;
w17096 <= w4781 and w4924;
w17097 <= w17095 and not w17096;
w17098 <= a(38) and not w17097;
w17099 <= a(38) and not w17098;
w17100 <= not w17097 and not w17098;
w17101 <= not w17099 and not w17100;
w17102 <= not w16747 and not w16904;
w17103 <= not w16901 and not w17102;
w17104 <= b(34) and w5520;
w17105 <= b(32) and w5802;
w17106 <= b(33) and w5515;
w17107 <= not w17105 and not w17106;
w17108 <= not w17104 and w17107;
w17109 <= w4209 and w5523;
w17110 <= w17108 and not w17109;
w17111 <= a(41) and not w17110;
w17112 <= a(41) and not w17111;
w17113 <= not w17110 and not w17111;
w17114 <= not w17112 and not w17113;
w17115 <= b(13) and w12411;
w17116 <= b(11) and w12790;
w17117 <= b(12) and w12406;
w17118 <= not w17116 and not w17117;
w17119 <= not w17115 and w17118;
w17120 <= w751 and w12414;
w17121 <= w17119 and not w17120;
w17122 <= a(62) and not w17121;
w17123 <= a(62) and not w17122;
w17124 <= not w17121 and not w17122;
w17125 <= not w17123 and not w17124;
w17126 <= b(9) and w13646;
w17127 <= b(10) and not w13231;
w17128 <= not w17126 and not w17127;
w17129 <= not a(8) and not w16376;
w17130 <= not w16791 and not w17129;
w17131 <= w17128 and not w17130;
w17132 <= w17128 and not w17131;
w17133 <= not w17130 and not w17131;
w17134 <= not w17132 and not w17133;
w17135 <= not w17125 and not w17134;
w17136 <= not w17125 and not w17135;
w17137 <= not w17134 and not w17135;
w17138 <= not w17136 and not w17137;
w17139 <= not w16784 and w16796;
w17140 <= not w16794 and not w17139;
w17141 <= not w17138 and not w17140;
w17142 <= not w17138 and not w17141;
w17143 <= not w17140 and not w17141;
w17144 <= not w17142 and not w17143;
w17145 <= b(16) and w11274;
w17146 <= b(14) and w11639;
w17147 <= b(15) and w11269;
w17148 <= not w17146 and not w17147;
w17149 <= not w17145 and w17148;
w17150 <= w980 and w11277;
w17151 <= w17149 and not w17150;
w17152 <= a(59) and not w17151;
w17153 <= a(59) and not w17152;
w17154 <= not w17151 and not w17152;
w17155 <= not w17153 and not w17154;
w17156 <= not w17144 and not w17155;
w17157 <= not w17144 and not w17156;
w17158 <= not w17155 and not w17156;
w17159 <= not w17157 and not w17158;
w17160 <= not w16811 and not w16814;
w17161 <= w17159 and w17160;
w17162 <= not w17159 and not w17160;
w17163 <= not w17161 and not w17162;
w17164 <= b(19) and w10169;
w17165 <= b(17) and w10539;
w17166 <= b(18) and w10164;
w17167 <= not w17165 and not w17166;
w17168 <= not w17164 and w17167;
w17169 <= w1451 and w10172;
w17170 <= w17168 and not w17169;
w17171 <= a(56) and not w17170;
w17172 <= a(56) and not w17171;
w17173 <= not w17170 and not w17171;
w17174 <= not w17172 and not w17173;
w17175 <= w17163 and not w17174;
w17176 <= w17163 and not w17175;
w17177 <= not w17174 and not w17175;
w17178 <= not w17176 and not w17177;
w17179 <= not w16817 and not w16823;
w17180 <= w17178 and w17179;
w17181 <= not w17178 and not w17179;
w17182 <= not w17180 and not w17181;
w17183 <= b(22) and w9082;
w17184 <= b(20) and w9475;
w17185 <= b(21) and w9077;
w17186 <= not w17184 and not w17185;
w17187 <= not w17183 and w17186;
w17188 <= w1888 and w9085;
w17189 <= w17187 and not w17188;
w17190 <= a(53) and not w17189;
w17191 <= a(53) and not w17190;
w17192 <= not w17189 and not w17190;
w17193 <= not w17191 and not w17192;
w17194 <= w17182 and not w17193;
w17195 <= w17182 and not w17194;
w17196 <= not w17193 and not w17194;
w17197 <= not w17195 and not w17196;
w17198 <= not w16836 and not w16841;
w17199 <= w17197 and w17198;
w17200 <= not w17197 and not w17198;
w17201 <= not w17199 and not w17200;
w17202 <= b(25) and w8105;
w17203 <= b(23) and w8458;
w17204 <= b(24) and w8100;
w17205 <= not w17203 and not w17204;
w17206 <= not w17202 and w17205;
w17207 <= w2228 and w8108;
w17208 <= w17206 and not w17207;
w17209 <= a(50) and not w17208;
w17210 <= a(50) and not w17209;
w17211 <= not w17208 and not w17209;
w17212 <= not w17210 and not w17211;
w17213 <= w17201 and not w17212;
w17214 <= w17201 and not w17213;
w17215 <= not w17212 and not w17213;
w17216 <= not w17214 and not w17215;
w17217 <= not w16844 and not w16848;
w17218 <= w17216 and w17217;
w17219 <= not w17216 and not w17217;
w17220 <= not w17218 and not w17219;
w17221 <= b(28) and w7189;
w17222 <= b(26) and w7530;
w17223 <= b(27) and w7184;
w17224 <= not w17222 and not w17223;
w17225 <= not w17221 and w17224;
w17226 <= w2932 and w7192;
w17227 <= w17225 and not w17226;
w17228 <= a(47) and not w17227;
w17229 <= a(47) and not w17228;
w17230 <= not w17227 and not w17228;
w17231 <= not w17229 and not w17230;
w17232 <= w17220 and not w17231;
w17233 <= w17220 and not w17232;
w17234 <= not w17231 and not w17232;
w17235 <= not w17233 and not w17234;
w17236 <= not w16863 and not w16869;
w17237 <= w17235 and w17236;
w17238 <= not w17235 and not w17236;
w17239 <= not w17237 and not w17238;
w17240 <= b(31) and w6338;
w17241 <= b(29) and w6645;
w17242 <= b(30) and w6333;
w17243 <= not w17241 and not w17242;
w17244 <= not w17240 and w17243;
w17245 <= w3539 and w6341;
w17246 <= w17244 and not w17245;
w17247 <= a(44) and not w17246;
w17248 <= a(44) and not w17247;
w17249 <= not w17246 and not w17247;
w17250 <= not w17248 and not w17249;
w17251 <= not w17239 and w17250;
w17252 <= w17239 and not w17250;
w17253 <= not w17251 and not w17252;
w17254 <= not w16887 and w17253;
w17255 <= w16887 and not w17253;
w17256 <= not w17254 and not w17255;
w17257 <= not w17114 and w17256;
w17258 <= w17114 and not w17256;
w17259 <= not w17257 and not w17258;
w17260 <= not w17103 and w17259;
w17261 <= not w17103 and not w17260;
w17262 <= w17259 and not w17260;
w17263 <= not w17261 and not w17262;
w17264 <= not w17101 and not w17263;
w17265 <= w17101 and not w17262;
w17266 <= not w17261 and w17265;
w17267 <= not w17264 and not w17266;
w17268 <= not w17090 and w17267;
w17269 <= not w17090 and not w17268;
w17270 <= w17267 and not w17268;
w17271 <= not w17269 and not w17270;
w17272 <= not w17089 and not w17271;
w17273 <= not w17089 and not w17272;
w17274 <= not w17271 and not w17272;
w17275 <= not w17273 and not w17274;
w17276 <= w17078 and not w17275;
w17277 <= w17078 and not w17276;
w17278 <= not w17275 and not w17276;
w17279 <= not w17277 and not w17278;
w17280 <= not w16742 and not w16945;
w17281 <= b(46) and w2793;
w17282 <= b(44) and w2986;
w17283 <= b(45) and w2788;
w17284 <= not w17282 and not w17283;
w17285 <= not w17281 and w17284;
w17286 <= not w2796 and w17285;
w17287 <= not w7420 and w17285;
w17288 <= not w17286 and not w17287;
w17289 <= a(29) and not w17288;
w17290 <= not a(29) and w17288;
w17291 <= not w17289 and not w17290;
w17292 <= not w17280 and not w17291;
w17293 <= not w17280 and not w17292;
w17294 <= not w17291 and not w17292;
w17295 <= not w17293 and not w17294;
w17296 <= not w17279 and not w17295;
w17297 <= not w17279 and not w17296;
w17298 <= not w17295 and not w17296;
w17299 <= not w17297 and not w17298;
w17300 <= not w17063 and not w17299;
w17301 <= not w17063 and not w17300;
w17302 <= not w17299 and not w17300;
w17303 <= not w17301 and not w17302;
w17304 <= w17046 and not w17303;
w17305 <= not w17046 and w17303;
w17306 <= w17031 and not w17305;
w17307 <= not w17304 and w17306;
w17308 <= w17031 and not w17307;
w17309 <= not w17305 and not w17307;
w17310 <= not w17304 and w17309;
w17311 <= not w17308 and not w17310;
w17312 <= not w16695 and not w16975;
w17313 <= b(58) and w1045;
w17314 <= b(56) and w1134;
w17315 <= b(57) and w1040;
w17316 <= not w17314 and not w17315;
w17317 <= not w17313 and w17316;
w17318 <= not w1048 and w17317;
w17319 <= not w11179 and w17317;
w17320 <= not w17318 and not w17319;
w17321 <= a(17) and not w17320;
w17322 <= not a(17) and w17320;
w17323 <= not w17321 and not w17322;
w17324 <= not w17312 and not w17323;
w17325 <= not w17312 and not w17324;
w17326 <= not w17323 and not w17324;
w17327 <= not w17325 and not w17326;
w17328 <= not w17311 and not w17327;
w17329 <= not w17311 and not w17328;
w17330 <= not w17327 and not w17328;
w17331 <= not w17329 and not w17330;
w17332 <= not w17016 and not w17331;
w17333 <= not w17016 and not w17332;
w17334 <= not w17331 and not w17332;
w17335 <= not w17333 and not w17334;
w17336 <= not w16653 and not w16664;
w17337 <= not w16982 and not w17336;
w17338 <= b(62) and w510;
w17339 <= b(63) and w438;
w17340 <= not w17338 and not w17339;
w17341 <= not w446 and w17340;
w17342 <= w13543 and w17340;
w17343 <= not w17341 and not w17342;
w17344 <= a(11) and not w17343;
w17345 <= not a(11) and w17343;
w17346 <= not w17344 and not w17345;
w17347 <= not w17337 and not w17346;
w17348 <= not w17337 and not w17347;
w17349 <= not w17346 and not w17347;
w17350 <= not w17348 and not w17349;
w17351 <= not w17335 and not w17350;
w17352 <= w17335 and not w17349;
w17353 <= not w17348 and w17352;
w17354 <= not w17351 and not w17353;
w17355 <= not w17000 and w17354;
w17356 <= not w17000 and not w17355;
w17357 <= w17354 and not w17355;
w17358 <= not w17356 and not w17357;
w17359 <= not w16998 and not w17358;
w17360 <= w16998 and not w17357;
w17361 <= not w17356 and w17360;
w17362 <= not w17359 and not w17361;
w17363 <= not w17355 and not w17359;
w17364 <= not w17347 and not w17351;
w17365 <= not w17013 and not w17332;
w17366 <= b(63) and w510;
w17367 <= w446 and w13540;
w17368 <= not w17366 and not w17367;
w17369 <= a(11) and not w17368;
w17370 <= a(11) and not w17369;
w17371 <= not w17368 and not w17369;
w17372 <= not w17370 and not w17371;
w17373 <= not w17365 and not w17372;
w17374 <= not w17365 and not w17373;
w17375 <= not w17372 and not w17373;
w17376 <= not w17374 and not w17375;
w17377 <= not w17324 and not w17328;
w17378 <= b(62) and w694;
w17379 <= b(60) and w799;
w17380 <= b(61) and w689;
w17381 <= not w17379 and not w17380;
w17382 <= not w17378 and w17381;
w17383 <= not w697 and w17382;
w17384 <= not w13113 and w17382;
w17385 <= not w17383 and not w17384;
w17386 <= a(14) and not w17385;
w17387 <= not a(14) and w17385;
w17388 <= not w17386 and not w17387;
w17389 <= not w17377 and not w17388;
w17390 <= w17377 and w17388;
w17391 <= not w17389 and not w17390;
w17392 <= b(59) and w1045;
w17393 <= b(57) and w1134;
w17394 <= b(58) and w1040;
w17395 <= not w17393 and not w17394;
w17396 <= not w17392 and w17395;
w17397 <= w1048 and w11922;
w17398 <= w17396 and not w17397;
w17399 <= a(17) and not w17398;
w17400 <= a(17) and not w17399;
w17401 <= not w17398 and not w17399;
w17402 <= not w17400 and not w17401;
w17403 <= not w17030 and not w17307;
w17404 <= w17402 and w17403;
w17405 <= not w17402 and not w17403;
w17406 <= not w17404 and not w17405;
w17407 <= b(56) and w1370;
w17408 <= b(54) and w1506;
w17409 <= b(55) and w1365;
w17410 <= not w17408 and not w17409;
w17411 <= not w17407 and w17410;
w17412 <= w1373 and w10451;
w17413 <= w17411 and not w17412;
w17414 <= a(20) and not w17413;
w17415 <= a(20) and not w17414;
w17416 <= not w17413 and not w17414;
w17417 <= not w17415 and not w17416;
w17418 <= not w17045 and not w17304;
w17419 <= not w17417 and not w17418;
w17420 <= not w17417 and not w17419;
w17421 <= not w17418 and not w17419;
w17422 <= not w17420 and not w17421;
w17423 <= not w17292 and not w17296;
w17424 <= b(50) and w2282;
w17425 <= b(48) and w2428;
w17426 <= b(49) and w2277;
w17427 <= not w17425 and not w17426;
w17428 <= not w17424 and w17427;
w17429 <= not w2285 and w17428;
w17430 <= not w8692 and w17428;
w17431 <= not w17429 and not w17430;
w17432 <= a(26) and not w17431;
w17433 <= not a(26) and w17431;
w17434 <= not w17432 and not w17433;
w17435 <= not w17423 and not w17434;
w17436 <= w17423 and w17434;
w17437 <= not w17435 and not w17436;
w17438 <= b(47) and w2793;
w17439 <= b(45) and w2986;
w17440 <= b(46) and w2788;
w17441 <= not w17439 and not w17440;
w17442 <= not w17438 and w17441;
w17443 <= w2796 and w7446;
w17444 <= w17442 and not w17443;
w17445 <= a(29) and not w17444;
w17446 <= a(29) and not w17445;
w17447 <= not w17444 and not w17445;
w17448 <= not w17446 and not w17447;
w17449 <= not w17077 and not w17276;
w17450 <= w17448 and w17449;
w17451 <= not w17448 and not w17449;
w17452 <= not w17450 and not w17451;
w17453 <= not w17268 and not w17272;
w17454 <= b(44) and w3381;
w17455 <= b(42) and w3586;
w17456 <= b(43) and w3376;
w17457 <= not w17455 and not w17456;
w17458 <= not w17454 and w17457;
w17459 <= not w3384 and w17458;
w17460 <= not w6815 and w17458;
w17461 <= not w17459 and not w17460;
w17462 <= a(32) and not w17461;
w17463 <= not a(32) and w17461;
w17464 <= not w17462 and not w17463;
w17465 <= not w17453 and not w17464;
w17466 <= w17453 and w17464;
w17467 <= not w17465 and not w17466;
w17468 <= b(41) and w4030;
w17469 <= b(39) and w4275;
w17470 <= b(40) and w4025;
w17471 <= not w17469 and not w17470;
w17472 <= not w17468 and w17471;
w17473 <= w4033 and w5962;
w17474 <= w17472 and not w17473;
w17475 <= a(35) and not w17474;
w17476 <= a(35) and not w17475;
w17477 <= not w17474 and not w17475;
w17478 <= not w17476 and not w17477;
w17479 <= not w17260 and not w17264;
w17480 <= b(35) and w5520;
w17481 <= b(33) and w5802;
w17482 <= b(34) and w5515;
w17483 <= not w17481 and not w17482;
w17484 <= not w17480 and w17483;
w17485 <= w4439 and w5523;
w17486 <= w17484 and not w17485;
w17487 <= a(41) and not w17486;
w17488 <= a(41) and not w17487;
w17489 <= not w17486 and not w17487;
w17490 <= not w17488 and not w17489;
w17491 <= not w17200 and not w17213;
w17492 <= b(26) and w8105;
w17493 <= b(24) and w8458;
w17494 <= b(25) and w8100;
w17495 <= not w17493 and not w17494;
w17496 <= not w17492 and w17495;
w17497 <= w2556 and w8108;
w17498 <= w17496 and not w17497;
w17499 <= a(50) and not w17498;
w17500 <= a(50) and not w17499;
w17501 <= not w17498 and not w17499;
w17502 <= not w17500 and not w17501;
w17503 <= not w17181 and not w17194;
w17504 <= b(23) and w9082;
w17505 <= b(21) and w9475;
w17506 <= b(22) and w9077;
w17507 <= not w17505 and not w17506;
w17508 <= not w17504 and w17507;
w17509 <= w2043 and w9085;
w17510 <= w17508 and not w17509;
w17511 <= a(53) and not w17510;
w17512 <= a(53) and not w17511;
w17513 <= not w17510 and not w17511;
w17514 <= not w17512 and not w17513;
w17515 <= not w17162 and not w17175;
w17516 <= not w17131 and not w17135;
w17517 <= b(10) and w13646;
w17518 <= b(11) and not w13231;
w17519 <= not w17517 and not w17518;
w17520 <= w17128 and not w17519;
w17521 <= w17128 and not w17520;
w17522 <= not w17519 and not w17520;
w17523 <= not w17521 and not w17522;
w17524 <= not w17516 and not w17523;
w17525 <= not w17516 and not w17524;
w17526 <= not w17523 and not w17524;
w17527 <= not w17525 and not w17526;
w17528 <= b(14) and w12411;
w17529 <= b(12) and w12790;
w17530 <= b(13) and w12406;
w17531 <= not w17529 and not w17530;
w17532 <= not w17528 and w17531;
w17533 <= w777 and w12414;
w17534 <= w17532 and not w17533;
w17535 <= a(62) and not w17534;
w17536 <= a(62) and not w17535;
w17537 <= not w17534 and not w17535;
w17538 <= not w17536 and not w17537;
w17539 <= not w17527 and not w17538;
w17540 <= not w17527 and not w17539;
w17541 <= not w17538 and not w17539;
w17542 <= not w17540 and not w17541;
w17543 <= b(17) and w11274;
w17544 <= b(15) and w11639;
w17545 <= b(16) and w11269;
w17546 <= not w17544 and not w17545;
w17547 <= not w17543 and w17546;
w17548 <= w1099 and w11277;
w17549 <= w17547 and not w17548;
w17550 <= a(59) and not w17549;
w17551 <= a(59) and not w17550;
w17552 <= not w17549 and not w17550;
w17553 <= not w17551 and not w17552;
w17554 <= not w17542 and not w17553;
w17555 <= not w17542 and not w17554;
w17556 <= not w17553 and not w17554;
w17557 <= not w17555 and not w17556;
w17558 <= not w17141 and not w17156;
w17559 <= w17557 and w17558;
w17560 <= not w17557 and not w17558;
w17561 <= not w17559 and not w17560;
w17562 <= b(20) and w10169;
w17563 <= b(18) and w10539;
w17564 <= b(19) and w10164;
w17565 <= not w17563 and not w17564;
w17566 <= not w17562 and w17565;
w17567 <= w1589 and w10172;
w17568 <= w17566 and not w17567;
w17569 <= a(56) and not w17568;
w17570 <= a(56) and not w17569;
w17571 <= not w17568 and not w17569;
w17572 <= not w17570 and not w17571;
w17573 <= not w17561 and w17572;
w17574 <= w17561 and not w17572;
w17575 <= not w17573 and not w17574;
w17576 <= not w17515 and w17575;
w17577 <= not w17515 and not w17576;
w17578 <= w17575 and not w17576;
w17579 <= not w17577 and not w17578;
w17580 <= not w17514 and not w17579;
w17581 <= w17514 and not w17578;
w17582 <= not w17577 and w17581;
w17583 <= not w17580 and not w17582;
w17584 <= not w17503 and w17583;
w17585 <= w17503 and not w17583;
w17586 <= not w17584 and not w17585;
w17587 <= not w17502 and w17586;
w17588 <= w17502 and not w17586;
w17589 <= not w17587 and not w17588;
w17590 <= not w17491 and w17589;
w17591 <= w17491 and not w17589;
w17592 <= not w17590 and not w17591;
w17593 <= b(29) and w7189;
w17594 <= b(27) and w7530;
w17595 <= b(28) and w7184;
w17596 <= not w17594 and not w17595;
w17597 <= not w17593 and w17596;
w17598 <= w3126 and w7192;
w17599 <= w17597 and not w17598;
w17600 <= a(47) and not w17599;
w17601 <= a(47) and not w17600;
w17602 <= not w17599 and not w17600;
w17603 <= not w17601 and not w17602;
w17604 <= w17592 and not w17603;
w17605 <= w17592 and not w17604;
w17606 <= not w17603 and not w17604;
w17607 <= not w17605 and not w17606;
w17608 <= not w17219 and not w17232;
w17609 <= w17607 and w17608;
w17610 <= not w17607 and not w17608;
w17611 <= not w17609 and not w17610;
w17612 <= b(32) and w6338;
w17613 <= b(30) and w6645;
w17614 <= b(31) and w6333;
w17615 <= not w17613 and not w17614;
w17616 <= not w17612 and w17615;
w17617 <= w3756 and w6341;
w17618 <= w17616 and not w17617;
w17619 <= a(44) and not w17618;
w17620 <= a(44) and not w17619;
w17621 <= not w17618 and not w17619;
w17622 <= not w17620 and not w17621;
w17623 <= not w17611 and w17622;
w17624 <= w17611 and not w17622;
w17625 <= not w17623 and not w17624;
w17626 <= not w17238 and not w17252;
w17627 <= w17625 and not w17626;
w17628 <= not w17625 and w17626;
w17629 <= not w17627 and not w17628;
w17630 <= not w17490 and w17629;
w17631 <= w17629 and not w17630;
w17632 <= not w17490 and not w17630;
w17633 <= not w17631 and not w17632;
w17634 <= not w17254 and not w17257;
w17635 <= w17633 and w17634;
w17636 <= not w17633 and not w17634;
w17637 <= not w17635 and not w17636;
w17638 <= b(38) and w4778;
w17639 <= b(36) and w5020;
w17640 <= b(37) and w4773;
w17641 <= not w17639 and not w17640;
w17642 <= not w17638 and w17641;
w17643 <= w4781 and w4948;
w17644 <= w17642 and not w17643;
w17645 <= a(38) and not w17644;
w17646 <= a(38) and not w17645;
w17647 <= not w17644 and not w17645;
w17648 <= not w17646 and not w17647;
w17649 <= not w17637 and w17648;
w17650 <= w17637 and not w17648;
w17651 <= not w17649 and not w17650;
w17652 <= not w17479 and w17651;
w17653 <= w17479 and not w17651;
w17654 <= not w17652 and not w17653;
w17655 <= not w17478 and w17654;
w17656 <= not w17478 and not w17655;
w17657 <= w17654 and not w17655;
w17658 <= not w17656 and not w17657;
w17659 <= w17467 and not w17658;
w17660 <= w17467 and not w17659;
w17661 <= not w17658 and not w17659;
w17662 <= not w17660 and not w17661;
w17663 <= w17452 and not w17662;
w17664 <= not w17452 and w17662;
w17665 <= w17437 and not w17664;
w17666 <= not w17663 and w17665;
w17667 <= w17437 and not w17666;
w17668 <= not w17664 and not w17666;
w17669 <= not w17663 and w17668;
w17670 <= not w17667 and not w17669;
w17671 <= not w17060 and not w17300;
w17672 <= b(53) and w1791;
w17673 <= b(51) and w1941;
w17674 <= b(52) and w1786;
w17675 <= not w17673 and not w17674;
w17676 <= not w17672 and w17675;
w17677 <= not w1794 and w17676;
w17678 <= not w9715 and w17676;
w17679 <= not w17677 and not w17678;
w17680 <= a(23) and not w17679;
w17681 <= not a(23) and w17679;
w17682 <= not w17680 and not w17681;
w17683 <= not w17671 and not w17682;
w17684 <= not w17671 and not w17683;
w17685 <= not w17682 and not w17683;
w17686 <= not w17684 and not w17685;
w17687 <= not w17670 and not w17686;
w17688 <= not w17670 and not w17687;
w17689 <= not w17686 and not w17687;
w17690 <= not w17688 and not w17689;
w17691 <= not w17422 and not w17690;
w17692 <= not w17422 and not w17691;
w17693 <= not w17690 and not w17691;
w17694 <= not w17692 and not w17693;
w17695 <= w17406 and not w17694;
w17696 <= not w17406 and w17694;
w17697 <= w17391 and not w17696;
w17698 <= not w17695 and w17697;
w17699 <= w17391 and not w17698;
w17700 <= not w17696 and not w17698;
w17701 <= not w17695 and w17700;
w17702 <= not w17699 and not w17701;
w17703 <= not w17376 and w17702;
w17704 <= w17376 and not w17702;
w17705 <= not w17703 and not w17704;
w17706 <= not w17364 and not w17705;
w17707 <= not w17364 and not w17706;
w17708 <= not w17705 and not w17706;
w17709 <= not w17707 and not w17708;
w17710 <= not w17363 and not w17709;
w17711 <= w17363 and not w17708;
w17712 <= not w17707 and w17711;
w17713 <= not w17710 and not w17712;
w17714 <= not w17706 and not w17710;
w17715 <= not w17376 and not w17702;
w17716 <= not w17373 and not w17715;
w17717 <= not w17389 and not w17698;
w17718 <= b(63) and w694;
w17719 <= b(61) and w799;
w17720 <= b(62) and w689;
w17721 <= not w17719 and not w17720;
w17722 <= not w17718 and w17721;
w17723 <= w697 and w13514;
w17724 <= w17722 and not w17723;
w17725 <= a(14) and not w17724;
w17726 <= a(14) and not w17725;
w17727 <= not w17724 and not w17725;
w17728 <= not w17726 and not w17727;
w17729 <= not w17717 and not w17728;
w17730 <= not w17717 and not w17729;
w17731 <= not w17728 and not w17729;
w17732 <= not w17730 and not w17731;
w17733 <= not w17405 and not w17695;
w17734 <= b(60) and w1045;
w17735 <= b(58) and w1134;
w17736 <= b(59) and w1040;
w17737 <= not w17735 and not w17736;
w17738 <= not w17734 and w17737;
w17739 <= w1048 and w11954;
w17740 <= w17738 and not w17739;
w17741 <= a(17) and not w17740;
w17742 <= a(17) and not w17741;
w17743 <= not w17740 and not w17741;
w17744 <= not w17742 and not w17743;
w17745 <= not w17733 and w17744;
w17746 <= w17733 and not w17744;
w17747 <= not w17745 and not w17746;
w17748 <= b(57) and w1370;
w17749 <= b(55) and w1506;
w17750 <= b(56) and w1365;
w17751 <= not w17749 and not w17750;
w17752 <= not w17748 and w17751;
w17753 <= w1373 and w11153;
w17754 <= w17752 and not w17753;
w17755 <= a(20) and not w17754;
w17756 <= a(20) and not w17755;
w17757 <= not w17754 and not w17755;
w17758 <= not w17756 and not w17757;
w17759 <= not w17419 and not w17691;
w17760 <= w17758 and w17759;
w17761 <= not w17758 and not w17759;
w17762 <= not w17760 and not w17761;
w17763 <= not w17683 and not w17687;
w17764 <= b(54) and w1791;
w17765 <= b(52) and w1941;
w17766 <= b(53) and w1786;
w17767 <= not w17765 and not w17766;
w17768 <= not w17764 and w17767;
w17769 <= w1794 and w9741;
w17770 <= w17768 and not w17769;
w17771 <= a(23) and not w17770;
w17772 <= a(23) and not w17771;
w17773 <= not w17770 and not w17771;
w17774 <= not w17772 and not w17773;
w17775 <= not w17763 and not w17774;
w17776 <= not w17763 and not w17775;
w17777 <= not w17774 and not w17775;
w17778 <= not w17776 and not w17777;
w17779 <= b(51) and w2282;
w17780 <= b(49) and w2428;
w17781 <= b(50) and w2277;
w17782 <= not w17780 and not w17781;
w17783 <= not w17779 and w17782;
w17784 <= w2285 and w8719;
w17785 <= w17783 and not w17784;
w17786 <= a(26) and not w17785;
w17787 <= a(26) and not w17786;
w17788 <= not w17785 and not w17786;
w17789 <= not w17787 and not w17788;
w17790 <= not w17435 and not w17666;
w17791 <= w17789 and w17790;
w17792 <= not w17789 and not w17790;
w17793 <= not w17791 and not w17792;
w17794 <= not w17451 and not w17663;
w17795 <= b(48) and w2793;
w17796 <= b(46) and w2986;
w17797 <= b(47) and w2788;
w17798 <= not w17796 and not w17797;
w17799 <= not w17795 and w17798;
w17800 <= w2796 and w7752;
w17801 <= w17799 and not w17800;
w17802 <= a(29) and not w17801;
w17803 <= a(29) and not w17802;
w17804 <= not w17801 and not w17802;
w17805 <= not w17803 and not w17804;
w17806 <= not w17794 and w17805;
w17807 <= w17794 and not w17805;
w17808 <= not w17806 and not w17807;
w17809 <= not w17652 and not w17655;
w17810 <= not w17636 and not w17650;
w17811 <= not w17627 and not w17630;
w17812 <= not w17610 and not w17624;
w17813 <= not w17590 and not w17604;
w17814 <= not w17576 and not w17580;
w17815 <= b(24) and w9082;
w17816 <= b(22) and w9475;
w17817 <= b(23) and w9077;
w17818 <= not w17816 and not w17817;
w17819 <= not w17815 and w17818;
w17820 <= w2201 and w9085;
w17821 <= w17819 and not w17820;
w17822 <= a(53) and not w17821;
w17823 <= a(53) and not w17822;
w17824 <= not w17821 and not w17822;
w17825 <= not w17823 and not w17824;
w17826 <= not w17520 and not w17524;
w17827 <= b(15) and w12411;
w17828 <= b(13) and w12790;
w17829 <= b(14) and w12406;
w17830 <= not w17828 and not w17829;
w17831 <= not w17827 and w17830;
w17832 <= w874 and w12414;
w17833 <= w17831 and not w17832;
w17834 <= a(62) and not w17833;
w17835 <= a(62) and not w17834;
w17836 <= not w17833 and not w17834;
w17837 <= not w17835 and not w17836;
w17838 <= b(11) and w13646;
w17839 <= b(12) and not w13231;
w17840 <= not w17838 and not w17839;
w17841 <= a(11) and not w17128;
w17842 <= not a(11) and w17128;
w17843 <= not w17841 and not w17842;
w17844 <= not w17840 and not w17843;
w17845 <= w17840 and w17843;
w17846 <= not w17844 and not w17845;
w17847 <= not w17837 and w17846;
w17848 <= not w17837 and not w17847;
w17849 <= w17846 and not w17847;
w17850 <= not w17848 and not w17849;
w17851 <= not w17826 and not w17850;
w17852 <= not w17826 and not w17851;
w17853 <= not w17850 and not w17851;
w17854 <= not w17852 and not w17853;
w17855 <= b(18) and w11274;
w17856 <= b(16) and w11639;
w17857 <= b(17) and w11269;
w17858 <= not w17856 and not w17857;
w17859 <= not w17855 and w17858;
w17860 <= w1309 and w11277;
w17861 <= w17859 and not w17860;
w17862 <= a(59) and not w17861;
w17863 <= a(59) and not w17862;
w17864 <= not w17861 and not w17862;
w17865 <= not w17863 and not w17864;
w17866 <= not w17854 and not w17865;
w17867 <= not w17854 and not w17866;
w17868 <= not w17865 and not w17866;
w17869 <= not w17867 and not w17868;
w17870 <= not w17539 and not w17554;
w17871 <= w17869 and w17870;
w17872 <= not w17869 and not w17870;
w17873 <= not w17871 and not w17872;
w17874 <= b(21) and w10169;
w17875 <= b(19) and w10539;
w17876 <= b(20) and w10164;
w17877 <= not w17875 and not w17876;
w17878 <= not w17874 and w17877;
w17879 <= w1727 and w10172;
w17880 <= w17878 and not w17879;
w17881 <= a(56) and not w17880;
w17882 <= a(56) and not w17881;
w17883 <= not w17880 and not w17881;
w17884 <= not w17882 and not w17883;
w17885 <= w17873 and not w17884;
w17886 <= w17873 and not w17885;
w17887 <= not w17884 and not w17885;
w17888 <= not w17886 and not w17887;
w17889 <= not w17560 and not w17574;
w17890 <= not w17888 and not w17889;
w17891 <= w17888 and w17889;
w17892 <= not w17890 and not w17891;
w17893 <= not w17825 and w17892;
w17894 <= not w17825 and not w17893;
w17895 <= w17892 and not w17893;
w17896 <= not w17894 and not w17895;
w17897 <= not w17814 and not w17896;
w17898 <= not w17814 and not w17897;
w17899 <= not w17896 and not w17897;
w17900 <= not w17898 and not w17899;
w17901 <= b(27) and w8105;
w17902 <= b(25) and w8458;
w17903 <= b(26) and w8100;
w17904 <= not w17902 and not w17903;
w17905 <= not w17901 and w17904;
w17906 <= w2733 and w8108;
w17907 <= w17905 and not w17906;
w17908 <= a(50) and not w17907;
w17909 <= a(50) and not w17908;
w17910 <= not w17907 and not w17908;
w17911 <= not w17909 and not w17910;
w17912 <= not w17900 and not w17911;
w17913 <= not w17900 and not w17912;
w17914 <= not w17911 and not w17912;
w17915 <= not w17913 and not w17914;
w17916 <= not w17584 and not w17587;
w17917 <= w17915 and w17916;
w17918 <= not w17915 and not w17916;
w17919 <= not w17917 and not w17918;
w17920 <= b(30) and w7189;
w17921 <= b(28) and w7530;
w17922 <= b(29) and w7184;
w17923 <= not w17921 and not w17922;
w17924 <= not w17920 and w17923;
w17925 <= w3320 and w7192;
w17926 <= w17924 and not w17925;
w17927 <= a(47) and not w17926;
w17928 <= a(47) and not w17927;
w17929 <= not w17926 and not w17927;
w17930 <= not w17928 and not w17929;
w17931 <= w17919 and not w17930;
w17932 <= not w17919 and w17930;
w17933 <= not w17813 and not w17932;
w17934 <= not w17931 and w17933;
w17935 <= not w17813 and not w17934;
w17936 <= not w17931 and not w17934;
w17937 <= not w17932 and w17936;
w17938 <= not w17935 and not w17937;
w17939 <= b(33) and w6338;
w17940 <= b(31) and w6645;
w17941 <= b(32) and w6333;
w17942 <= not w17940 and not w17941;
w17943 <= not w17939 and w17942;
w17944 <= w3966 and w6341;
w17945 <= w17943 and not w17944;
w17946 <= a(44) and not w17945;
w17947 <= a(44) and not w17946;
w17948 <= not w17945 and not w17946;
w17949 <= not w17947 and not w17948;
w17950 <= not w17938 and not w17949;
w17951 <= not w17938 and not w17950;
w17952 <= not w17949 and not w17950;
w17953 <= not w17951 and not w17952;
w17954 <= not w17812 and w17953;
w17955 <= w17812 and not w17953;
w17956 <= not w17954 and not w17955;
w17957 <= b(36) and w5520;
w17958 <= b(34) and w5802;
w17959 <= b(35) and w5515;
w17960 <= not w17958 and not w17959;
w17961 <= not w17957 and w17960;
w17962 <= w4665 and w5523;
w17963 <= w17961 and not w17962;
w17964 <= a(41) and not w17963;
w17965 <= a(41) and not w17964;
w17966 <= not w17963 and not w17964;
w17967 <= not w17965 and not w17966;
w17968 <= not w17956 and not w17967;
w17969 <= w17956 and w17967;
w17970 <= not w17968 and not w17969;
w17971 <= w17811 and not w17970;
w17972 <= not w17811 and w17970;
w17973 <= not w17971 and not w17972;
w17974 <= b(39) and w4778;
w17975 <= b(37) and w5020;
w17976 <= b(38) and w4773;
w17977 <= not w17975 and not w17976;
w17978 <= not w17974 and w17977;
w17979 <= w4781 and w5194;
w17980 <= w17978 and not w17979;
w17981 <= a(38) and not w17980;
w17982 <= a(38) and not w17981;
w17983 <= not w17980 and not w17981;
w17984 <= not w17982 and not w17983;
w17985 <= w17973 and not w17984;
w17986 <= w17973 and not w17985;
w17987 <= not w17984 and not w17985;
w17988 <= not w17986 and not w17987;
w17989 <= not w17810 and w17988;
w17990 <= w17810 and not w17988;
w17991 <= not w17989 and not w17990;
w17992 <= b(42) and w4030;
w17993 <= b(40) and w4275;
w17994 <= b(41) and w4025;
w17995 <= not w17993 and not w17994;
w17996 <= not w17992 and w17995;
w17997 <= w4033 and w6232;
w17998 <= w17996 and not w17997;
w17999 <= a(35) and not w17998;
w18000 <= a(35) and not w17999;
w18001 <= not w17998 and not w17999;
w18002 <= not w18000 and not w18001;
w18003 <= not w17991 and not w18002;
w18004 <= w17991 and w18002;
w18005 <= not w18003 and not w18004;
w18006 <= w17809 and not w18005;
w18007 <= not w17809 and w18005;
w18008 <= not w18006 and not w18007;
w18009 <= not w17465 and not w17659;
w18010 <= b(45) and w3381;
w18011 <= b(43) and w3586;
w18012 <= b(44) and w3376;
w18013 <= not w18011 and not w18012;
w18014 <= not w18010 and w18013;
w18015 <= w3384 and w7104;
w18016 <= w18014 and not w18015;
w18017 <= a(32) and not w18016;
w18018 <= a(32) and not w18017;
w18019 <= not w18016 and not w18017;
w18020 <= not w18018 and not w18019;
w18021 <= not w18009 and not w18020;
w18022 <= not w18009 and not w18021;
w18023 <= not w18020 and not w18021;
w18024 <= not w18022 and not w18023;
w18025 <= w18008 and not w18024;
w18026 <= not w18008 and w18024;
w18027 <= not w17808 and not w18026;
w18028 <= not w18025 and w18027;
w18029 <= not w17808 and not w18028;
w18030 <= not w18026 and not w18028;
w18031 <= not w18025 and w18030;
w18032 <= not w18029 and not w18031;
w18033 <= w17793 and not w18032;
w18034 <= not w17793 and w18032;
w18035 <= not w17778 and not w18034;
w18036 <= not w18033 and w18035;
w18037 <= not w17778 and not w18036;
w18038 <= not w18034 and not w18036;
w18039 <= not w18033 and w18038;
w18040 <= not w18037 and not w18039;
w18041 <= w17762 and not w18040;
w18042 <= not w17762 and w18040;
w18043 <= not w17747 and not w18042;
w18044 <= not w18041 and w18043;
w18045 <= not w17747 and not w18044;
w18046 <= not w18042 and not w18044;
w18047 <= not w18041 and w18046;
w18048 <= not w18045 and not w18047;
w18049 <= not w17732 and w18048;
w18050 <= w17732 and not w18048;
w18051 <= not w18049 and not w18050;
w18052 <= not w17716 and not w18051;
w18053 <= not w17716 and not w18052;
w18054 <= not w18051 and not w18052;
w18055 <= not w18053 and not w18054;
w18056 <= not w17714 and not w18055;
w18057 <= w17714 and not w18054;
w18058 <= not w18053 and w18057;
w18059 <= not w18056 and not w18058;
w18060 <= not w18052 and not w18056;
w18061 <= not w17732 and not w18048;
w18062 <= not w17729 and not w18061;
w18063 <= b(61) and w1045;
w18064 <= b(59) and w1134;
w18065 <= b(60) and w1040;
w18066 <= not w18064 and not w18065;
w18067 <= not w18063 and w18066;
w18068 <= w1048 and w12712;
w18069 <= w18067 and not w18068;
w18070 <= a(17) and not w18069;
w18071 <= a(17) and not w18070;
w18072 <= not w18069 and not w18070;
w18073 <= not w18071 and not w18072;
w18074 <= not w17761 and not w18041;
w18075 <= not w18073 and not w18074;
w18076 <= not w18073 and not w18075;
w18077 <= not w18074 and not w18075;
w18078 <= not w18076 and not w18077;
w18079 <= b(55) and w1791;
w18080 <= b(53) and w1941;
w18081 <= b(54) and w1786;
w18082 <= not w18080 and not w18081;
w18083 <= not w18079 and w18082;
w18084 <= w1794 and w10427;
w18085 <= w18083 and not w18084;
w18086 <= a(23) and not w18085;
w18087 <= a(23) and not w18086;
w18088 <= not w18085 and not w18086;
w18089 <= not w18087 and not w18088;
w18090 <= not w17792 and not w18033;
w18091 <= not w18089 and not w18090;
w18092 <= not w18089 and not w18091;
w18093 <= not w18090 and not w18091;
w18094 <= not w18092 and not w18093;
w18095 <= b(49) and w2793;
w18096 <= b(47) and w2986;
w18097 <= b(48) and w2788;
w18098 <= not w18096 and not w18097;
w18099 <= not w18095 and w18098;
w18100 <= w2796 and w8368;
w18101 <= w18099 and not w18100;
w18102 <= a(29) and not w18101;
w18103 <= a(29) and not w18102;
w18104 <= not w18101 and not w18102;
w18105 <= not w18103 and not w18104;
w18106 <= not w18021 and not w18025;
w18107 <= not w18105 and not w18106;
w18108 <= not w18105 and not w18107;
w18109 <= not w18106 and not w18107;
w18110 <= not w18108 and not w18109;
w18111 <= b(43) and w4030;
w18112 <= b(41) and w4275;
w18113 <= b(42) and w4025;
w18114 <= not w18112 and not w18113;
w18115 <= not w18111 and w18114;
w18116 <= w4033 and w6258;
w18117 <= w18115 and not w18116;
w18118 <= a(35) and not w18117;
w18119 <= a(35) and not w18118;
w18120 <= not w18117 and not w18118;
w18121 <= not w18119 and not w18120;
w18122 <= not w17810 and not w17988;
w18123 <= not w17985 and not w18122;
w18124 <= b(40) and w4778;
w18125 <= b(38) and w5020;
w18126 <= b(39) and w4773;
w18127 <= not w18125 and not w18126;
w18128 <= not w18124 and w18127;
w18129 <= w4781 and w5698;
w18130 <= w18128 and not w18129;
w18131 <= a(38) and not w18130;
w18132 <= a(38) and not w18131;
w18133 <= not w18130 and not w18131;
w18134 <= not w18132 and not w18133;
w18135 <= not w17968 and not w17972;
w18136 <= b(37) and w5520;
w18137 <= b(35) and w5802;
w18138 <= b(36) and w5515;
w18139 <= not w18137 and not w18138;
w18140 <= not w18136 and w18139;
w18141 <= w4924 and w5523;
w18142 <= w18140 and not w18141;
w18143 <= a(41) and not w18142;
w18144 <= a(41) and not w18143;
w18145 <= not w18142 and not w18143;
w18146 <= not w18144 and not w18145;
w18147 <= not w17812 and not w17953;
w18148 <= not w17950 and not w18147;
w18149 <= b(34) and w6338;
w18150 <= b(32) and w6645;
w18151 <= b(33) and w6333;
w18152 <= not w18150 and not w18151;
w18153 <= not w18149 and w18152;
w18154 <= w4209 and w6341;
w18155 <= w18153 and not w18154;
w18156 <= a(44) and not w18155;
w18157 <= a(44) and not w18156;
w18158 <= not w18155 and not w18156;
w18159 <= not w18157 and not w18158;
w18160 <= b(31) and w7189;
w18161 <= b(29) and w7530;
w18162 <= b(30) and w7184;
w18163 <= not w18161 and not w18162;
w18164 <= not w18160 and w18163;
w18165 <= w3539 and w7192;
w18166 <= w18164 and not w18165;
w18167 <= a(47) and not w18166;
w18168 <= a(47) and not w18167;
w18169 <= not w18166 and not w18167;
w18170 <= not w18168 and not w18169;
w18171 <= not w17912 and not w17918;
w18172 <= b(12) and w13646;
w18173 <= b(13) and not w13231;
w18174 <= not w18172 and not w18173;
w18175 <= not a(11) and not w17128;
w18176 <= not w17844 and not w18175;
w18177 <= w18174 and not w18176;
w18178 <= w18174 and not w18177;
w18179 <= not w18176 and not w18177;
w18180 <= not w18178 and not w18179;
w18181 <= b(16) and w12411;
w18182 <= b(14) and w12790;
w18183 <= b(15) and w12406;
w18184 <= not w18182 and not w18183;
w18185 <= not w18181 and w18184;
w18186 <= w980 and w12414;
w18187 <= w18185 and not w18186;
w18188 <= a(62) and not w18187;
w18189 <= a(62) and not w18188;
w18190 <= not w18187 and not w18188;
w18191 <= not w18189 and not w18190;
w18192 <= not w18180 and w18191;
w18193 <= w18180 and not w18191;
w18194 <= not w18192 and not w18193;
w18195 <= not w17847 and not w17851;
w18196 <= w18194 and w18195;
w18197 <= not w18194 and not w18195;
w18198 <= not w18196 and not w18197;
w18199 <= b(19) and w11274;
w18200 <= b(17) and w11639;
w18201 <= b(18) and w11269;
w18202 <= not w18200 and not w18201;
w18203 <= not w18199 and w18202;
w18204 <= w1451 and w11277;
w18205 <= w18203 and not w18204;
w18206 <= a(59) and not w18205;
w18207 <= a(59) and not w18206;
w18208 <= not w18205 and not w18206;
w18209 <= not w18207 and not w18208;
w18210 <= w18198 and not w18209;
w18211 <= w18198 and not w18210;
w18212 <= not w18209 and not w18210;
w18213 <= not w18211 and not w18212;
w18214 <= not w17866 and not w17872;
w18215 <= w18213 and w18214;
w18216 <= not w18213 and not w18214;
w18217 <= not w18215 and not w18216;
w18218 <= b(22) and w10169;
w18219 <= b(20) and w10539;
w18220 <= b(21) and w10164;
w18221 <= not w18219 and not w18220;
w18222 <= not w18218 and w18221;
w18223 <= w1888 and w10172;
w18224 <= w18222 and not w18223;
w18225 <= a(56) and not w18224;
w18226 <= a(56) and not w18225;
w18227 <= not w18224 and not w18225;
w18228 <= not w18226 and not w18227;
w18229 <= w18217 and not w18228;
w18230 <= w18217 and not w18229;
w18231 <= not w18228 and not w18229;
w18232 <= not w18230 and not w18231;
w18233 <= not w17885 and not w17890;
w18234 <= w18232 and w18233;
w18235 <= not w18232 and not w18233;
w18236 <= not w18234 and not w18235;
w18237 <= b(25) and w9082;
w18238 <= b(23) and w9475;
w18239 <= b(24) and w9077;
w18240 <= not w18238 and not w18239;
w18241 <= not w18237 and w18240;
w18242 <= w2228 and w9085;
w18243 <= w18241 and not w18242;
w18244 <= a(53) and not w18243;
w18245 <= a(53) and not w18244;
w18246 <= not w18243 and not w18244;
w18247 <= not w18245 and not w18246;
w18248 <= w18236 and not w18247;
w18249 <= w18236 and not w18248;
w18250 <= not w18247 and not w18248;
w18251 <= not w18249 and not w18250;
w18252 <= not w17893 and not w17897;
w18253 <= w18251 and w18252;
w18254 <= not w18251 and not w18252;
w18255 <= not w18253 and not w18254;
w18256 <= b(28) and w8105;
w18257 <= b(26) and w8458;
w18258 <= b(27) and w8100;
w18259 <= not w18257 and not w18258;
w18260 <= not w18256 and w18259;
w18261 <= w2932 and w8108;
w18262 <= w18260 and not w18261;
w18263 <= a(50) and not w18262;
w18264 <= a(50) and not w18263;
w18265 <= not w18262 and not w18263;
w18266 <= not w18264 and not w18265;
w18267 <= not w18255 and w18266;
w18268 <= w18255 and not w18266;
w18269 <= not w18267 and not w18268;
w18270 <= not w18171 and w18269;
w18271 <= not w18171 and not w18270;
w18272 <= w18269 and not w18270;
w18273 <= not w18271 and not w18272;
w18274 <= not w18170 and not w18273;
w18275 <= w18170 and not w18272;
w18276 <= not w18271 and w18275;
w18277 <= not w18274 and not w18276;
w18278 <= not w17936 and w18277;
w18279 <= w17936 and not w18277;
w18280 <= not w18278 and not w18279;
w18281 <= not w18159 and w18280;
w18282 <= w18159 and not w18280;
w18283 <= not w18281 and not w18282;
w18284 <= not w18148 and w18283;
w18285 <= not w18148 and not w18284;
w18286 <= w18283 and not w18284;
w18287 <= not w18285 and not w18286;
w18288 <= not w18146 and not w18287;
w18289 <= w18146 and not w18286;
w18290 <= not w18285 and w18289;
w18291 <= not w18288 and not w18290;
w18292 <= not w18135 and w18291;
w18293 <= not w18135 and not w18292;
w18294 <= w18291 and not w18292;
w18295 <= not w18293 and not w18294;
w18296 <= not w18134 and not w18295;
w18297 <= w18134 and not w18294;
w18298 <= not w18293 and w18297;
w18299 <= not w18296 and not w18298;
w18300 <= not w18123 and w18299;
w18301 <= w18123 and not w18299;
w18302 <= not w18300 and not w18301;
w18303 <= not w18121 and w18302;
w18304 <= w18302 and not w18303;
w18305 <= not w18121 and not w18303;
w18306 <= not w18304 and not w18305;
w18307 <= not w18003 and not w18007;
w18308 <= b(46) and w3381;
w18309 <= b(44) and w3586;
w18310 <= b(45) and w3376;
w18311 <= not w18309 and not w18310;
w18312 <= not w18308 and w18311;
w18313 <= not w3384 and w18312;
w18314 <= not w7420 and w18312;
w18315 <= not w18313 and not w18314;
w18316 <= a(32) and not w18315;
w18317 <= not a(32) and w18315;
w18318 <= not w18316 and not w18317;
w18319 <= not w18307 and not w18318;
w18320 <= not w18307 and not w18319;
w18321 <= not w18318 and not w18319;
w18322 <= not w18320 and not w18321;
w18323 <= not w18306 and not w18322;
w18324 <= not w18306 and not w18323;
w18325 <= not w18322 and not w18323;
w18326 <= not w18324 and not w18325;
w18327 <= not w18110 and not w18326;
w18328 <= not w18110 and not w18327;
w18329 <= not w18326 and not w18327;
w18330 <= not w18328 and not w18329;
w18331 <= not w17794 and not w17805;
w18332 <= not w18028 and not w18331;
w18333 <= b(52) and w2282;
w18334 <= b(50) and w2428;
w18335 <= b(51) and w2277;
w18336 <= not w18334 and not w18335;
w18337 <= not w18333 and w18336;
w18338 <= not w2285 and w18337;
w18339 <= not w9371 and w18337;
w18340 <= not w18338 and not w18339;
w18341 <= a(26) and not w18340;
w18342 <= not a(26) and w18340;
w18343 <= not w18341 and not w18342;
w18344 <= not w18332 and not w18343;
w18345 <= w18332 and w18343;
w18346 <= not w18344 and not w18345;
w18347 <= not w18330 and w18346;
w18348 <= not w18330 and not w18347;
w18349 <= w18346 and not w18347;
w18350 <= not w18348 and not w18349;
w18351 <= not w18094 and not w18350;
w18352 <= not w18094 and not w18351;
w18353 <= not w18350 and not w18351;
w18354 <= not w18352 and not w18353;
w18355 <= not w17775 and not w18036;
w18356 <= b(58) and w1370;
w18357 <= b(56) and w1506;
w18358 <= b(57) and w1365;
w18359 <= not w18357 and not w18358;
w18360 <= not w18356 and w18359;
w18361 <= not w1373 and w18360;
w18362 <= not w11179 and w18360;
w18363 <= not w18361 and not w18362;
w18364 <= a(20) and not w18363;
w18365 <= not a(20) and w18363;
w18366 <= not w18364 and not w18365;
w18367 <= not w18355 and not w18366;
w18368 <= not w18355 and not w18367;
w18369 <= not w18366 and not w18367;
w18370 <= not w18368 and not w18369;
w18371 <= not w18354 and not w18370;
w18372 <= not w18354 and not w18371;
w18373 <= not w18370 and not w18371;
w18374 <= not w18372 and not w18373;
w18375 <= not w18078 and not w18374;
w18376 <= not w18078 and not w18375;
w18377 <= not w18374 and not w18375;
w18378 <= not w18376 and not w18377;
w18379 <= not w17733 and not w17744;
w18380 <= not w18044 and not w18379;
w18381 <= b(62) and w799;
w18382 <= b(63) and w689;
w18383 <= not w18381 and not w18382;
w18384 <= not w697 and w18383;
w18385 <= w13543 and w18383;
w18386 <= not w18384 and not w18385;
w18387 <= a(14) and not w18386;
w18388 <= not a(14) and w18386;
w18389 <= not w18387 and not w18388;
w18390 <= not w18380 and not w18389;
w18391 <= not w18380 and not w18390;
w18392 <= not w18389 and not w18390;
w18393 <= not w18391 and not w18392;
w18394 <= not w18378 and not w18393;
w18395 <= w18378 and not w18392;
w18396 <= not w18391 and w18395;
w18397 <= not w18394 and not w18396;
w18398 <= not w18062 and w18397;
w18399 <= not w18062 and not w18398;
w18400 <= w18397 and not w18398;
w18401 <= not w18399 and not w18400;
w18402 <= not w18060 and not w18401;
w18403 <= w18060 and not w18400;
w18404 <= not w18399 and w18403;
w18405 <= not w18402 and not w18404;
w18406 <= not w18398 and not w18402;
w18407 <= not w18390 and not w18394;
w18408 <= not w18075 and not w18375;
w18409 <= b(63) and w799;
w18410 <= w697 and w13540;
w18411 <= not w18409 and not w18410;
w18412 <= a(14) and not w18411;
w18413 <= a(14) and not w18412;
w18414 <= not w18411 and not w18412;
w18415 <= not w18413 and not w18414;
w18416 <= not w18408 and not w18415;
w18417 <= not w18408 and not w18416;
w18418 <= not w18415 and not w18416;
w18419 <= not w18417 and not w18418;
w18420 <= b(59) and w1370;
w18421 <= b(57) and w1506;
w18422 <= b(58) and w1365;
w18423 <= not w18421 and not w18422;
w18424 <= not w18420 and w18423;
w18425 <= w1373 and w11922;
w18426 <= w18424 and not w18425;
w18427 <= a(20) and not w18426;
w18428 <= a(20) and not w18427;
w18429 <= not w18426 and not w18427;
w18430 <= not w18428 and not w18429;
w18431 <= not w18091 and not w18351;
w18432 <= w18430 and w18431;
w18433 <= not w18430 and not w18431;
w18434 <= not w18432 and not w18433;
w18435 <= b(56) and w1791;
w18436 <= b(54) and w1941;
w18437 <= b(55) and w1786;
w18438 <= not w18436 and not w18437;
w18439 <= not w18435 and w18438;
w18440 <= w1794 and w10451;
w18441 <= w18439 and not w18440;
w18442 <= a(23) and not w18441;
w18443 <= a(23) and not w18442;
w18444 <= not w18441 and not w18442;
w18445 <= not w18443 and not w18444;
w18446 <= not w18344 and not w18347;
w18447 <= w18445 and w18446;
w18448 <= not w18445 and not w18446;
w18449 <= not w18447 and not w18448;
w18450 <= b(53) and w2282;
w18451 <= b(51) and w2428;
w18452 <= b(52) and w2277;
w18453 <= not w18451 and not w18452;
w18454 <= not w18450 and w18453;
w18455 <= w2285 and w9715;
w18456 <= w18454 and not w18455;
w18457 <= a(26) and not w18456;
w18458 <= a(26) and not w18457;
w18459 <= not w18456 and not w18457;
w18460 <= not w18458 and not w18459;
w18461 <= not w18107 and not w18327;
w18462 <= w18460 and w18461;
w18463 <= not w18460 and not w18461;
w18464 <= not w18462 and not w18463;
w18465 <= not w18300 and not w18303;
w18466 <= b(47) and w3381;
w18467 <= b(45) and w3586;
w18468 <= b(46) and w3376;
w18469 <= not w18467 and not w18468;
w18470 <= not w18466 and w18469;
w18471 <= not w3384 and w18470;
w18472 <= not w7446 and w18470;
w18473 <= not w18471 and not w18472;
w18474 <= a(32) and not w18473;
w18475 <= not a(32) and w18473;
w18476 <= not w18474 and not w18475;
w18477 <= not w18465 and not w18476;
w18478 <= w18465 and w18476;
w18479 <= not w18477 and not w18478;
w18480 <= b(44) and w4030;
w18481 <= b(42) and w4275;
w18482 <= b(43) and w4025;
w18483 <= not w18481 and not w18482;
w18484 <= not w18480 and w18483;
w18485 <= w4033 and w6815;
w18486 <= w18484 and not w18485;
w18487 <= a(35) and not w18486;
w18488 <= a(35) and not w18487;
w18489 <= not w18486 and not w18487;
w18490 <= not w18488 and not w18489;
w18491 <= not w18292 and not w18296;
w18492 <= b(41) and w4778;
w18493 <= b(39) and w5020;
w18494 <= b(40) and w4773;
w18495 <= not w18493 and not w18494;
w18496 <= not w18492 and w18495;
w18497 <= w4781 and w5962;
w18498 <= w18496 and not w18497;
w18499 <= a(38) and not w18498;
w18500 <= a(38) and not w18499;
w18501 <= not w18498 and not w18499;
w18502 <= not w18500 and not w18501;
w18503 <= not w18284 and not w18288;
w18504 <= not w18270 and not w18274;
w18505 <= not w18235 and not w18248;
w18506 <= b(26) and w9082;
w18507 <= b(24) and w9475;
w18508 <= b(25) and w9077;
w18509 <= not w18507 and not w18508;
w18510 <= not w18506 and w18509;
w18511 <= w2556 and w9085;
w18512 <= w18510 and not w18511;
w18513 <= a(53) and not w18512;
w18514 <= a(53) and not w18513;
w18515 <= not w18512 and not w18513;
w18516 <= not w18514 and not w18515;
w18517 <= not w18216 and not w18229;
w18518 <= not w18180 and not w18191;
w18519 <= not w18177 and not w18518;
w18520 <= b(13) and w13646;
w18521 <= b(14) and not w13231;
w18522 <= not w18520 and not w18521;
w18523 <= w18174 and not w18522;
w18524 <= not w18174 and w18522;
w18525 <= not w18523 and not w18524;
w18526 <= b(17) and w12411;
w18527 <= b(15) and w12790;
w18528 <= b(16) and w12406;
w18529 <= not w18527 and not w18528;
w18530 <= not w18526 and w18529;
w18531 <= not w12414 and w18530;
w18532 <= not w1099 and w18530;
w18533 <= not w18531 and not w18532;
w18534 <= a(62) and not w18533;
w18535 <= not a(62) and w18533;
w18536 <= not w18534 and not w18535;
w18537 <= w18525 and not w18536;
w18538 <= not w18525 and w18536;
w18539 <= not w18537 and not w18538;
w18540 <= not w18519 and w18539;
w18541 <= w18519 and not w18539;
w18542 <= not w18540 and not w18541;
w18543 <= b(20) and w11274;
w18544 <= b(18) and w11639;
w18545 <= b(19) and w11269;
w18546 <= not w18544 and not w18545;
w18547 <= not w18543 and w18546;
w18548 <= w1589 and w11277;
w18549 <= w18547 and not w18548;
w18550 <= a(59) and not w18549;
w18551 <= a(59) and not w18550;
w18552 <= not w18549 and not w18550;
w18553 <= not w18551 and not w18552;
w18554 <= w18542 and not w18553;
w18555 <= w18542 and not w18554;
w18556 <= not w18553 and not w18554;
w18557 <= not w18555 and not w18556;
w18558 <= not w18197 and not w18210;
w18559 <= w18557 and w18558;
w18560 <= not w18557 and not w18558;
w18561 <= not w18559 and not w18560;
w18562 <= b(23) and w10169;
w18563 <= b(21) and w10539;
w18564 <= b(22) and w10164;
w18565 <= not w18563 and not w18564;
w18566 <= not w18562 and w18565;
w18567 <= w2043 and w10172;
w18568 <= w18566 and not w18567;
w18569 <= a(56) and not w18568;
w18570 <= a(56) and not w18569;
w18571 <= not w18568 and not w18569;
w18572 <= not w18570 and not w18571;
w18573 <= not w18561 and w18572;
w18574 <= w18561 and not w18572;
w18575 <= not w18573 and not w18574;
w18576 <= not w18517 and w18575;
w18577 <= w18517 and not w18575;
w18578 <= not w18576 and not w18577;
w18579 <= not w18516 and w18578;
w18580 <= w18516 and not w18578;
w18581 <= not w18579 and not w18580;
w18582 <= not w18505 and w18581;
w18583 <= w18505 and not w18581;
w18584 <= not w18582 and not w18583;
w18585 <= b(29) and w8105;
w18586 <= b(27) and w8458;
w18587 <= b(28) and w8100;
w18588 <= not w18586 and not w18587;
w18589 <= not w18585 and w18588;
w18590 <= w3126 and w8108;
w18591 <= w18589 and not w18590;
w18592 <= a(50) and not w18591;
w18593 <= a(50) and not w18592;
w18594 <= not w18591 and not w18592;
w18595 <= not w18593 and not w18594;
w18596 <= w18584 and not w18595;
w18597 <= w18584 and not w18596;
w18598 <= not w18595 and not w18596;
w18599 <= not w18597 and not w18598;
w18600 <= not w18254 and not w18268;
w18601 <= not w18599 and not w18600;
w18602 <= not w18599 and not w18601;
w18603 <= not w18600 and not w18601;
w18604 <= not w18602 and not w18603;
w18605 <= b(32) and w7189;
w18606 <= b(30) and w7530;
w18607 <= b(31) and w7184;
w18608 <= not w18606 and not w18607;
w18609 <= not w18605 and w18608;
w18610 <= w3756 and w7192;
w18611 <= w18609 and not w18610;
w18612 <= a(47) and not w18611;
w18613 <= a(47) and not w18612;
w18614 <= not w18611 and not w18612;
w18615 <= not w18613 and not w18614;
w18616 <= not w18604 and w18615;
w18617 <= w18604 and not w18615;
w18618 <= not w18616 and not w18617;
w18619 <= w18504 and w18618;
w18620 <= not w18504 and not w18618;
w18621 <= not w18619 and not w18620;
w18622 <= b(35) and w6338;
w18623 <= b(33) and w6645;
w18624 <= b(34) and w6333;
w18625 <= not w18623 and not w18624;
w18626 <= not w18622 and w18625;
w18627 <= w4439 and w6341;
w18628 <= w18626 and not w18627;
w18629 <= a(44) and not w18628;
w18630 <= a(44) and not w18629;
w18631 <= not w18628 and not w18629;
w18632 <= not w18630 and not w18631;
w18633 <= w18621 and not w18632;
w18634 <= w18621 and not w18633;
w18635 <= not w18632 and not w18633;
w18636 <= not w18634 and not w18635;
w18637 <= not w18278 and not w18281;
w18638 <= w18636 and w18637;
w18639 <= not w18636 and not w18637;
w18640 <= not w18638 and not w18639;
w18641 <= b(38) and w5520;
w18642 <= b(36) and w5802;
w18643 <= b(37) and w5515;
w18644 <= not w18642 and not w18643;
w18645 <= not w18641 and w18644;
w18646 <= w4948 and w5523;
w18647 <= w18645 and not w18646;
w18648 <= a(41) and not w18647;
w18649 <= a(41) and not w18648;
w18650 <= not w18647 and not w18648;
w18651 <= not w18649 and not w18650;
w18652 <= not w18640 and w18651;
w18653 <= w18640 and not w18651;
w18654 <= not w18652 and not w18653;
w18655 <= not w18503 and w18654;
w18656 <= w18503 and not w18654;
w18657 <= not w18655 and not w18656;
w18658 <= not w18502 and w18657;
w18659 <= w18502 and not w18657;
w18660 <= not w18658 and not w18659;
w18661 <= not w18491 and w18660;
w18662 <= w18491 and not w18660;
w18663 <= not w18661 and not w18662;
w18664 <= not w18490 and w18663;
w18665 <= not w18490 and not w18664;
w18666 <= w18663 and not w18664;
w18667 <= not w18665 and not w18666;
w18668 <= w18479 and not w18667;
w18669 <= w18479 and not w18668;
w18670 <= not w18667 and not w18668;
w18671 <= not w18669 and not w18670;
w18672 <= not w18319 and not w18323;
w18673 <= b(50) and w2793;
w18674 <= b(48) and w2986;
w18675 <= b(49) and w2788;
w18676 <= not w18674 and not w18675;
w18677 <= not w18673 and w18676;
w18678 <= not w2796 and w18677;
w18679 <= not w8692 and w18677;
w18680 <= not w18678 and not w18679;
w18681 <= a(29) and not w18680;
w18682 <= not a(29) and w18680;
w18683 <= not w18681 and not w18682;
w18684 <= not w18672 and not w18683;
w18685 <= w18672 and w18683;
w18686 <= not w18684 and not w18685;
w18687 <= not w18671 and w18686;
w18688 <= not w18671 and not w18687;
w18689 <= w18686 and not w18687;
w18690 <= not w18688 and not w18689;
w18691 <= w18464 and not w18690;
w18692 <= w18464 and not w18691;
w18693 <= not w18690 and not w18691;
w18694 <= not w18692 and not w18693;
w18695 <= w18449 and not w18694;
w18696 <= not w18449 and w18694;
w18697 <= w18434 and not w18696;
w18698 <= not w18695 and w18697;
w18699 <= w18434 and not w18698;
w18700 <= not w18696 and not w18698;
w18701 <= not w18695 and w18700;
w18702 <= not w18699 and not w18701;
w18703 <= not w18367 and not w18371;
w18704 <= b(62) and w1045;
w18705 <= b(60) and w1134;
w18706 <= b(61) and w1040;
w18707 <= not w18705 and not w18706;
w18708 <= not w18704 and w18707;
w18709 <= not w1048 and w18708;
w18710 <= not w13113 and w18708;
w18711 <= not w18709 and not w18710;
w18712 <= a(17) and not w18711;
w18713 <= not a(17) and w18711;
w18714 <= not w18712 and not w18713;
w18715 <= not w18703 and not w18714;
w18716 <= not w18703 and not w18715;
w18717 <= not w18714 and not w18715;
w18718 <= not w18716 and not w18717;
w18719 <= not w18702 and not w18718;
w18720 <= w18702 and not w18717;
w18721 <= not w18716 and w18720;
w18722 <= not w18719 and not w18721;
w18723 <= not w18419 and w18722;
w18724 <= w18419 and not w18722;
w18725 <= not w18723 and not w18724;
w18726 <= not w18407 and w18725;
w18727 <= w18407 and not w18725;
w18728 <= not w18726 and not w18727;
w18729 <= not w18406 and w18728;
w18730 <= w18406 and not w18728;
w18731 <= not w18729 and not w18730;
w18732 <= not w18715 and not w18719;
w18733 <= b(63) and w1045;
w18734 <= b(61) and w1134;
w18735 <= b(62) and w1040;
w18736 <= not w18734 and not w18735;
w18737 <= not w18733 and w18736;
w18738 <= w1048 and w13514;
w18739 <= w18737 and not w18738;
w18740 <= a(17) and not w18739;
w18741 <= a(17) and not w18740;
w18742 <= not w18739 and not w18740;
w18743 <= not w18741 and not w18742;
w18744 <= not w18732 and not w18743;
w18745 <= not w18732 and not w18744;
w18746 <= not w18743 and not w18744;
w18747 <= not w18745 and not w18746;
w18748 <= b(60) and w1370;
w18749 <= b(58) and w1506;
w18750 <= b(59) and w1365;
w18751 <= not w18749 and not w18750;
w18752 <= not w18748 and w18751;
w18753 <= w1373 and w11954;
w18754 <= w18752 and not w18753;
w18755 <= a(20) and not w18754;
w18756 <= a(20) and not w18755;
w18757 <= not w18754 and not w18755;
w18758 <= not w18756 and not w18757;
w18759 <= not w18433 and not w18698;
w18760 <= w18758 and w18759;
w18761 <= not w18758 and not w18759;
w18762 <= not w18760 and not w18761;
w18763 <= not w18448 and not w18695;
w18764 <= b(57) and w1791;
w18765 <= b(55) and w1941;
w18766 <= b(56) and w1786;
w18767 <= not w18765 and not w18766;
w18768 <= not w18764 and w18767;
w18769 <= w1794 and w11153;
w18770 <= w18768 and not w18769;
w18771 <= a(23) and not w18770;
w18772 <= a(23) and not w18771;
w18773 <= not w18770 and not w18771;
w18774 <= not w18772 and not w18773;
w18775 <= not w18763 and w18774;
w18776 <= w18763 and not w18774;
w18777 <= not w18775 and not w18776;
w18778 <= b(54) and w2282;
w18779 <= b(52) and w2428;
w18780 <= b(53) and w2277;
w18781 <= not w18779 and not w18780;
w18782 <= not w18778 and w18781;
w18783 <= w2285 and w9741;
w18784 <= w18782 and not w18783;
w18785 <= a(26) and not w18784;
w18786 <= a(26) and not w18785;
w18787 <= not w18784 and not w18785;
w18788 <= not w18786 and not w18787;
w18789 <= not w18463 and not w18691;
w18790 <= w18788 and w18789;
w18791 <= not w18788 and not w18789;
w18792 <= not w18790 and not w18791;
w18793 <= b(51) and w2793;
w18794 <= b(49) and w2986;
w18795 <= b(50) and w2788;
w18796 <= not w18794 and not w18795;
w18797 <= not w18793 and w18796;
w18798 <= w2796 and w8719;
w18799 <= w18797 and not w18798;
w18800 <= a(29) and not w18799;
w18801 <= a(29) and not w18800;
w18802 <= not w18799 and not w18800;
w18803 <= not w18801 and not w18802;
w18804 <= not w18684 and not w18687;
w18805 <= w18803 and w18804;
w18806 <= not w18803 and not w18804;
w18807 <= not w18805 and not w18806;
w18808 <= not w18655 and not w18658;
w18809 <= not w18639 and not w18653;
w18810 <= not w18620 and not w18633;
w18811 <= not w18604 and not w18615;
w18812 <= not w18601 and not w18811;
w18813 <= not w18560 and not w18574;
w18814 <= b(14) and w13646;
w18815 <= b(15) and not w13231;
w18816 <= not w18814 and not w18815;
w18817 <= not a(14) and not w18816;
w18818 <= not a(14) and not w18817;
w18819 <= not w18816 and not w18817;
w18820 <= not w18818 and not w18819;
w18821 <= not w18174 and not w18820;
w18822 <= not w18174 and not w18821;
w18823 <= not w18820 and not w18821;
w18824 <= not w18822 and not w18823;
w18825 <= b(18) and w12411;
w18826 <= b(16) and w12790;
w18827 <= b(17) and w12406;
w18828 <= not w18826 and not w18827;
w18829 <= not w18825 and w18828;
w18830 <= w1309 and w12414;
w18831 <= w18829 and not w18830;
w18832 <= a(62) and not w18831;
w18833 <= a(62) and not w18832;
w18834 <= not w18831 and not w18832;
w18835 <= not w18833 and not w18834;
w18836 <= not w18824 and not w18835;
w18837 <= not w18824 and not w18836;
w18838 <= not w18835 and not w18836;
w18839 <= not w18837 and not w18838;
w18840 <= not w18523 and not w18537;
w18841 <= w18839 and w18840;
w18842 <= not w18839 and not w18840;
w18843 <= not w18841 and not w18842;
w18844 <= b(21) and w11274;
w18845 <= b(19) and w11639;
w18846 <= b(20) and w11269;
w18847 <= not w18845 and not w18846;
w18848 <= not w18844 and w18847;
w18849 <= w1727 and w11277;
w18850 <= w18848 and not w18849;
w18851 <= a(59) and not w18850;
w18852 <= a(59) and not w18851;
w18853 <= not w18850 and not w18851;
w18854 <= not w18852 and not w18853;
w18855 <= w18843 and not w18854;
w18856 <= w18843 and not w18855;
w18857 <= not w18854 and not w18855;
w18858 <= not w18856 and not w18857;
w18859 <= not w18540 and not w18554;
w18860 <= w18858 and w18859;
w18861 <= not w18858 and not w18859;
w18862 <= not w18860 and not w18861;
w18863 <= b(24) and w10169;
w18864 <= b(22) and w10539;
w18865 <= b(23) and w10164;
w18866 <= not w18864 and not w18865;
w18867 <= not w18863 and w18866;
w18868 <= w2201 and w10172;
w18869 <= w18867 and not w18868;
w18870 <= a(56) and not w18869;
w18871 <= a(56) and not w18870;
w18872 <= not w18869 and not w18870;
w18873 <= not w18871 and not w18872;
w18874 <= w18862 and not w18873;
w18875 <= not w18862 and w18873;
w18876 <= not w18813 and not w18875;
w18877 <= not w18874 and w18876;
w18878 <= not w18813 and not w18877;
w18879 <= not w18874 and not w18877;
w18880 <= not w18875 and w18879;
w18881 <= not w18878 and not w18880;
w18882 <= b(27) and w9082;
w18883 <= b(25) and w9475;
w18884 <= b(26) and w9077;
w18885 <= not w18883 and not w18884;
w18886 <= not w18882 and w18885;
w18887 <= w2733 and w9085;
w18888 <= w18886 and not w18887;
w18889 <= a(53) and not w18888;
w18890 <= a(53) and not w18889;
w18891 <= not w18888 and not w18889;
w18892 <= not w18890 and not w18891;
w18893 <= not w18881 and not w18892;
w18894 <= not w18881 and not w18893;
w18895 <= not w18892 and not w18893;
w18896 <= not w18894 and not w18895;
w18897 <= not w18576 and not w18579;
w18898 <= w18896 and w18897;
w18899 <= not w18896 and not w18897;
w18900 <= not w18898 and not w18899;
w18901 <= b(30) and w8105;
w18902 <= b(28) and w8458;
w18903 <= b(29) and w8100;
w18904 <= not w18902 and not w18903;
w18905 <= not w18901 and w18904;
w18906 <= w3320 and w8108;
w18907 <= w18905 and not w18906;
w18908 <= a(50) and not w18907;
w18909 <= a(50) and not w18908;
w18910 <= not w18907 and not w18908;
w18911 <= not w18909 and not w18910;
w18912 <= w18900 and not w18911;
w18913 <= w18900 and not w18912;
w18914 <= not w18911 and not w18912;
w18915 <= not w18913 and not w18914;
w18916 <= not w18582 and not w18596;
w18917 <= w18915 and w18916;
w18918 <= not w18915 and not w18916;
w18919 <= not w18917 and not w18918;
w18920 <= b(33) and w7189;
w18921 <= b(31) and w7530;
w18922 <= b(32) and w7184;
w18923 <= not w18921 and not w18922;
w18924 <= not w18920 and w18923;
w18925 <= w3966 and w7192;
w18926 <= w18924 and not w18925;
w18927 <= a(47) and not w18926;
w18928 <= a(47) and not w18927;
w18929 <= not w18926 and not w18927;
w18930 <= not w18928 and not w18929;
w18931 <= w18919 and not w18930;
w18932 <= w18919 and not w18931;
w18933 <= not w18930 and not w18931;
w18934 <= not w18932 and not w18933;
w18935 <= not w18812 and w18934;
w18936 <= w18812 and not w18934;
w18937 <= not w18935 and not w18936;
w18938 <= b(36) and w6338;
w18939 <= b(34) and w6645;
w18940 <= b(35) and w6333;
w18941 <= not w18939 and not w18940;
w18942 <= not w18938 and w18941;
w18943 <= w4665 and w6341;
w18944 <= w18942 and not w18943;
w18945 <= a(44) and not w18944;
w18946 <= a(44) and not w18945;
w18947 <= not w18944 and not w18945;
w18948 <= not w18946 and not w18947;
w18949 <= not w18937 and not w18948;
w18950 <= w18937 and w18948;
w18951 <= not w18949 and not w18950;
w18952 <= w18810 and not w18951;
w18953 <= not w18810 and w18951;
w18954 <= not w18952 and not w18953;
w18955 <= b(39) and w5520;
w18956 <= b(37) and w5802;
w18957 <= b(38) and w5515;
w18958 <= not w18956 and not w18957;
w18959 <= not w18955 and w18958;
w18960 <= w5194 and w5523;
w18961 <= w18959 and not w18960;
w18962 <= a(41) and not w18961;
w18963 <= a(41) and not w18962;
w18964 <= not w18961 and not w18962;
w18965 <= not w18963 and not w18964;
w18966 <= w18954 and not w18965;
w18967 <= w18954 and not w18966;
w18968 <= not w18965 and not w18966;
w18969 <= not w18967 and not w18968;
w18970 <= not w18809 and w18969;
w18971 <= w18809 and not w18969;
w18972 <= not w18970 and not w18971;
w18973 <= b(42) and w4778;
w18974 <= b(40) and w5020;
w18975 <= b(41) and w4773;
w18976 <= not w18974 and not w18975;
w18977 <= not w18973 and w18976;
w18978 <= w4781 and w6232;
w18979 <= w18977 and not w18978;
w18980 <= a(38) and not w18979;
w18981 <= a(38) and not w18980;
w18982 <= not w18979 and not w18980;
w18983 <= not w18981 and not w18982;
w18984 <= not w18972 and not w18983;
w18985 <= w18972 and w18983;
w18986 <= not w18984 and not w18985;
w18987 <= w18808 and not w18986;
w18988 <= not w18808 and w18986;
w18989 <= not w18987 and not w18988;
w18990 <= b(45) and w4030;
w18991 <= b(43) and w4275;
w18992 <= b(44) and w4025;
w18993 <= not w18991 and not w18992;
w18994 <= not w18990 and w18993;
w18995 <= w4033 and w7104;
w18996 <= w18994 and not w18995;
w18997 <= a(35) and not w18996;
w18998 <= a(35) and not w18997;
w18999 <= not w18996 and not w18997;
w19000 <= not w18998 and not w18999;
w19001 <= w18989 and not w19000;
w19002 <= w18989 and not w19001;
w19003 <= not w19000 and not w19001;
w19004 <= not w19002 and not w19003;
w19005 <= not w18661 and not w18664;
w19006 <= w19004 and w19005;
w19007 <= not w19004 and not w19005;
w19008 <= not w19006 and not w19007;
w19009 <= not w18477 and not w18668;
w19010 <= b(48) and w3381;
w19011 <= b(46) and w3586;
w19012 <= b(47) and w3376;
w19013 <= not w19011 and not w19012;
w19014 <= not w19010 and w19013;
w19015 <= w3384 and w7752;
w19016 <= w19014 and not w19015;
w19017 <= a(32) and not w19016;
w19018 <= a(32) and not w19017;
w19019 <= not w19016 and not w19017;
w19020 <= not w19018 and not w19019;
w19021 <= not w19009 and not w19020;
w19022 <= not w19009 and not w19021;
w19023 <= not w19020 and not w19021;
w19024 <= not w19022 and not w19023;
w19025 <= w19008 and not w19024;
w19026 <= not w19008 and w19024;
w19027 <= w18807 and not w19026;
w19028 <= not w19025 and w19027;
w19029 <= w18807 and not w19028;
w19030 <= not w19026 and not w19028;
w19031 <= not w19025 and w19030;
w19032 <= not w19029 and not w19031;
w19033 <= w18792 and not w19032;
w19034 <= not w18792 and w19032;
w19035 <= not w18777 and not w19034;
w19036 <= not w19033 and w19035;
w19037 <= not w18777 and not w19036;
w19038 <= not w19034 and not w19036;
w19039 <= not w19033 and w19038;
w19040 <= not w19037 and not w19039;
w19041 <= w18762 and not w19040;
w19042 <= not w18762 and w19040;
w19043 <= not w18747 and not w19042;
w19044 <= not w19041 and w19043;
w19045 <= not w18747 and not w19044;
w19046 <= not w19042 and not w19044;
w19047 <= not w19041 and w19046;
w19048 <= not w19045 and not w19047;
w19049 <= not w18416 and not w18723;
w19050 <= w19048 and w19049;
w19051 <= not w19048 and not w19049;
w19052 <= not w19050 and not w19051;
w19053 <= not w18726 and not w18729;
w19054 <= w19052 and not w19053;
w19055 <= not w19052 and w19053;
w19056 <= not w19054 and not w19055;
w19057 <= not w18761 and not w19041;
w19058 <= b(62) and w1134;
w19059 <= b(63) and w1040;
w19060 <= not w19058 and not w19059;
w19061 <= not w1048 and w19060;
w19062 <= w13543 and w19060;
w19063 <= not w19061 and not w19062;
w19064 <= a(17) and not w19063;
w19065 <= not a(17) and w19063;
w19066 <= not w19064 and not w19065;
w19067 <= not w19057 and not w19066;
w19068 <= w19057 and w19066;
w19069 <= not w19067 and not w19068;
w19070 <= b(61) and w1370;
w19071 <= b(59) and w1506;
w19072 <= b(60) and w1365;
w19073 <= not w19071 and not w19072;
w19074 <= not w19070 and w19073;
w19075 <= w1373 and w12712;
w19076 <= w19074 and not w19075;
w19077 <= a(20) and not w19076;
w19078 <= a(20) and not w19077;
w19079 <= not w19076 and not w19077;
w19080 <= not w19078 and not w19079;
w19081 <= not w18763 and not w18774;
w19082 <= not w19036 and not w19081;
w19083 <= w19080 and w19082;
w19084 <= not w19080 and not w19082;
w19085 <= not w19083 and not w19084;
w19086 <= not w18791 and not w19033;
w19087 <= b(58) and w1791;
w19088 <= b(56) and w1941;
w19089 <= b(57) and w1786;
w19090 <= not w19088 and not w19089;
w19091 <= not w19087 and w19090;
w19092 <= not w1794 and w19091;
w19093 <= not w11179 and w19091;
w19094 <= not w19092 and not w19093;
w19095 <= a(23) and not w19094;
w19096 <= not a(23) and w19094;
w19097 <= not w19095 and not w19096;
w19098 <= not w19086 and not w19097;
w19099 <= w19086 and w19097;
w19100 <= not w19098 and not w19099;
w19101 <= b(55) and w2282;
w19102 <= b(53) and w2428;
w19103 <= b(54) and w2277;
w19104 <= not w19102 and not w19103;
w19105 <= not w19101 and w19104;
w19106 <= w2285 and w10427;
w19107 <= w19105 and not w19106;
w19108 <= a(26) and not w19107;
w19109 <= a(26) and not w19108;
w19110 <= not w19107 and not w19108;
w19111 <= not w19109 and not w19110;
w19112 <= not w18806 and not w19028;
w19113 <= w19111 and w19112;
w19114 <= not w19111 and not w19112;
w19115 <= not w19113 and not w19114;
w19116 <= b(52) and w2793;
w19117 <= b(50) and w2986;
w19118 <= b(51) and w2788;
w19119 <= not w19117 and not w19118;
w19120 <= not w19116 and w19119;
w19121 <= w2796 and w9371;
w19122 <= w19120 and not w19121;
w19123 <= a(29) and not w19122;
w19124 <= a(29) and not w19123;
w19125 <= not w19122 and not w19123;
w19126 <= not w19124 and not w19125;
w19127 <= not w19021 and not w19025;
w19128 <= not w19126 and not w19127;
w19129 <= not w19126 and not w19128;
w19130 <= not w19127 and not w19128;
w19131 <= not w19129 and not w19130;
w19132 <= b(49) and w3381;
w19133 <= b(47) and w3586;
w19134 <= b(48) and w3376;
w19135 <= not w19133 and not w19134;
w19136 <= not w19132 and w19135;
w19137 <= w3384 and w8368;
w19138 <= w19136 and not w19137;
w19139 <= a(32) and not w19138;
w19140 <= a(32) and not w19139;
w19141 <= not w19138 and not w19139;
w19142 <= not w19140 and not w19141;
w19143 <= not w19001 and not w19007;
w19144 <= w19142 and w19143;
w19145 <= not w19142 and not w19143;
w19146 <= not w19144 and not w19145;
w19147 <= b(43) and w4778;
w19148 <= b(41) and w5020;
w19149 <= b(42) and w4773;
w19150 <= not w19148 and not w19149;
w19151 <= not w19147 and w19150;
w19152 <= w4781 and w6258;
w19153 <= w19151 and not w19152;
w19154 <= a(38) and not w19153;
w19155 <= a(38) and not w19154;
w19156 <= not w19153 and not w19154;
w19157 <= not w19155 and not w19156;
w19158 <= not w18809 and not w18969;
w19159 <= not w18966 and not w19158;
w19160 <= b(40) and w5520;
w19161 <= b(38) and w5802;
w19162 <= b(39) and w5515;
w19163 <= not w19161 and not w19162;
w19164 <= not w19160 and w19163;
w19165 <= w5523 and w5698;
w19166 <= w19164 and not w19165;
w19167 <= a(41) and not w19166;
w19168 <= a(41) and not w19167;
w19169 <= not w19166 and not w19167;
w19170 <= not w19168 and not w19169;
w19171 <= not w18949 and not w18953;
w19172 <= b(37) and w6338;
w19173 <= b(35) and w6645;
w19174 <= b(36) and w6333;
w19175 <= not w19173 and not w19174;
w19176 <= not w19172 and w19175;
w19177 <= w4924 and w6341;
w19178 <= w19176 and not w19177;
w19179 <= a(44) and not w19178;
w19180 <= a(44) and not w19179;
w19181 <= not w19178 and not w19179;
w19182 <= not w19180 and not w19181;
w19183 <= not w18812 and not w18934;
w19184 <= not w18931 and not w19183;
w19185 <= b(31) and w8105;
w19186 <= b(29) and w8458;
w19187 <= b(30) and w8100;
w19188 <= not w19186 and not w19187;
w19189 <= not w19185 and w19188;
w19190 <= w3539 and w8108;
w19191 <= w19189 and not w19190;
w19192 <= a(50) and not w19191;
w19193 <= a(50) and not w19192;
w19194 <= not w19191 and not w19192;
w19195 <= not w19193 and not w19194;
w19196 <= not w18836 and not w18842;
w19197 <= b(15) and w13646;
w19198 <= b(16) and not w13231;
w19199 <= not w19197 and not w19198;
w19200 <= not w18817 and not w18821;
w19201 <= not w19199 and w19200;
w19202 <= w19199 and not w19200;
w19203 <= not w19201 and not w19202;
w19204 <= b(19) and w12411;
w19205 <= b(17) and w12790;
w19206 <= b(18) and w12406;
w19207 <= not w19205 and not w19206;
w19208 <= not w19204 and w19207;
w19209 <= not w12414 and w19208;
w19210 <= not w1451 and w19208;
w19211 <= not w19209 and not w19210;
w19212 <= a(62) and not w19211;
w19213 <= not a(62) and w19211;
w19214 <= not w19212 and not w19213;
w19215 <= w19203 and not w19214;
w19216 <= not w19203 and w19214;
w19217 <= not w19215 and not w19216;
w19218 <= not w19196 and w19217;
w19219 <= w19196 and not w19217;
w19220 <= not w19218 and not w19219;
w19221 <= b(22) and w11274;
w19222 <= b(20) and w11639;
w19223 <= b(21) and w11269;
w19224 <= not w19222 and not w19223;
w19225 <= not w19221 and w19224;
w19226 <= w1888 and w11277;
w19227 <= w19225 and not w19226;
w19228 <= a(59) and not w19227;
w19229 <= a(59) and not w19228;
w19230 <= not w19227 and not w19228;
w19231 <= not w19229 and not w19230;
w19232 <= w19220 and not w19231;
w19233 <= w19220 and not w19232;
w19234 <= not w19231 and not w19232;
w19235 <= not w19233 and not w19234;
w19236 <= not w18855 and not w18861;
w19237 <= w19235 and w19236;
w19238 <= not w19235 and not w19236;
w19239 <= not w19237 and not w19238;
w19240 <= b(25) and w10169;
w19241 <= b(23) and w10539;
w19242 <= b(24) and w10164;
w19243 <= not w19241 and not w19242;
w19244 <= not w19240 and w19243;
w19245 <= w2228 and w10172;
w19246 <= w19244 and not w19245;
w19247 <= a(56) and not w19246;
w19248 <= a(56) and not w19247;
w19249 <= not w19246 and not w19247;
w19250 <= not w19248 and not w19249;
w19251 <= w19239 and not w19250;
w19252 <= w19239 and not w19251;
w19253 <= not w19250 and not w19251;
w19254 <= not w19252 and not w19253;
w19255 <= not w18879 and w19254;
w19256 <= w18879 and not w19254;
w19257 <= not w19255 and not w19256;
w19258 <= b(28) and w9082;
w19259 <= b(26) and w9475;
w19260 <= b(27) and w9077;
w19261 <= not w19259 and not w19260;
w19262 <= not w19258 and w19261;
w19263 <= w2932 and w9085;
w19264 <= w19262 and not w19263;
w19265 <= a(53) and not w19264;
w19266 <= a(53) and not w19265;
w19267 <= not w19264 and not w19265;
w19268 <= not w19266 and not w19267;
w19269 <= w19257 and w19268;
w19270 <= not w19257 and not w19268;
w19271 <= not w19269 and not w19270;
w19272 <= not w18893 and not w18899;
w19273 <= w19271 and not w19272;
w19274 <= not w19271 and w19272;
w19275 <= not w19273 and not w19274;
w19276 <= not w19195 and w19275;
w19277 <= w19275 and not w19276;
w19278 <= not w19195 and not w19276;
w19279 <= not w19277 and not w19278;
w19280 <= not w18912 and not w18918;
w19281 <= w19279 and w19280;
w19282 <= not w19279 and not w19280;
w19283 <= not w19281 and not w19282;
w19284 <= b(34) and w7189;
w19285 <= b(32) and w7530;
w19286 <= b(33) and w7184;
w19287 <= not w19285 and not w19286;
w19288 <= not w19284 and w19287;
w19289 <= w4209 and w7192;
w19290 <= w19288 and not w19289;
w19291 <= a(47) and not w19290;
w19292 <= a(47) and not w19291;
w19293 <= not w19290 and not w19291;
w19294 <= not w19292 and not w19293;
w19295 <= not w19283 and w19294;
w19296 <= w19283 and not w19294;
w19297 <= not w19295 and not w19296;
w19298 <= not w19184 and w19297;
w19299 <= not w19184 and not w19298;
w19300 <= w19297 and not w19298;
w19301 <= not w19299 and not w19300;
w19302 <= not w19182 and not w19301;
w19303 <= w19182 and not w19300;
w19304 <= not w19299 and w19303;
w19305 <= not w19302 and not w19304;
w19306 <= not w19171 and w19305;
w19307 <= not w19171 and not w19306;
w19308 <= w19305 and not w19306;
w19309 <= not w19307 and not w19308;
w19310 <= not w19170 and not w19309;
w19311 <= w19170 and not w19308;
w19312 <= not w19307 and w19311;
w19313 <= not w19310 and not w19312;
w19314 <= not w19159 and w19313;
w19315 <= w19159 and not w19313;
w19316 <= not w19314 and not w19315;
w19317 <= not w19157 and w19316;
w19318 <= w19316 and not w19317;
w19319 <= not w19157 and not w19317;
w19320 <= not w19318 and not w19319;
w19321 <= not w18984 and not w18988;
w19322 <= w19320 and w19321;
w19323 <= not w19320 and not w19321;
w19324 <= not w19322 and not w19323;
w19325 <= b(46) and w4030;
w19326 <= b(44) and w4275;
w19327 <= b(45) and w4025;
w19328 <= not w19326 and not w19327;
w19329 <= not w19325 and w19328;
w19330 <= w4033 and w7420;
w19331 <= w19329 and not w19330;
w19332 <= a(35) and not w19331;
w19333 <= a(35) and not w19332;
w19334 <= not w19331 and not w19332;
w19335 <= not w19333 and not w19334;
w19336 <= w19324 and not w19335;
w19337 <= w19324 and not w19336;
w19338 <= not w19335 and not w19336;
w19339 <= not w19337 and not w19338;
w19340 <= w19146 and not w19339;
w19341 <= not w19146 and w19339;
w19342 <= not w19131 and not w19341;
w19343 <= not w19340 and w19342;
w19344 <= not w19131 and not w19343;
w19345 <= not w19341 and not w19343;
w19346 <= not w19340 and w19345;
w19347 <= not w19344 and not w19346;
w19348 <= w19115 and not w19347;
w19349 <= not w19115 and w19347;
w19350 <= w19100 and not w19349;
w19351 <= not w19348 and w19350;
w19352 <= w19100 and not w19351;
w19353 <= not w19349 and not w19351;
w19354 <= not w19348 and w19353;
w19355 <= not w19352 and not w19354;
w19356 <= w19085 and not w19355;
w19357 <= not w19085 and w19355;
w19358 <= w19069 and not w19357;
w19359 <= not w19356 and w19358;
w19360 <= w19069 and not w19359;
w19361 <= not w19357 and not w19359;
w19362 <= not w19356 and w19361;
w19363 <= not w19360 and not w19362;
w19364 <= not w18744 and not w19044;
w19365 <= w19363 and w19364;
w19366 <= not w19363 and not w19364;
w19367 <= not w19365 and not w19366;
w19368 <= not w19051 and not w19054;
w19369 <= w19367 and not w19368;
w19370 <= not w19367 and w19368;
w19371 <= not w19369 and not w19370;
w19372 <= not w19366 and not w19369;
w19373 <= not w19067 and not w19359;
w19374 <= not w19084 and not w19356;
w19375 <= b(63) and w1134;
w19376 <= w1048 and w13540;
w19377 <= not w19375 and not w19376;
w19378 <= a(17) and not w19377;
w19379 <= a(17) and not w19378;
w19380 <= not w19377 and not w19378;
w19381 <= not w19379 and not w19380;
w19382 <= not w19374 and not w19381;
w19383 <= not w19374 and not w19382;
w19384 <= not w19381 and not w19382;
w19385 <= not w19383 and not w19384;
w19386 <= b(62) and w1370;
w19387 <= b(60) and w1506;
w19388 <= b(61) and w1365;
w19389 <= not w19387 and not w19388;
w19390 <= not w19386 and w19389;
w19391 <= w1373 and w13113;
w19392 <= w19390 and not w19391;
w19393 <= a(20) and not w19392;
w19394 <= a(20) and not w19393;
w19395 <= not w19392 and not w19393;
w19396 <= not w19394 and not w19395;
w19397 <= not w19098 and not w19351;
w19398 <= w19396 and w19397;
w19399 <= not w19396 and not w19397;
w19400 <= not w19398 and not w19399;
w19401 <= b(59) and w1791;
w19402 <= b(57) and w1941;
w19403 <= b(58) and w1786;
w19404 <= not w19402 and not w19403;
w19405 <= not w19401 and w19404;
w19406 <= w1794 and w11922;
w19407 <= w19405 and not w19406;
w19408 <= a(23) and not w19407;
w19409 <= a(23) and not w19408;
w19410 <= not w19407 and not w19408;
w19411 <= not w19409 and not w19410;
w19412 <= not w19114 and not w19348;
w19413 <= not w19411 and not w19412;
w19414 <= not w19411 and not w19413;
w19415 <= not w19412 and not w19413;
w19416 <= not w19414 and not w19415;
w19417 <= b(56) and w2282;
w19418 <= b(54) and w2428;
w19419 <= b(55) and w2277;
w19420 <= not w19418 and not w19419;
w19421 <= not w19417 and w19420;
w19422 <= w2285 and w10451;
w19423 <= w19421 and not w19422;
w19424 <= a(26) and not w19423;
w19425 <= a(26) and not w19424;
w19426 <= not w19423 and not w19424;
w19427 <= not w19425 and not w19426;
w19428 <= not w19128 and not w19343;
w19429 <= w19427 and w19428;
w19430 <= not w19427 and not w19428;
w19431 <= not w19429 and not w19430;
w19432 <= b(53) and w2793;
w19433 <= b(51) and w2986;
w19434 <= b(52) and w2788;
w19435 <= not w19433 and not w19434;
w19436 <= not w19432 and w19435;
w19437 <= w2796 and w9715;
w19438 <= w19436 and not w19437;
w19439 <= a(29) and not w19438;
w19440 <= a(29) and not w19439;
w19441 <= not w19438 and not w19439;
w19442 <= not w19440 and not w19441;
w19443 <= not w19145 and not w19340;
w19444 <= not w19442 and not w19443;
w19445 <= not w19442 and not w19444;
w19446 <= not w19443 and not w19444;
w19447 <= not w19445 and not w19446;
w19448 <= b(50) and w3381;
w19449 <= b(48) and w3586;
w19450 <= b(49) and w3376;
w19451 <= not w19449 and not w19450;
w19452 <= not w19448 and w19451;
w19453 <= w3384 and w8692;
w19454 <= w19452 and not w19453;
w19455 <= a(32) and not w19454;
w19456 <= a(32) and not w19455;
w19457 <= not w19454 and not w19455;
w19458 <= not w19456 and not w19457;
w19459 <= not w19323 and not w19336;
w19460 <= w19458 and w19459;
w19461 <= not w19458 and not w19459;
w19462 <= not w19460 and not w19461;
w19463 <= not w19314 and not w19317;
w19464 <= b(44) and w4778;
w19465 <= b(42) and w5020;
w19466 <= b(43) and w4773;
w19467 <= not w19465 and not w19466;
w19468 <= not w19464 and w19467;
w19469 <= w4781 and w6815;
w19470 <= w19468 and not w19469;
w19471 <= a(38) and not w19470;
w19472 <= a(38) and not w19471;
w19473 <= not w19470 and not w19471;
w19474 <= not w19472 and not w19473;
w19475 <= not w19306 and not w19310;
w19476 <= b(41) and w5520;
w19477 <= b(39) and w5802;
w19478 <= b(40) and w5515;
w19479 <= not w19477 and not w19478;
w19480 <= not w19476 and w19479;
w19481 <= w5523 and w5962;
w19482 <= w19480 and not w19481;
w19483 <= a(41) and not w19482;
w19484 <= a(41) and not w19483;
w19485 <= not w19482 and not w19483;
w19486 <= not w19484 and not w19485;
w19487 <= not w19298 and not w19302;
w19488 <= not w19238 and not w19251;
w19489 <= b(26) and w10169;
w19490 <= b(24) and w10539;
w19491 <= b(25) and w10164;
w19492 <= not w19490 and not w19491;
w19493 <= not w19489 and w19492;
w19494 <= w2556 and w10172;
w19495 <= w19493 and not w19494;
w19496 <= a(56) and not w19495;
w19497 <= a(56) and not w19496;
w19498 <= not w19495 and not w19496;
w19499 <= not w19497 and not w19498;
w19500 <= not w19218 and not w19232;
w19501 <= b(20) and w12411;
w19502 <= b(18) and w12790;
w19503 <= b(19) and w12406;
w19504 <= not w19502 and not w19503;
w19505 <= not w19501 and w19504;
w19506 <= w1589 and w12414;
w19507 <= w19505 and not w19506;
w19508 <= a(62) and not w19507;
w19509 <= a(62) and not w19508;
w19510 <= not w19507 and not w19508;
w19511 <= not w19509 and not w19510;
w19512 <= b(16) and w13646;
w19513 <= b(17) and not w13231;
w19514 <= not w19512 and not w19513;
w19515 <= w19199 and not w19514;
w19516 <= not w19199 and w19514;
w19517 <= not w19511 and not w19516;
w19518 <= not w19515 and w19517;
w19519 <= not w19511 and not w19518;
w19520 <= not w19516 and not w19518;
w19521 <= not w19515 and w19520;
w19522 <= not w19519 and not w19521;
w19523 <= not w19202 and not w19215;
w19524 <= w19522 and w19523;
w19525 <= not w19522 and not w19523;
w19526 <= not w19524 and not w19525;
w19527 <= b(23) and w11274;
w19528 <= b(21) and w11639;
w19529 <= b(22) and w11269;
w19530 <= not w19528 and not w19529;
w19531 <= not w19527 and w19530;
w19532 <= w2043 and w11277;
w19533 <= w19531 and not w19532;
w19534 <= a(59) and not w19533;
w19535 <= a(59) and not w19534;
w19536 <= not w19533 and not w19534;
w19537 <= not w19535 and not w19536;
w19538 <= not w19526 and w19537;
w19539 <= w19526 and not w19537;
w19540 <= not w19538 and not w19539;
w19541 <= not w19500 and w19540;
w19542 <= w19500 and not w19540;
w19543 <= not w19541 and not w19542;
w19544 <= not w19499 and w19543;
w19545 <= w19499 and not w19543;
w19546 <= not w19544 and not w19545;
w19547 <= not w19488 and w19546;
w19548 <= w19488 and not w19546;
w19549 <= not w19547 and not w19548;
w19550 <= b(29) and w9082;
w19551 <= b(27) and w9475;
w19552 <= b(28) and w9077;
w19553 <= not w19551 and not w19552;
w19554 <= not w19550 and w19553;
w19555 <= w3126 and w9085;
w19556 <= w19554 and not w19555;
w19557 <= a(53) and not w19556;
w19558 <= a(53) and not w19557;
w19559 <= not w19556 and not w19557;
w19560 <= not w19558 and not w19559;
w19561 <= w19549 and not w19560;
w19562 <= w19549 and not w19561;
w19563 <= not w19560 and not w19561;
w19564 <= not w19562 and not w19563;
w19565 <= not w18879 and not w19254;
w19566 <= not w19270 and not w19565;
w19567 <= not w19564 and not w19566;
w19568 <= not w19564 and not w19567;
w19569 <= not w19566 and not w19567;
w19570 <= not w19568 and not w19569;
w19571 <= b(32) and w8105;
w19572 <= b(30) and w8458;
w19573 <= b(31) and w8100;
w19574 <= not w19572 and not w19573;
w19575 <= not w19571 and w19574;
w19576 <= w3756 and w8108;
w19577 <= w19575 and not w19576;
w19578 <= a(50) and not w19577;
w19579 <= a(50) and not w19578;
w19580 <= not w19577 and not w19578;
w19581 <= not w19579 and not w19580;
w19582 <= not w19570 and w19581;
w19583 <= w19570 and not w19581;
w19584 <= not w19582 and not w19583;
w19585 <= not w19273 and not w19276;
w19586 <= w19584 and w19585;
w19587 <= not w19584 and not w19585;
w19588 <= not w19586 and not w19587;
w19589 <= b(35) and w7189;
w19590 <= b(33) and w7530;
w19591 <= b(34) and w7184;
w19592 <= not w19590 and not w19591;
w19593 <= not w19589 and w19592;
w19594 <= w4439 and w7192;
w19595 <= w19593 and not w19594;
w19596 <= a(47) and not w19595;
w19597 <= a(47) and not w19596;
w19598 <= not w19595 and not w19596;
w19599 <= not w19597 and not w19598;
w19600 <= w19588 and not w19599;
w19601 <= w19588 and not w19600;
w19602 <= not w19599 and not w19600;
w19603 <= not w19601 and not w19602;
w19604 <= not w19282 and not w19296;
w19605 <= not w19603 and not w19604;
w19606 <= not w19603 and not w19605;
w19607 <= not w19604 and not w19605;
w19608 <= not w19606 and not w19607;
w19609 <= b(38) and w6338;
w19610 <= b(36) and w6645;
w19611 <= b(37) and w6333;
w19612 <= not w19610 and not w19611;
w19613 <= not w19609 and w19612;
w19614 <= w4948 and w6341;
w19615 <= w19613 and not w19614;
w19616 <= a(44) and not w19615;
w19617 <= a(44) and not w19616;
w19618 <= not w19615 and not w19616;
w19619 <= not w19617 and not w19618;
w19620 <= not w19608 and w19619;
w19621 <= w19608 and not w19619;
w19622 <= not w19620 and not w19621;
w19623 <= not w19487 and not w19622;
w19624 <= w19487 and w19622;
w19625 <= not w19623 and not w19624;
w19626 <= not w19486 and w19625;
w19627 <= w19486 and not w19625;
w19628 <= not w19626 and not w19627;
w19629 <= not w19475 and w19628;
w19630 <= w19475 and not w19628;
w19631 <= not w19629 and not w19630;
w19632 <= not w19474 and w19631;
w19633 <= w19474 and not w19631;
w19634 <= not w19632 and not w19633;
w19635 <= not w19463 and w19634;
w19636 <= w19463 and not w19634;
w19637 <= not w19635 and not w19636;
w19638 <= b(47) and w4030;
w19639 <= b(45) and w4275;
w19640 <= b(46) and w4025;
w19641 <= not w19639 and not w19640;
w19642 <= not w19638 and w19641;
w19643 <= w4033 and w7446;
w19644 <= w19642 and not w19643;
w19645 <= a(35) and not w19644;
w19646 <= a(35) and not w19645;
w19647 <= not w19644 and not w19645;
w19648 <= not w19646 and not w19647;
w19649 <= w19637 and not w19648;
w19650 <= w19637 and not w19649;
w19651 <= not w19648 and not w19649;
w19652 <= not w19650 and not w19651;
w19653 <= w19462 and not w19652;
w19654 <= not w19462 and w19652;
w19655 <= not w19447 and not w19654;
w19656 <= not w19653 and w19655;
w19657 <= not w19447 and not w19656;
w19658 <= not w19654 and not w19656;
w19659 <= not w19653 and w19658;
w19660 <= not w19657 and not w19659;
w19661 <= w19431 and not w19660;
w19662 <= not w19431 and w19660;
w19663 <= not w19416 and not w19662;
w19664 <= not w19661 and w19663;
w19665 <= not w19416 and not w19664;
w19666 <= not w19662 and not w19664;
w19667 <= not w19661 and w19666;
w19668 <= not w19665 and not w19667;
w19669 <= not w19400 and w19668;
w19670 <= w19400 and not w19668;
w19671 <= not w19669 and not w19670;
w19672 <= not w19385 and w19671;
w19673 <= w19385 and not w19671;
w19674 <= not w19672 and not w19673;
w19675 <= not w19373 and w19674;
w19676 <= not w19373 and not w19675;
w19677 <= w19674 and not w19675;
w19678 <= not w19676 and not w19677;
w19679 <= not w19372 and not w19678;
w19680 <= w19372 and not w19677;
w19681 <= not w19676 and w19680;
w19682 <= not w19679 and not w19681;
w19683 <= not w19675 and not w19679;
w19684 <= not w19382 and not w19672;
w19685 <= not w19399 and not w19670;
w19686 <= b(63) and w1370;
w19687 <= b(61) and w1506;
w19688 <= b(62) and w1365;
w19689 <= not w19687 and not w19688;
w19690 <= not w19686 and w19689;
w19691 <= w1373 and w13514;
w19692 <= w19690 and not w19691;
w19693 <= a(20) and not w19692;
w19694 <= a(20) and not w19693;
w19695 <= not w19692 and not w19693;
w19696 <= not w19694 and not w19695;
w19697 <= not w19685 and not w19696;
w19698 <= not w19685 and not w19697;
w19699 <= not w19696 and not w19697;
w19700 <= not w19698 and not w19699;
w19701 <= b(60) and w1791;
w19702 <= b(58) and w1941;
w19703 <= b(59) and w1786;
w19704 <= not w19702 and not w19703;
w19705 <= not w19701 and w19704;
w19706 <= w1794 and w11954;
w19707 <= w19705 and not w19706;
w19708 <= a(23) and not w19707;
w19709 <= a(23) and not w19708;
w19710 <= not w19707 and not w19708;
w19711 <= not w19709 and not w19710;
w19712 <= not w19413 and not w19664;
w19713 <= w19711 and w19712;
w19714 <= not w19711 and not w19712;
w19715 <= not w19713 and not w19714;
w19716 <= b(54) and w2793;
w19717 <= b(52) and w2986;
w19718 <= b(53) and w2788;
w19719 <= not w19717 and not w19718;
w19720 <= not w19716 and w19719;
w19721 <= w2796 and w9741;
w19722 <= w19720 and not w19721;
w19723 <= a(29) and not w19722;
w19724 <= a(29) and not w19723;
w19725 <= not w19722 and not w19723;
w19726 <= not w19724 and not w19725;
w19727 <= not w19444 and not w19656;
w19728 <= w19726 and w19727;
w19729 <= not w19726 and not w19727;
w19730 <= not w19728 and not w19729;
w19731 <= not w19623 and not w19626;
w19732 <= not w19608 and not w19619;
w19733 <= not w19605 and not w19732;
w19734 <= not w19587 and not w19600;
w19735 <= b(27) and w10169;
w19736 <= b(25) and w10539;
w19737 <= b(26) and w10164;
w19738 <= not w19736 and not w19737;
w19739 <= not w19735 and w19738;
w19740 <= w2733 and w10172;
w19741 <= w19739 and not w19740;
w19742 <= a(56) and not w19741;
w19743 <= a(56) and not w19742;
w19744 <= not w19741 and not w19742;
w19745 <= not w19743 and not w19744;
w19746 <= not w19525 and not w19539;
w19747 <= b(21) and w12411;
w19748 <= b(19) and w12790;
w19749 <= b(20) and w12406;
w19750 <= not w19748 and not w19749;
w19751 <= not w19747 and w19750;
w19752 <= w1727 and w12414;
w19753 <= w19751 and not w19752;
w19754 <= a(62) and not w19753;
w19755 <= a(62) and not w19754;
w19756 <= not w19753 and not w19754;
w19757 <= not w19755 and not w19756;
w19758 <= b(17) and w13646;
w19759 <= b(18) and not w13231;
w19760 <= not w19758 and not w19759;
w19761 <= not a(17) and not w19760;
w19762 <= a(17) and w19760;
w19763 <= not w19761 and not w19762;
w19764 <= not w19514 and w19763;
w19765 <= w19514 and not w19763;
w19766 <= not w19764 and not w19765;
w19767 <= not w19757 and w19766;
w19768 <= not w19757 and not w19767;
w19769 <= w19766 and not w19767;
w19770 <= not w19768 and not w19769;
w19771 <= not w19520 and not w19770;
w19772 <= not w19520 and not w19771;
w19773 <= not w19770 and not w19771;
w19774 <= not w19772 and not w19773;
w19775 <= b(24) and w11274;
w19776 <= b(22) and w11639;
w19777 <= b(23) and w11269;
w19778 <= not w19776 and not w19777;
w19779 <= not w19775 and w19778;
w19780 <= w2201 and w11277;
w19781 <= w19779 and not w19780;
w19782 <= a(59) and not w19781;
w19783 <= a(59) and not w19782;
w19784 <= not w19781 and not w19782;
w19785 <= not w19783 and not w19784;
w19786 <= w19774 and w19785;
w19787 <= not w19774 and not w19785;
w19788 <= not w19786 and not w19787;
w19789 <= not w19746 and w19788;
w19790 <= w19746 and not w19788;
w19791 <= not w19789 and not w19790;
w19792 <= not w19745 and w19791;
w19793 <= w19791 and not w19792;
w19794 <= not w19745 and not w19792;
w19795 <= not w19793 and not w19794;
w19796 <= not w19541 and not w19544;
w19797 <= w19795 and w19796;
w19798 <= not w19795 and not w19796;
w19799 <= not w19797 and not w19798;
w19800 <= b(30) and w9082;
w19801 <= b(28) and w9475;
w19802 <= b(29) and w9077;
w19803 <= not w19801 and not w19802;
w19804 <= not w19800 and w19803;
w19805 <= w3320 and w9085;
w19806 <= w19804 and not w19805;
w19807 <= a(53) and not w19806;
w19808 <= a(53) and not w19807;
w19809 <= not w19806 and not w19807;
w19810 <= not w19808 and not w19809;
w19811 <= w19799 and not w19810;
w19812 <= w19799 and not w19811;
w19813 <= not w19810 and not w19811;
w19814 <= not w19812 and not w19813;
w19815 <= not w19547 and not w19561;
w19816 <= w19814 and w19815;
w19817 <= not w19814 and not w19815;
w19818 <= not w19816 and not w19817;
w19819 <= b(33) and w8105;
w19820 <= b(31) and w8458;
w19821 <= b(32) and w8100;
w19822 <= not w19820 and not w19821;
w19823 <= not w19819 and w19822;
w19824 <= w3966 and w8108;
w19825 <= w19823 and not w19824;
w19826 <= a(50) and not w19825;
w19827 <= a(50) and not w19826;
w19828 <= not w19825 and not w19826;
w19829 <= not w19827 and not w19828;
w19830 <= not w19570 and not w19581;
w19831 <= not w19567 and not w19830;
w19832 <= not w19829 and not w19831;
w19833 <= w19829 and w19831;
w19834 <= not w19832 and not w19833;
w19835 <= not w19818 and w19834;
w19836 <= w19818 and not w19834;
w19837 <= not w19835 and not w19836;
w19838 <= b(36) and w7189;
w19839 <= b(34) and w7530;
w19840 <= b(35) and w7184;
w19841 <= not w19839 and not w19840;
w19842 <= not w19838 and w19841;
w19843 <= w4665 and w7192;
w19844 <= w19842 and not w19843;
w19845 <= a(47) and not w19844;
w19846 <= a(47) and not w19845;
w19847 <= not w19844 and not w19845;
w19848 <= not w19846 and not w19847;
w19849 <= not w19837 and not w19848;
w19850 <= w19837 and w19848;
w19851 <= not w19849 and not w19850;
w19852 <= w19734 and not w19851;
w19853 <= not w19734 and w19851;
w19854 <= not w19852 and not w19853;
w19855 <= b(39) and w6338;
w19856 <= b(37) and w6645;
w19857 <= b(38) and w6333;
w19858 <= not w19856 and not w19857;
w19859 <= not w19855 and w19858;
w19860 <= w5194 and w6341;
w19861 <= w19859 and not w19860;
w19862 <= a(44) and not w19861;
w19863 <= a(44) and not w19862;
w19864 <= not w19861 and not w19862;
w19865 <= not w19863 and not w19864;
w19866 <= w19854 and not w19865;
w19867 <= w19854 and not w19866;
w19868 <= not w19865 and not w19866;
w19869 <= not w19867 and not w19868;
w19870 <= not w19733 and w19869;
w19871 <= w19733 and not w19869;
w19872 <= not w19870 and not w19871;
w19873 <= b(42) and w5520;
w19874 <= b(40) and w5802;
w19875 <= b(41) and w5515;
w19876 <= not w19874 and not w19875;
w19877 <= not w19873 and w19876;
w19878 <= w5523 and w6232;
w19879 <= w19877 and not w19878;
w19880 <= a(41) and not w19879;
w19881 <= a(41) and not w19880;
w19882 <= not w19879 and not w19880;
w19883 <= not w19881 and not w19882;
w19884 <= not w19872 and not w19883;
w19885 <= w19872 and w19883;
w19886 <= not w19884 and not w19885;
w19887 <= w19731 and not w19886;
w19888 <= not w19731 and w19886;
w19889 <= not w19887 and not w19888;
w19890 <= b(45) and w4778;
w19891 <= b(43) and w5020;
w19892 <= b(44) and w4773;
w19893 <= not w19891 and not w19892;
w19894 <= not w19890 and w19893;
w19895 <= w4781 and w7104;
w19896 <= w19894 and not w19895;
w19897 <= a(38) and not w19896;
w19898 <= a(38) and not w19897;
w19899 <= not w19896 and not w19897;
w19900 <= not w19898 and not w19899;
w19901 <= w19889 and not w19900;
w19902 <= w19889 and not w19901;
w19903 <= not w19900 and not w19901;
w19904 <= not w19902 and not w19903;
w19905 <= not w19629 and not w19632;
w19906 <= w19904 and w19905;
w19907 <= not w19904 and not w19905;
w19908 <= not w19906 and not w19907;
w19909 <= b(48) and w4030;
w19910 <= b(46) and w4275;
w19911 <= b(47) and w4025;
w19912 <= not w19910 and not w19911;
w19913 <= not w19909 and w19912;
w19914 <= w4033 and w7752;
w19915 <= w19913 and not w19914;
w19916 <= a(35) and not w19915;
w19917 <= a(35) and not w19916;
w19918 <= not w19915 and not w19916;
w19919 <= not w19917 and not w19918;
w19920 <= w19908 and not w19919;
w19921 <= w19908 and not w19920;
w19922 <= not w19919 and not w19920;
w19923 <= not w19921 and not w19922;
w19924 <= not w19635 and not w19649;
w19925 <= w19923 and w19924;
w19926 <= not w19923 and not w19924;
w19927 <= not w19925 and not w19926;
w19928 <= b(51) and w3381;
w19929 <= b(49) and w3586;
w19930 <= b(50) and w3376;
w19931 <= not w19929 and not w19930;
w19932 <= not w19928 and w19931;
w19933 <= w3384 and w8719;
w19934 <= w19932 and not w19933;
w19935 <= a(32) and not w19934;
w19936 <= a(32) and not w19935;
w19937 <= not w19934 and not w19935;
w19938 <= not w19936 and not w19937;
w19939 <= not w19461 and not w19653;
w19940 <= not w19938 and not w19939;
w19941 <= w19938 and w19939;
w19942 <= not w19940 and not w19941;
w19943 <= w19927 and w19942;
w19944 <= w19927 and not w19943;
w19945 <= w19942 and not w19943;
w19946 <= not w19944 and not w19945;
w19947 <= w19730 and not w19946;
w19948 <= w19730 and not w19947;
w19949 <= not w19946 and not w19947;
w19950 <= not w19948 and not w19949;
w19951 <= b(57) and w2282;
w19952 <= b(55) and w2428;
w19953 <= b(56) and w2277;
w19954 <= not w19952 and not w19953;
w19955 <= not w19951 and w19954;
w19956 <= w2285 and w11153;
w19957 <= w19955 and not w19956;
w19958 <= a(26) and not w19957;
w19959 <= a(26) and not w19958;
w19960 <= not w19957 and not w19958;
w19961 <= not w19959 and not w19960;
w19962 <= not w19430 and not w19661;
w19963 <= not w19961 and not w19962;
w19964 <= w19961 and w19962;
w19965 <= not w19963 and not w19964;
w19966 <= not w19950 and w19965;
w19967 <= not w19950 and not w19966;
w19968 <= w19965 and not w19966;
w19969 <= not w19967 and not w19968;
w19970 <= w19715 and not w19969;
w19971 <= w19715 and not w19970;
w19972 <= not w19969 and not w19970;
w19973 <= not w19971 and not w19972;
w19974 <= not w19700 and w19973;
w19975 <= w19700 and not w19973;
w19976 <= not w19974 and not w19975;
w19977 <= not w19684 and not w19976;
w19978 <= not w19684 and not w19977;
w19979 <= not w19976 and not w19977;
w19980 <= not w19978 and not w19979;
w19981 <= not w19683 and not w19980;
w19982 <= w19683 and not w19979;
w19983 <= not w19978 and w19982;
w19984 <= not w19981 and not w19983;
w19985 <= not w19977 and not w19981;
w19986 <= not w19700 and not w19973;
w19987 <= not w19697 and not w19986;
w19988 <= b(61) and w1791;
w19989 <= b(59) and w1941;
w19990 <= b(60) and w1786;
w19991 <= not w19989 and not w19990;
w19992 <= not w19988 and w19991;
w19993 <= w1794 and w12712;
w19994 <= w19992 and not w19993;
w19995 <= a(23) and not w19994;
w19996 <= a(23) and not w19995;
w19997 <= not w19994 and not w19995;
w19998 <= not w19996 and not w19997;
w19999 <= not w19963 and not w19966;
w20000 <= w19998 and w19999;
w20001 <= not w19998 and not w19999;
w20002 <= not w20000 and not w20001;
w20003 <= b(58) and w2282;
w20004 <= b(56) and w2428;
w20005 <= b(57) and w2277;
w20006 <= not w20004 and not w20005;
w20007 <= not w20003 and w20006;
w20008 <= w2285 and w11179;
w20009 <= w20007 and not w20008;
w20010 <= a(26) and not w20009;
w20011 <= a(26) and not w20010;
w20012 <= not w20009 and not w20010;
w20013 <= not w20011 and not w20012;
w20014 <= not w19729 and not w19947;
w20015 <= w20013 and w20014;
w20016 <= not w20013 and not w20014;
w20017 <= not w20015 and not w20016;
w20018 <= b(55) and w2793;
w20019 <= b(53) and w2986;
w20020 <= b(54) and w2788;
w20021 <= not w20019 and not w20020;
w20022 <= not w20018 and w20021;
w20023 <= w2796 and w10427;
w20024 <= w20022 and not w20023;
w20025 <= a(29) and not w20024;
w20026 <= a(29) and not w20025;
w20027 <= not w20024 and not w20025;
w20028 <= not w20026 and not w20027;
w20029 <= not w19940 and not w19943;
w20030 <= w20028 and w20029;
w20031 <= not w20028 and not w20029;
w20032 <= not w20030 and not w20031;
w20033 <= b(52) and w3381;
w20034 <= b(50) and w3586;
w20035 <= b(51) and w3376;
w20036 <= not w20034 and not w20035;
w20037 <= not w20033 and w20036;
w20038 <= w3384 and w9371;
w20039 <= w20037 and not w20038;
w20040 <= a(32) and not w20039;
w20041 <= a(32) and not w20040;
w20042 <= not w20039 and not w20040;
w20043 <= not w20041 and not w20042;
w20044 <= not w19920 and not w19926;
w20045 <= w20043 and w20044;
w20046 <= not w20043 and not w20044;
w20047 <= not w20045 and not w20046;
w20048 <= b(43) and w5520;
w20049 <= b(41) and w5802;
w20050 <= b(42) and w5515;
w20051 <= not w20049 and not w20050;
w20052 <= not w20048 and w20051;
w20053 <= w5523 and w6258;
w20054 <= w20052 and not w20053;
w20055 <= a(41) and not w20054;
w20056 <= a(41) and not w20055;
w20057 <= not w20054 and not w20055;
w20058 <= not w20056 and not w20057;
w20059 <= not w19733 and not w19869;
w20060 <= not w19866 and not w20059;
w20061 <= b(40) and w6338;
w20062 <= b(38) and w6645;
w20063 <= b(39) and w6333;
w20064 <= not w20062 and not w20063;
w20065 <= not w20061 and w20064;
w20066 <= w5698 and w6341;
w20067 <= w20065 and not w20066;
w20068 <= a(44) and not w20067;
w20069 <= a(44) and not w20068;
w20070 <= not w20067 and not w20068;
w20071 <= not w20069 and not w20070;
w20072 <= not w19849 and not w19853;
w20073 <= b(31) and w9082;
w20074 <= b(29) and w9475;
w20075 <= b(30) and w9077;
w20076 <= not w20074 and not w20075;
w20077 <= not w20073 and w20076;
w20078 <= w3539 and w9085;
w20079 <= w20077 and not w20078;
w20080 <= a(53) and not w20079;
w20081 <= a(53) and not w20080;
w20082 <= not w20079 and not w20080;
w20083 <= not w20081 and not w20082;
w20084 <= not w19787 and not w19789;
w20085 <= b(25) and w11274;
w20086 <= b(23) and w11639;
w20087 <= b(24) and w11269;
w20088 <= not w20086 and not w20087;
w20089 <= not w20085 and w20088;
w20090 <= w2228 and w11277;
w20091 <= w20089 and not w20090;
w20092 <= a(59) and not w20091;
w20093 <= a(59) and not w20092;
w20094 <= not w20091 and not w20092;
w20095 <= not w20093 and not w20094;
w20096 <= b(18) and w13646;
w20097 <= b(19) and not w13231;
w20098 <= not w20096 and not w20097;
w20099 <= not w19761 and not w19764;
w20100 <= not w20098 and w20099;
w20101 <= w20098 and not w20099;
w20102 <= not w20100 and not w20101;
w20103 <= b(22) and w12411;
w20104 <= b(20) and w12790;
w20105 <= b(21) and w12406;
w20106 <= not w20104 and not w20105;
w20107 <= not w20103 and w20106;
w20108 <= w1888 and w12414;
w20109 <= w20107 and not w20108;
w20110 <= a(62) and not w20109;
w20111 <= a(62) and not w20110;
w20112 <= not w20109 and not w20110;
w20113 <= not w20111 and not w20112;
w20114 <= not w20102 and w20113;
w20115 <= w20102 and not w20113;
w20116 <= not w20114 and not w20115;
w20117 <= not w19767 and not w19771;
w20118 <= w20116 and not w20117;
w20119 <= not w20116 and w20117;
w20120 <= not w20118 and not w20119;
w20121 <= not w20095 and w20120;
w20122 <= w20120 and not w20121;
w20123 <= not w20095 and not w20121;
w20124 <= not w20122 and not w20123;
w20125 <= not w20084 and w20124;
w20126 <= w20084 and not w20124;
w20127 <= not w20125 and not w20126;
w20128 <= b(28) and w10169;
w20129 <= b(26) and w10539;
w20130 <= b(27) and w10164;
w20131 <= not w20129 and not w20130;
w20132 <= not w20128 and w20131;
w20133 <= w2932 and w10172;
w20134 <= w20132 and not w20133;
w20135 <= a(56) and not w20134;
w20136 <= a(56) and not w20135;
w20137 <= not w20134 and not w20135;
w20138 <= not w20136 and not w20137;
w20139 <= w20127 and w20138;
w20140 <= not w20127 and not w20138;
w20141 <= not w20139 and not w20140;
w20142 <= not w19792 and not w19798;
w20143 <= w20141 and not w20142;
w20144 <= not w20141 and w20142;
w20145 <= not w20143 and not w20144;
w20146 <= not w20083 and w20145;
w20147 <= w20145 and not w20146;
w20148 <= not w20083 and not w20146;
w20149 <= not w20147 and not w20148;
w20150 <= not w19811 and not w19817;
w20151 <= w20149 and w20150;
w20152 <= not w20149 and not w20150;
w20153 <= not w20151 and not w20152;
w20154 <= b(34) and w8105;
w20155 <= b(32) and w8458;
w20156 <= b(33) and w8100;
w20157 <= not w20155 and not w20156;
w20158 <= not w20154 and w20157;
w20159 <= w4209 and w8108;
w20160 <= w20158 and not w20159;
w20161 <= a(50) and not w20160;
w20162 <= a(50) and not w20161;
w20163 <= not w20160 and not w20161;
w20164 <= not w20162 and not w20163;
w20165 <= w20153 and not w20164;
w20166 <= w20153 and not w20165;
w20167 <= not w20164 and not w20165;
w20168 <= not w20166 and not w20167;
w20169 <= w19818 and w19834;
w20170 <= not w19832 and not w20169;
w20171 <= w20168 and w20170;
w20172 <= not w20168 and not w20170;
w20173 <= not w20171 and not w20172;
w20174 <= b(37) and w7189;
w20175 <= b(35) and w7530;
w20176 <= b(36) and w7184;
w20177 <= not w20175 and not w20176;
w20178 <= not w20174 and w20177;
w20179 <= w4924 and w7192;
w20180 <= w20178 and not w20179;
w20181 <= a(47) and not w20180;
w20182 <= a(47) and not w20181;
w20183 <= not w20180 and not w20181;
w20184 <= not w20182 and not w20183;
w20185 <= not w20173 and w20184;
w20186 <= w20173 and not w20184;
w20187 <= not w20185 and not w20186;
w20188 <= not w20072 and w20187;
w20189 <= not w20072 and not w20188;
w20190 <= w20187 and not w20188;
w20191 <= not w20189 and not w20190;
w20192 <= not w20071 and not w20191;
w20193 <= w20071 and not w20190;
w20194 <= not w20189 and w20193;
w20195 <= not w20192 and not w20194;
w20196 <= not w20060 and w20195;
w20197 <= w20060 and not w20195;
w20198 <= not w20196 and not w20197;
w20199 <= not w20058 and w20198;
w20200 <= w20198 and not w20199;
w20201 <= not w20058 and not w20199;
w20202 <= not w20200 and not w20201;
w20203 <= not w19884 and not w19888;
w20204 <= w20202 and w20203;
w20205 <= not w20202 and not w20203;
w20206 <= not w20204 and not w20205;
w20207 <= b(46) and w4778;
w20208 <= b(44) and w5020;
w20209 <= b(45) and w4773;
w20210 <= not w20208 and not w20209;
w20211 <= not w20207 and w20210;
w20212 <= w4781 and w7420;
w20213 <= w20211 and not w20212;
w20214 <= a(38) and not w20213;
w20215 <= a(38) and not w20214;
w20216 <= not w20213 and not w20214;
w20217 <= not w20215 and not w20216;
w20218 <= w20206 and not w20217;
w20219 <= w20206 and not w20218;
w20220 <= not w20217 and not w20218;
w20221 <= not w20219 and not w20220;
w20222 <= not w19901 and not w19907;
w20223 <= w20221 and w20222;
w20224 <= not w20221 and not w20222;
w20225 <= not w20223 and not w20224;
w20226 <= b(49) and w4030;
w20227 <= b(47) and w4275;
w20228 <= b(48) and w4025;
w20229 <= not w20227 and not w20228;
w20230 <= not w20226 and w20229;
w20231 <= w4033 and w8368;
w20232 <= w20230 and not w20231;
w20233 <= a(35) and not w20232;
w20234 <= a(35) and not w20233;
w20235 <= not w20232 and not w20233;
w20236 <= not w20234 and not w20235;
w20237 <= w20225 and not w20236;
w20238 <= w20225 and not w20237;
w20239 <= not w20236 and not w20237;
w20240 <= not w20238 and not w20239;
w20241 <= w20047 and not w20240;
w20242 <= not w20047 and w20240;
w20243 <= w20032 and not w20242;
w20244 <= not w20241 and w20243;
w20245 <= w20032 and not w20244;
w20246 <= not w20242 and not w20244;
w20247 <= not w20241 and w20246;
w20248 <= not w20245 and not w20247;
w20249 <= w20017 and not w20248;
w20250 <= not w20017 and w20248;
w20251 <= w20002 and not w20250;
w20252 <= not w20249 and w20251;
w20253 <= w20002 and not w20252;
w20254 <= not w20250 and not w20252;
w20255 <= not w20249 and w20254;
w20256 <= not w20253 and not w20255;
w20257 <= not w19714 and not w19970;
w20258 <= b(62) and w1506;
w20259 <= b(63) and w1365;
w20260 <= not w20258 and not w20259;
w20261 <= not w1373 and w20260;
w20262 <= w13543 and w20260;
w20263 <= not w20261 and not w20262;
w20264 <= a(20) and not w20263;
w20265 <= not a(20) and w20263;
w20266 <= not w20264 and not w20265;
w20267 <= not w20257 and not w20266;
w20268 <= not w20257 and not w20267;
w20269 <= not w20266 and not w20267;
w20270 <= not w20268 and not w20269;
w20271 <= not w20256 and not w20270;
w20272 <= w20256 and not w20269;
w20273 <= not w20268 and w20272;
w20274 <= not w20271 and not w20273;
w20275 <= not w19987 and w20274;
w20276 <= not w19987 and not w20275;
w20277 <= w20274 and not w20275;
w20278 <= not w20276 and not w20277;
w20279 <= not w19985 and not w20278;
w20280 <= w19985 and not w20277;
w20281 <= not w20276 and w20280;
w20282 <= not w20279 and not w20281;
w20283 <= not w20275 and not w20279;
w20284 <= not w20267 and not w20271;
w20285 <= not w20001 and not w20252;
w20286 <= b(63) and w1506;
w20287 <= w1373 and w13540;
w20288 <= not w20286 and not w20287;
w20289 <= a(20) and not w20288;
w20290 <= a(20) and not w20289;
w20291 <= not w20288 and not w20289;
w20292 <= not w20290 and not w20291;
w20293 <= not w20285 and not w20292;
w20294 <= not w20285 and not w20293;
w20295 <= not w20292 and not w20293;
w20296 <= not w20294 and not w20295;
w20297 <= b(62) and w1791;
w20298 <= b(60) and w1941;
w20299 <= b(61) and w1786;
w20300 <= not w20298 and not w20299;
w20301 <= not w20297 and w20300;
w20302 <= w1794 and w13113;
w20303 <= w20301 and not w20302;
w20304 <= a(23) and not w20303;
w20305 <= a(23) and not w20304;
w20306 <= not w20303 and not w20304;
w20307 <= not w20305 and not w20306;
w20308 <= not w20016 and not w20249;
w20309 <= not w20307 and not w20308;
w20310 <= not w20307 and not w20309;
w20311 <= not w20308 and not w20309;
w20312 <= not w20310 and not w20311;
w20313 <= b(59) and w2282;
w20314 <= b(57) and w2428;
w20315 <= b(58) and w2277;
w20316 <= not w20314 and not w20315;
w20317 <= not w20313 and w20316;
w20318 <= w2285 and w11922;
w20319 <= w20317 and not w20318;
w20320 <= a(26) and not w20319;
w20321 <= a(26) and not w20320;
w20322 <= not w20319 and not w20320;
w20323 <= not w20321 and not w20322;
w20324 <= not w20031 and not w20244;
w20325 <= w20323 and w20324;
w20326 <= not w20323 and not w20324;
w20327 <= not w20325 and not w20326;
w20328 <= b(56) and w2793;
w20329 <= b(54) and w2986;
w20330 <= b(55) and w2788;
w20331 <= not w20329 and not w20330;
w20332 <= not w20328 and w20331;
w20333 <= w2796 and w10451;
w20334 <= w20332 and not w20333;
w20335 <= a(29) and not w20334;
w20336 <= a(29) and not w20335;
w20337 <= not w20334 and not w20335;
w20338 <= not w20336 and not w20337;
w20339 <= not w20046 and not w20241;
w20340 <= not w20338 and not w20339;
w20341 <= not w20338 and not w20340;
w20342 <= not w20339 and not w20340;
w20343 <= not w20341 and not w20342;
w20344 <= b(53) and w3381;
w20345 <= b(51) and w3586;
w20346 <= b(52) and w3376;
w20347 <= not w20345 and not w20346;
w20348 <= not w20344 and w20347;
w20349 <= w3384 and w9715;
w20350 <= w20348 and not w20349;
w20351 <= a(32) and not w20350;
w20352 <= a(32) and not w20351;
w20353 <= not w20350 and not w20351;
w20354 <= not w20352 and not w20353;
w20355 <= not w20224 and not w20237;
w20356 <= w20354 and w20355;
w20357 <= not w20354 and not w20355;
w20358 <= not w20356 and not w20357;
w20359 <= not w20196 and not w20199;
w20360 <= b(44) and w5520;
w20361 <= b(42) and w5802;
w20362 <= b(43) and w5515;
w20363 <= not w20361 and not w20362;
w20364 <= not w20360 and w20363;
w20365 <= w5523 and w6815;
w20366 <= w20364 and not w20365;
w20367 <= a(41) and not w20366;
w20368 <= a(41) and not w20367;
w20369 <= not w20366 and not w20367;
w20370 <= not w20368 and not w20369;
w20371 <= not w20188 and not w20192;
w20372 <= b(41) and w6338;
w20373 <= b(39) and w6645;
w20374 <= b(40) and w6333;
w20375 <= not w20373 and not w20374;
w20376 <= not w20372 and w20375;
w20377 <= w5962 and w6341;
w20378 <= w20376 and not w20377;
w20379 <= a(44) and not w20378;
w20380 <= a(44) and not w20379;
w20381 <= not w20378 and not w20379;
w20382 <= not w20380 and not w20381;
w20383 <= not w20172 and not w20186;
w20384 <= b(38) and w7189;
w20385 <= b(36) and w7530;
w20386 <= b(37) and w7184;
w20387 <= not w20385 and not w20386;
w20388 <= not w20384 and w20387;
w20389 <= w4948 and w7192;
w20390 <= w20388 and not w20389;
w20391 <= a(47) and not w20390;
w20392 <= a(47) and not w20391;
w20393 <= not w20390 and not w20391;
w20394 <= not w20392 and not w20393;
w20395 <= not w20152 and not w20165;
w20396 <= b(35) and w8105;
w20397 <= b(33) and w8458;
w20398 <= b(34) and w8100;
w20399 <= not w20397 and not w20398;
w20400 <= not w20396 and w20399;
w20401 <= w4439 and w8108;
w20402 <= w20400 and not w20401;
w20403 <= a(50) and not w20402;
w20404 <= a(50) and not w20403;
w20405 <= not w20402 and not w20403;
w20406 <= not w20404 and not w20405;
w20407 <= not w20143 and not w20146;
w20408 <= not w20118 and not w20121;
w20409 <= b(26) and w11274;
w20410 <= b(24) and w11639;
w20411 <= b(25) and w11269;
w20412 <= not w20410 and not w20411;
w20413 <= not w20409 and w20412;
w20414 <= w2556 and w11277;
w20415 <= w20413 and not w20414;
w20416 <= a(59) and not w20415;
w20417 <= a(59) and not w20416;
w20418 <= not w20415 and not w20416;
w20419 <= not w20417 and not w20418;
w20420 <= not w20101 and not w20115;
w20421 <= b(19) and w13646;
w20422 <= b(20) and not w13231;
w20423 <= not w20421 and not w20422;
w20424 <= not w20098 and w20423;
w20425 <= w20098 and not w20423;
w20426 <= not w20424 and not w20425;
w20427 <= b(23) and w12411;
w20428 <= b(21) and w12790;
w20429 <= b(22) and w12406;
w20430 <= not w20428 and not w20429;
w20431 <= not w20427 and w20430;
w20432 <= not w12414 and w20431;
w20433 <= not w2043 and w20431;
w20434 <= not w20432 and not w20433;
w20435 <= a(62) and not w20434;
w20436 <= not a(62) and w20434;
w20437 <= not w20435 and not w20436;
w20438 <= w20426 and not w20437;
w20439 <= not w20426 and w20437;
w20440 <= not w20438 and not w20439;
w20441 <= not w20420 and w20440;
w20442 <= w20420 and not w20440;
w20443 <= not w20441 and not w20442;
w20444 <= not w20419 and w20443;
w20445 <= w20419 and not w20443;
w20446 <= not w20444 and not w20445;
w20447 <= not w20408 and w20446;
w20448 <= w20408 and not w20446;
w20449 <= not w20447 and not w20448;
w20450 <= b(29) and w10169;
w20451 <= b(27) and w10539;
w20452 <= b(28) and w10164;
w20453 <= not w20451 and not w20452;
w20454 <= not w20450 and w20453;
w20455 <= w3126 and w10172;
w20456 <= w20454 and not w20455;
w20457 <= a(56) and not w20456;
w20458 <= a(56) and not w20457;
w20459 <= not w20456 and not w20457;
w20460 <= not w20458 and not w20459;
w20461 <= w20449 and not w20460;
w20462 <= w20449 and not w20461;
w20463 <= not w20460 and not w20461;
w20464 <= not w20462 and not w20463;
w20465 <= not w20084 and not w20124;
w20466 <= not w20140 and not w20465;
w20467 <= not w20464 and not w20466;
w20468 <= not w20464 and not w20467;
w20469 <= not w20466 and not w20467;
w20470 <= not w20468 and not w20469;
w20471 <= b(32) and w9082;
w20472 <= b(30) and w9475;
w20473 <= b(31) and w9077;
w20474 <= not w20472 and not w20473;
w20475 <= not w20471 and w20474;
w20476 <= w3756 and w9085;
w20477 <= w20475 and not w20476;
w20478 <= a(53) and not w20477;
w20479 <= a(53) and not w20478;
w20480 <= not w20477 and not w20478;
w20481 <= not w20479 and not w20480;
w20482 <= not w20470 and w20481;
w20483 <= w20470 and not w20481;
w20484 <= not w20482 and not w20483;
w20485 <= not w20407 and not w20484;
w20486 <= w20407 and w20484;
w20487 <= not w20485 and not w20486;
w20488 <= not w20406 and w20487;
w20489 <= w20406 and not w20487;
w20490 <= not w20488 and not w20489;
w20491 <= not w20395 and w20490;
w20492 <= w20395 and not w20490;
w20493 <= not w20491 and not w20492;
w20494 <= not w20394 and w20493;
w20495 <= w20394 and not w20493;
w20496 <= not w20494 and not w20495;
w20497 <= not w20383 and w20496;
w20498 <= w20383 and not w20496;
w20499 <= not w20497 and not w20498;
w20500 <= not w20382 and w20499;
w20501 <= w20382 and not w20499;
w20502 <= not w20500 and not w20501;
w20503 <= not w20371 and w20502;
w20504 <= w20371 and not w20502;
w20505 <= not w20503 and not w20504;
w20506 <= not w20370 and w20505;
w20507 <= w20370 and not w20505;
w20508 <= not w20506 and not w20507;
w20509 <= not w20359 and w20508;
w20510 <= w20359 and not w20508;
w20511 <= not w20509 and not w20510;
w20512 <= b(47) and w4778;
w20513 <= b(45) and w5020;
w20514 <= b(46) and w4773;
w20515 <= not w20513 and not w20514;
w20516 <= not w20512 and w20515;
w20517 <= w4781 and w7446;
w20518 <= w20516 and not w20517;
w20519 <= a(38) and not w20518;
w20520 <= a(38) and not w20519;
w20521 <= not w20518 and not w20519;
w20522 <= not w20520 and not w20521;
w20523 <= w20511 and not w20522;
w20524 <= w20511 and not w20523;
w20525 <= not w20522 and not w20523;
w20526 <= not w20524 and not w20525;
w20527 <= not w20205 and not w20218;
w20528 <= w20526 and w20527;
w20529 <= not w20526 and not w20527;
w20530 <= not w20528 and not w20529;
w20531 <= b(50) and w4030;
w20532 <= b(48) and w4275;
w20533 <= b(49) and w4025;
w20534 <= not w20532 and not w20533;
w20535 <= not w20531 and w20534;
w20536 <= w4033 and w8692;
w20537 <= w20535 and not w20536;
w20538 <= a(35) and not w20537;
w20539 <= a(35) and not w20538;
w20540 <= not w20537 and not w20538;
w20541 <= not w20539 and not w20540;
w20542 <= w20530 and not w20541;
w20543 <= not w20530 and w20541;
w20544 <= w20358 and not w20543;
w20545 <= not w20542 and w20544;
w20546 <= w20358 and not w20545;
w20547 <= not w20543 and not w20545;
w20548 <= not w20542 and w20547;
w20549 <= not w20546 and not w20548;
w20550 <= not w20343 and w20549;
w20551 <= w20343 and not w20549;
w20552 <= not w20550 and not w20551;
w20553 <= w20327 and not w20552;
w20554 <= w20327 and not w20553;
w20555 <= not w20552 and not w20553;
w20556 <= not w20554 and not w20555;
w20557 <= not w20312 and w20556;
w20558 <= w20312 and not w20556;
w20559 <= not w20557 and not w20558;
w20560 <= not w20296 and not w20559;
w20561 <= w20296 and w20559;
w20562 <= not w20560 and not w20561;
w20563 <= not w20284 and w20562;
w20564 <= w20284 and not w20562;
w20565 <= not w20563 and not w20564;
w20566 <= not w20283 and w20565;
w20567 <= w20283 and not w20565;
w20568 <= not w20566 and not w20567;
w20569 <= not w20312 and not w20556;
w20570 <= not w20309 and not w20569;
w20571 <= b(63) and w1791;
w20572 <= b(61) and w1941;
w20573 <= b(62) and w1786;
w20574 <= not w20572 and not w20573;
w20575 <= not w20571 and w20574;
w20576 <= w1794 and w13514;
w20577 <= w20575 and not w20576;
w20578 <= a(23) and not w20577;
w20579 <= a(23) and not w20578;
w20580 <= not w20577 and not w20578;
w20581 <= not w20579 and not w20580;
w20582 <= not w20570 and not w20581;
w20583 <= not w20570 and not w20582;
w20584 <= not w20581 and not w20582;
w20585 <= not w20583 and not w20584;
w20586 <= b(60) and w2282;
w20587 <= b(58) and w2428;
w20588 <= b(59) and w2277;
w20589 <= not w20587 and not w20588;
w20590 <= not w20586 and w20589;
w20591 <= w2285 and w11954;
w20592 <= w20590 and not w20591;
w20593 <= a(26) and not w20592;
w20594 <= a(26) and not w20593;
w20595 <= not w20592 and not w20593;
w20596 <= not w20594 and not w20595;
w20597 <= not w20326 and not w20553;
w20598 <= w20596 and w20597;
w20599 <= not w20596 and not w20597;
w20600 <= not w20598 and not w20599;
w20601 <= not w20343 and not w20549;
w20602 <= not w20340 and not w20601;
w20603 <= b(57) and w2793;
w20604 <= b(55) and w2986;
w20605 <= b(56) and w2788;
w20606 <= not w20604 and not w20605;
w20607 <= not w20603 and w20606;
w20608 <= w2796 and w11153;
w20609 <= w20607 and not w20608;
w20610 <= a(29) and not w20609;
w20611 <= a(29) and not w20610;
w20612 <= not w20609 and not w20610;
w20613 <= not w20611 and not w20612;
w20614 <= not w20602 and w20613;
w20615 <= w20602 and not w20613;
w20616 <= not w20614 and not w20615;
w20617 <= b(54) and w3381;
w20618 <= b(52) and w3586;
w20619 <= b(53) and w3376;
w20620 <= not w20618 and not w20619;
w20621 <= not w20617 and w20620;
w20622 <= w3384 and w9741;
w20623 <= w20621 and not w20622;
w20624 <= a(32) and not w20623;
w20625 <= a(32) and not w20624;
w20626 <= not w20623 and not w20624;
w20627 <= not w20625 and not w20626;
w20628 <= not w20357 and not w20545;
w20629 <= w20627 and w20628;
w20630 <= not w20627 and not w20628;
w20631 <= not w20629 and not w20630;
w20632 <= not w20529 and not w20542;
w20633 <= not w20485 and not w20488;
w20634 <= b(20) and w13646;
w20635 <= b(21) and not w13231;
w20636 <= not w20634 and not w20635;
w20637 <= not a(20) and not w20636;
w20638 <= a(20) and w20636;
w20639 <= not w20637 and not w20638;
w20640 <= not w20423 and w20639;
w20641 <= w20423 and not w20639;
w20642 <= not w20640 and not w20641;
w20643 <= b(24) and w12411;
w20644 <= b(22) and w12790;
w20645 <= b(23) and w12406;
w20646 <= not w20644 and not w20645;
w20647 <= not w20643 and w20646;
w20648 <= w2201 and w12414;
w20649 <= w20647 and not w20648;
w20650 <= a(62) and not w20649;
w20651 <= a(62) and not w20650;
w20652 <= not w20649 and not w20650;
w20653 <= not w20651 and not w20652;
w20654 <= w20642 and not w20653;
w20655 <= w20642 and not w20654;
w20656 <= not w20653 and not w20654;
w20657 <= not w20655 and not w20656;
w20658 <= not w20424 and not w20438;
w20659 <= not w20657 and not w20658;
w20660 <= not w20657 and not w20659;
w20661 <= not w20658 and not w20659;
w20662 <= not w20660 and not w20661;
w20663 <= b(27) and w11274;
w20664 <= b(25) and w11639;
w20665 <= b(26) and w11269;
w20666 <= not w20664 and not w20665;
w20667 <= not w20663 and w20666;
w20668 <= w2733 and w11277;
w20669 <= w20667 and not w20668;
w20670 <= a(59) and not w20669;
w20671 <= a(59) and not w20670;
w20672 <= not w20669 and not w20670;
w20673 <= not w20671 and not w20672;
w20674 <= not w20662 and not w20673;
w20675 <= not w20662 and not w20674;
w20676 <= not w20673 and not w20674;
w20677 <= not w20675 and not w20676;
w20678 <= not w20441 and not w20444;
w20679 <= w20677 and w20678;
w20680 <= not w20677 and not w20678;
w20681 <= not w20679 and not w20680;
w20682 <= b(30) and w10169;
w20683 <= b(28) and w10539;
w20684 <= b(29) and w10164;
w20685 <= not w20683 and not w20684;
w20686 <= not w20682 and w20685;
w20687 <= w3320 and w10172;
w20688 <= w20686 and not w20687;
w20689 <= a(56) and not w20688;
w20690 <= a(56) and not w20689;
w20691 <= not w20688 and not w20689;
w20692 <= not w20690 and not w20691;
w20693 <= w20681 and not w20692;
w20694 <= w20681 and not w20693;
w20695 <= not w20692 and not w20693;
w20696 <= not w20694 and not w20695;
w20697 <= not w20447 and not w20461;
w20698 <= w20696 and w20697;
w20699 <= not w20696 and not w20697;
w20700 <= not w20698 and not w20699;
w20701 <= b(33) and w9082;
w20702 <= b(31) and w9475;
w20703 <= b(32) and w9077;
w20704 <= not w20702 and not w20703;
w20705 <= not w20701 and w20704;
w20706 <= w3966 and w9085;
w20707 <= w20705 and not w20706;
w20708 <= a(53) and not w20707;
w20709 <= a(53) and not w20708;
w20710 <= not w20707 and not w20708;
w20711 <= not w20709 and not w20710;
w20712 <= not w20470 and not w20481;
w20713 <= not w20467 and not w20712;
w20714 <= not w20711 and not w20713;
w20715 <= w20711 and w20713;
w20716 <= not w20714 and not w20715;
w20717 <= not w20700 and w20716;
w20718 <= w20700 and not w20716;
w20719 <= not w20717 and not w20718;
w20720 <= b(36) and w8105;
w20721 <= b(34) and w8458;
w20722 <= b(35) and w8100;
w20723 <= not w20721 and not w20722;
w20724 <= not w20720 and w20723;
w20725 <= w4665 and w8108;
w20726 <= w20724 and not w20725;
w20727 <= a(50) and not w20726;
w20728 <= a(50) and not w20727;
w20729 <= not w20726 and not w20727;
w20730 <= not w20728 and not w20729;
w20731 <= not w20719 and not w20730;
w20732 <= w20719 and w20730;
w20733 <= not w20731 and not w20732;
w20734 <= w20633 and not w20733;
w20735 <= not w20633 and w20733;
w20736 <= not w20734 and not w20735;
w20737 <= b(39) and w7189;
w20738 <= b(37) and w7530;
w20739 <= b(38) and w7184;
w20740 <= not w20738 and not w20739;
w20741 <= not w20737 and w20740;
w20742 <= w5194 and w7192;
w20743 <= w20741 and not w20742;
w20744 <= a(47) and not w20743;
w20745 <= a(47) and not w20744;
w20746 <= not w20743 and not w20744;
w20747 <= not w20745 and not w20746;
w20748 <= w20736 and not w20747;
w20749 <= w20736 and not w20748;
w20750 <= not w20747 and not w20748;
w20751 <= not w20749 and not w20750;
w20752 <= not w20491 and not w20494;
w20753 <= w20751 and w20752;
w20754 <= not w20751 and not w20752;
w20755 <= not w20753 and not w20754;
w20756 <= b(42) and w6338;
w20757 <= b(40) and w6645;
w20758 <= b(41) and w6333;
w20759 <= not w20757 and not w20758;
w20760 <= not w20756 and w20759;
w20761 <= w6232 and w6341;
w20762 <= w20760 and not w20761;
w20763 <= a(44) and not w20762;
w20764 <= a(44) and not w20763;
w20765 <= not w20762 and not w20763;
w20766 <= not w20764 and not w20765;
w20767 <= w20755 and not w20766;
w20768 <= w20755 and not w20767;
w20769 <= not w20766 and not w20767;
w20770 <= not w20768 and not w20769;
w20771 <= not w20497 and not w20500;
w20772 <= w20770 and w20771;
w20773 <= not w20770 and not w20771;
w20774 <= not w20772 and not w20773;
w20775 <= b(45) and w5520;
w20776 <= b(43) and w5802;
w20777 <= b(44) and w5515;
w20778 <= not w20776 and not w20777;
w20779 <= not w20775 and w20778;
w20780 <= w5523 and w7104;
w20781 <= w20779 and not w20780;
w20782 <= a(41) and not w20781;
w20783 <= a(41) and not w20782;
w20784 <= not w20781 and not w20782;
w20785 <= not w20783 and not w20784;
w20786 <= w20774 and not w20785;
w20787 <= w20774 and not w20786;
w20788 <= not w20785 and not w20786;
w20789 <= not w20787 and not w20788;
w20790 <= not w20503 and not w20506;
w20791 <= w20789 and w20790;
w20792 <= not w20789 and not w20790;
w20793 <= not w20791 and not w20792;
w20794 <= b(48) and w4778;
w20795 <= b(46) and w5020;
w20796 <= b(47) and w4773;
w20797 <= not w20795 and not w20796;
w20798 <= not w20794 and w20797;
w20799 <= w4781 and w7752;
w20800 <= w20798 and not w20799;
w20801 <= a(38) and not w20800;
w20802 <= a(38) and not w20801;
w20803 <= not w20800 and not w20801;
w20804 <= not w20802 and not w20803;
w20805 <= w20793 and not w20804;
w20806 <= w20793 and not w20805;
w20807 <= not w20804 and not w20805;
w20808 <= not w20806 and not w20807;
w20809 <= not w20509 and not w20523;
w20810 <= w20808 and w20809;
w20811 <= not w20808 and not w20809;
w20812 <= not w20810 and not w20811;
w20813 <= b(51) and w4030;
w20814 <= b(49) and w4275;
w20815 <= b(50) and w4025;
w20816 <= not w20814 and not w20815;
w20817 <= not w20813 and w20816;
w20818 <= w4033 and w8719;
w20819 <= w20817 and not w20818;
w20820 <= a(35) and not w20819;
w20821 <= a(35) and not w20820;
w20822 <= not w20819 and not w20820;
w20823 <= not w20821 and not w20822;
w20824 <= w20812 and not w20823;
w20825 <= not w20812 and w20823;
w20826 <= not w20632 and not w20825;
w20827 <= not w20824 and w20826;
w20828 <= not w20632 and not w20827;
w20829 <= not w20824 and not w20827;
w20830 <= not w20825 and w20829;
w20831 <= not w20828 and not w20830;
w20832 <= w20631 and not w20831;
w20833 <= not w20631 and w20831;
w20834 <= not w20616 and not w20833;
w20835 <= not w20832 and w20834;
w20836 <= not w20616 and not w20835;
w20837 <= not w20833 and not w20835;
w20838 <= not w20832 and w20837;
w20839 <= not w20836 and not w20838;
w20840 <= w20600 and not w20839;
w20841 <= not w20600 and w20839;
w20842 <= not w20585 and not w20841;
w20843 <= not w20840 and w20842;
w20844 <= not w20585 and not w20843;
w20845 <= not w20841 and not w20843;
w20846 <= not w20840 and w20845;
w20847 <= not w20844 and not w20846;
w20848 <= not w20293 and not w20560;
w20849 <= w20847 and w20848;
w20850 <= not w20847 and not w20848;
w20851 <= not w20849 and not w20850;
w20852 <= not w20563 and not w20566;
w20853 <= w20851 and not w20852;
w20854 <= not w20851 and w20852;
w20855 <= not w20853 and not w20854;
w20856 <= not w20599 and not w20840;
w20857 <= b(62) and w1941;
w20858 <= b(63) and w1786;
w20859 <= not w20857 and not w20858;
w20860 <= not w1794 and w20859;
w20861 <= w13543 and w20859;
w20862 <= not w20860 and not w20861;
w20863 <= a(23) and not w20862;
w20864 <= not a(23) and w20862;
w20865 <= not w20863 and not w20864;
w20866 <= not w20856 and not w20865;
w20867 <= w20856 and w20865;
w20868 <= not w20866 and not w20867;
w20869 <= b(61) and w2282;
w20870 <= b(59) and w2428;
w20871 <= b(60) and w2277;
w20872 <= not w20870 and not w20871;
w20873 <= not w20869 and w20872;
w20874 <= w2285 and w12712;
w20875 <= w20873 and not w20874;
w20876 <= a(26) and not w20875;
w20877 <= a(26) and not w20876;
w20878 <= not w20875 and not w20876;
w20879 <= not w20877 and not w20878;
w20880 <= not w20602 and not w20613;
w20881 <= not w20835 and not w20880;
w20882 <= w20879 and w20881;
w20883 <= not w20879 and not w20881;
w20884 <= not w20882 and not w20883;
w20885 <= not w20630 and not w20832;
w20886 <= b(58) and w2793;
w20887 <= b(56) and w2986;
w20888 <= b(57) and w2788;
w20889 <= not w20887 and not w20888;
w20890 <= not w20886 and w20889;
w20891 <= not w2796 and w20890;
w20892 <= not w11179 and w20890;
w20893 <= not w20891 and not w20892;
w20894 <= a(29) and not w20893;
w20895 <= not a(29) and w20893;
w20896 <= not w20894 and not w20895;
w20897 <= not w20885 and not w20896;
w20898 <= w20885 and w20896;
w20899 <= not w20897 and not w20898;
w20900 <= b(55) and w3381;
w20901 <= b(53) and w3586;
w20902 <= b(54) and w3376;
w20903 <= not w20901 and not w20902;
w20904 <= not w20900 and w20903;
w20905 <= w3384 and w10427;
w20906 <= w20904 and not w20905;
w20907 <= a(32) and not w20906;
w20908 <= a(32) and not w20907;
w20909 <= not w20906 and not w20907;
w20910 <= not w20908 and not w20909;
w20911 <= not w20829 and w20910;
w20912 <= w20829 and not w20910;
w20913 <= not w20911 and not w20912;
w20914 <= b(43) and w6338;
w20915 <= b(41) and w6645;
w20916 <= b(42) and w6333;
w20917 <= not w20915 and not w20916;
w20918 <= not w20914 and w20917;
w20919 <= w6258 and w6341;
w20920 <= w20918 and not w20919;
w20921 <= a(44) and not w20920;
w20922 <= a(44) and not w20921;
w20923 <= not w20920 and not w20921;
w20924 <= not w20922 and not w20923;
w20925 <= not w20748 and not w20754;
w20926 <= b(40) and w7189;
w20927 <= b(38) and w7530;
w20928 <= b(39) and w7184;
w20929 <= not w20927 and not w20928;
w20930 <= not w20926 and w20929;
w20931 <= w5698 and w7192;
w20932 <= w20930 and not w20931;
w20933 <= a(47) and not w20932;
w20934 <= a(47) and not w20933;
w20935 <= not w20932 and not w20933;
w20936 <= not w20934 and not w20935;
w20937 <= not w20731 and not w20735;
w20938 <= not w20674 and not w20680;
w20939 <= b(28) and w11274;
w20940 <= b(26) and w11639;
w20941 <= b(27) and w11269;
w20942 <= not w20940 and not w20941;
w20943 <= not w20939 and w20942;
w20944 <= w2932 and w11277;
w20945 <= w20943 and not w20944;
w20946 <= a(59) and not w20945;
w20947 <= a(59) and not w20946;
w20948 <= not w20945 and not w20946;
w20949 <= not w20947 and not w20948;
w20950 <= not w20654 and not w20659;
w20951 <= b(21) and w13646;
w20952 <= b(22) and not w13231;
w20953 <= not w20951 and not w20952;
w20954 <= not w20637 and not w20640;
w20955 <= not w20953 and w20954;
w20956 <= w20953 and not w20954;
w20957 <= not w20955 and not w20956;
w20958 <= b(25) and w12411;
w20959 <= b(23) and w12790;
w20960 <= b(24) and w12406;
w20961 <= not w20959 and not w20960;
w20962 <= not w20958 and w20961;
w20963 <= not w12414 and w20962;
w20964 <= not w2228 and w20962;
w20965 <= not w20963 and not w20964;
w20966 <= a(62) and not w20965;
w20967 <= not a(62) and w20965;
w20968 <= not w20966 and not w20967;
w20969 <= w20957 and not w20968;
w20970 <= not w20957 and w20968;
w20971 <= not w20969 and not w20970;
w20972 <= not w20950 and w20971;
w20973 <= w20950 and not w20971;
w20974 <= not w20972 and not w20973;
w20975 <= not w20949 and w20974;
w20976 <= w20949 and not w20974;
w20977 <= not w20975 and not w20976;
w20978 <= not w20938 and w20977;
w20979 <= w20938 and not w20977;
w20980 <= not w20978 and not w20979;
w20981 <= b(31) and w10169;
w20982 <= b(29) and w10539;
w20983 <= b(30) and w10164;
w20984 <= not w20982 and not w20983;
w20985 <= not w20981 and w20984;
w20986 <= w3539 and w10172;
w20987 <= w20985 and not w20986;
w20988 <= a(56) and not w20987;
w20989 <= a(56) and not w20988;
w20990 <= not w20987 and not w20988;
w20991 <= not w20989 and not w20990;
w20992 <= w20980 and not w20991;
w20993 <= w20980 and not w20992;
w20994 <= not w20991 and not w20992;
w20995 <= not w20993 and not w20994;
w20996 <= not w20693 and not w20699;
w20997 <= w20995 and w20996;
w20998 <= not w20995 and not w20996;
w20999 <= not w20997 and not w20998;
w21000 <= b(34) and w9082;
w21001 <= b(32) and w9475;
w21002 <= b(33) and w9077;
w21003 <= not w21001 and not w21002;
w21004 <= not w21000 and w21003;
w21005 <= w4209 and w9085;
w21006 <= w21004 and not w21005;
w21007 <= a(53) and not w21006;
w21008 <= a(53) and not w21007;
w21009 <= not w21006 and not w21007;
w21010 <= not w21008 and not w21009;
w21011 <= w20999 and not w21010;
w21012 <= w20999 and not w21011;
w21013 <= not w21010 and not w21011;
w21014 <= not w21012 and not w21013;
w21015 <= w20700 and w20716;
w21016 <= not w20714 and not w21015;
w21017 <= w21014 and w21016;
w21018 <= not w21014 and not w21016;
w21019 <= not w21017 and not w21018;
w21020 <= b(37) and w8105;
w21021 <= b(35) and w8458;
w21022 <= b(36) and w8100;
w21023 <= not w21021 and not w21022;
w21024 <= not w21020 and w21023;
w21025 <= w4924 and w8108;
w21026 <= w21024 and not w21025;
w21027 <= a(50) and not w21026;
w21028 <= a(50) and not w21027;
w21029 <= not w21026 and not w21027;
w21030 <= not w21028 and not w21029;
w21031 <= not w21019 and w21030;
w21032 <= w21019 and not w21030;
w21033 <= not w21031 and not w21032;
w21034 <= not w20937 and w21033;
w21035 <= not w20937 and not w21034;
w21036 <= w21033 and not w21034;
w21037 <= not w21035 and not w21036;
w21038 <= not w20936 and not w21037;
w21039 <= w20936 and not w21036;
w21040 <= not w21035 and w21039;
w21041 <= not w21038 and not w21040;
w21042 <= not w20925 and w21041;
w21043 <= w20925 and not w21041;
w21044 <= not w21042 and not w21043;
w21045 <= not w20924 and w21044;
w21046 <= w21044 and not w21045;
w21047 <= not w20924 and not w21045;
w21048 <= not w21046 and not w21047;
w21049 <= not w20767 and not w20773;
w21050 <= w21048 and w21049;
w21051 <= not w21048 and not w21049;
w21052 <= not w21050 and not w21051;
w21053 <= b(46) and w5520;
w21054 <= b(44) and w5802;
w21055 <= b(45) and w5515;
w21056 <= not w21054 and not w21055;
w21057 <= not w21053 and w21056;
w21058 <= w5523 and w7420;
w21059 <= w21057 and not w21058;
w21060 <= a(41) and not w21059;
w21061 <= a(41) and not w21060;
w21062 <= not w21059 and not w21060;
w21063 <= not w21061 and not w21062;
w21064 <= w21052 and not w21063;
w21065 <= w21052 and not w21064;
w21066 <= not w21063 and not w21064;
w21067 <= not w21065 and not w21066;
w21068 <= not w20786 and not w20792;
w21069 <= w21067 and w21068;
w21070 <= not w21067 and not w21068;
w21071 <= not w21069 and not w21070;
w21072 <= b(49) and w4778;
w21073 <= b(47) and w5020;
w21074 <= b(48) and w4773;
w21075 <= not w21073 and not w21074;
w21076 <= not w21072 and w21075;
w21077 <= w4781 and w8368;
w21078 <= w21076 and not w21077;
w21079 <= a(38) and not w21078;
w21080 <= a(38) and not w21079;
w21081 <= not w21078 and not w21079;
w21082 <= not w21080 and not w21081;
w21083 <= w21071 and not w21082;
w21084 <= w21071 and not w21083;
w21085 <= not w21082 and not w21083;
w21086 <= not w21084 and not w21085;
w21087 <= not w20805 and not w20811;
w21088 <= w21086 and w21087;
w21089 <= not w21086 and not w21087;
w21090 <= not w21088 and not w21089;
w21091 <= b(52) and w4030;
w21092 <= b(50) and w4275;
w21093 <= b(51) and w4025;
w21094 <= not w21092 and not w21093;
w21095 <= not w21091 and w21094;
w21096 <= w4033 and w9371;
w21097 <= w21095 and not w21096;
w21098 <= a(35) and not w21097;
w21099 <= a(35) and not w21098;
w21100 <= not w21097 and not w21098;
w21101 <= not w21099 and not w21100;
w21102 <= w21090 and not w21101;
w21103 <= w21090 and not w21102;
w21104 <= not w21101 and not w21102;
w21105 <= not w21103 and not w21104;
w21106 <= not w20913 and not w21105;
w21107 <= w20913 and w21105;
w21108 <= w20899 and not w21107;
w21109 <= not w21106 and w21108;
w21110 <= w20899 and not w21109;
w21111 <= not w21107 and not w21109;
w21112 <= not w21106 and w21111;
w21113 <= not w21110 and not w21112;
w21114 <= w20884 and not w21113;
w21115 <= not w20884 and w21113;
w21116 <= w20868 and not w21115;
w21117 <= not w21114 and w21116;
w21118 <= w20868 and not w21117;
w21119 <= not w21115 and not w21117;
w21120 <= not w21114 and w21119;
w21121 <= not w21118 and not w21120;
w21122 <= not w20582 and not w20843;
w21123 <= w21121 and w21122;
w21124 <= not w21121 and not w21122;
w21125 <= not w21123 and not w21124;
w21126 <= not w20850 and not w20853;
w21127 <= w21125 and not w21126;
w21128 <= not w21125 and w21126;
w21129 <= not w21127 and not w21128;
w21130 <= not w21124 and not w21127;
w21131 <= not w20866 and not w21117;
w21132 <= not w20883 and not w21114;
w21133 <= b(63) and w1941;
w21134 <= w1794 and w13540;
w21135 <= not w21133 and not w21134;
w21136 <= a(23) and not w21135;
w21137 <= a(23) and not w21136;
w21138 <= not w21135 and not w21136;
w21139 <= not w21137 and not w21138;
w21140 <= not w21132 and not w21139;
w21141 <= not w21132 and not w21140;
w21142 <= not w21139 and not w21140;
w21143 <= not w21141 and not w21142;
w21144 <= b(62) and w2282;
w21145 <= b(60) and w2428;
w21146 <= b(61) and w2277;
w21147 <= not w21145 and not w21146;
w21148 <= not w21144 and w21147;
w21149 <= w2285 and w13113;
w21150 <= w21148 and not w21149;
w21151 <= a(26) and not w21150;
w21152 <= a(26) and not w21151;
w21153 <= not w21150 and not w21151;
w21154 <= not w21152 and not w21153;
w21155 <= not w20897 and not w21109;
w21156 <= w21154 and w21155;
w21157 <= not w21154 and not w21155;
w21158 <= not w21156 and not w21157;
w21159 <= b(59) and w2793;
w21160 <= b(57) and w2986;
w21161 <= b(58) and w2788;
w21162 <= not w21160 and not w21161;
w21163 <= not w21159 and w21162;
w21164 <= w2796 and w11922;
w21165 <= w21163 and not w21164;
w21166 <= a(29) and not w21165;
w21167 <= a(29) and not w21166;
w21168 <= not w21165 and not w21166;
w21169 <= not w21167 and not w21168;
w21170 <= not w20829 and not w20910;
w21171 <= not w21106 and not w21170;
w21172 <= not w21169 and not w21171;
w21173 <= not w21169 and not w21172;
w21174 <= not w21171 and not w21172;
w21175 <= not w21173 and not w21174;
w21176 <= b(56) and w3381;
w21177 <= b(54) and w3586;
w21178 <= b(55) and w3376;
w21179 <= not w21177 and not w21178;
w21180 <= not w21176 and w21179;
w21181 <= w3384 and w10451;
w21182 <= w21180 and not w21181;
w21183 <= a(32) and not w21182;
w21184 <= a(32) and not w21183;
w21185 <= not w21182 and not w21183;
w21186 <= not w21184 and not w21185;
w21187 <= not w21089 and not w21102;
w21188 <= w21186 and w21187;
w21189 <= not w21186 and not w21187;
w21190 <= not w21188 and not w21189;
w21191 <= b(53) and w4030;
w21192 <= b(51) and w4275;
w21193 <= b(52) and w4025;
w21194 <= not w21192 and not w21193;
w21195 <= not w21191 and w21194;
w21196 <= w4033 and w9715;
w21197 <= w21195 and not w21196;
w21198 <= a(35) and not w21197;
w21199 <= a(35) and not w21198;
w21200 <= not w21197 and not w21198;
w21201 <= not w21199 and not w21200;
w21202 <= not w21070 and not w21083;
w21203 <= not w21042 and not w21045;
w21204 <= b(44) and w6338;
w21205 <= b(42) and w6645;
w21206 <= b(43) and w6333;
w21207 <= not w21205 and not w21206;
w21208 <= not w21204 and w21207;
w21209 <= w6341 and w6815;
w21210 <= w21208 and not w21209;
w21211 <= a(44) and not w21210;
w21212 <= a(44) and not w21211;
w21213 <= not w21210 and not w21211;
w21214 <= not w21212 and not w21213;
w21215 <= not w21034 and not w21038;
w21216 <= not w20998 and not w21011;
w21217 <= b(35) and w9082;
w21218 <= b(33) and w9475;
w21219 <= b(34) and w9077;
w21220 <= not w21218 and not w21219;
w21221 <= not w21217 and w21220;
w21222 <= w4439 and w9085;
w21223 <= w21221 and not w21222;
w21224 <= a(53) and not w21223;
w21225 <= a(53) and not w21224;
w21226 <= not w21223 and not w21224;
w21227 <= not w21225 and not w21226;
w21228 <= not w20978 and not w20992;
w21229 <= not w20956 and not w20969;
w21230 <= b(22) and w13646;
w21231 <= b(23) and not w13231;
w21232 <= not w21230 and not w21231;
w21233 <= not w20953 and w21232;
w21234 <= w20953 and not w21232;
w21235 <= not w21233 and not w21234;
w21236 <= b(26) and w12411;
w21237 <= b(24) and w12790;
w21238 <= b(25) and w12406;
w21239 <= not w21237 and not w21238;
w21240 <= not w21236 and w21239;
w21241 <= not w12414 and w21240;
w21242 <= not w2556 and w21240;
w21243 <= not w21241 and not w21242;
w21244 <= a(62) and not w21243;
w21245 <= not a(62) and w21243;
w21246 <= not w21244 and not w21245;
w21247 <= w21235 and not w21246;
w21248 <= not w21235 and w21246;
w21249 <= not w21247 and not w21248;
w21250 <= not w21229 and w21249;
w21251 <= w21229 and not w21249;
w21252 <= not w21250 and not w21251;
w21253 <= b(29) and w11274;
w21254 <= b(27) and w11639;
w21255 <= b(28) and w11269;
w21256 <= not w21254 and not w21255;
w21257 <= not w21253 and w21256;
w21258 <= w3126 and w11277;
w21259 <= w21257 and not w21258;
w21260 <= a(59) and not w21259;
w21261 <= a(59) and not w21260;
w21262 <= not w21259 and not w21260;
w21263 <= not w21261 and not w21262;
w21264 <= w21252 and not w21263;
w21265 <= w21252 and not w21264;
w21266 <= not w21263 and not w21264;
w21267 <= not w21265 and not w21266;
w21268 <= not w20972 and not w20975;
w21269 <= w21267 and w21268;
w21270 <= not w21267 and not w21268;
w21271 <= not w21269 and not w21270;
w21272 <= b(32) and w10169;
w21273 <= b(30) and w10539;
w21274 <= b(31) and w10164;
w21275 <= not w21273 and not w21274;
w21276 <= not w21272 and w21275;
w21277 <= w3756 and w10172;
w21278 <= w21276 and not w21277;
w21279 <= a(56) and not w21278;
w21280 <= a(56) and not w21279;
w21281 <= not w21278 and not w21279;
w21282 <= not w21280 and not w21281;
w21283 <= not w21271 and w21282;
w21284 <= w21271 and not w21282;
w21285 <= not w21283 and not w21284;
w21286 <= not w21228 and w21285;
w21287 <= w21228 and not w21285;
w21288 <= not w21286 and not w21287;
w21289 <= not w21227 and w21288;
w21290 <= w21227 and not w21288;
w21291 <= not w21289 and not w21290;
w21292 <= not w21216 and w21291;
w21293 <= w21216 and not w21291;
w21294 <= not w21292 and not w21293;
w21295 <= b(38) and w8105;
w21296 <= b(36) and w8458;
w21297 <= b(37) and w8100;
w21298 <= not w21296 and not w21297;
w21299 <= not w21295 and w21298;
w21300 <= w4948 and w8108;
w21301 <= w21299 and not w21300;
w21302 <= a(50) and not w21301;
w21303 <= a(50) and not w21302;
w21304 <= not w21301 and not w21302;
w21305 <= not w21303 and not w21304;
w21306 <= w21294 and not w21305;
w21307 <= w21294 and not w21306;
w21308 <= not w21305 and not w21306;
w21309 <= not w21307 and not w21308;
w21310 <= not w21018 and not w21032;
w21311 <= not w21309 and not w21310;
w21312 <= not w21309 and not w21311;
w21313 <= not w21310 and not w21311;
w21314 <= not w21312 and not w21313;
w21315 <= b(41) and w7189;
w21316 <= b(39) and w7530;
w21317 <= b(40) and w7184;
w21318 <= not w21316 and not w21317;
w21319 <= not w21315 and w21318;
w21320 <= w5962 and w7192;
w21321 <= w21319 and not w21320;
w21322 <= a(47) and not w21321;
w21323 <= a(47) and not w21322;
w21324 <= not w21321 and not w21322;
w21325 <= not w21323 and not w21324;
w21326 <= not w21314 and w21325;
w21327 <= w21314 and not w21325;
w21328 <= not w21326 and not w21327;
w21329 <= not w21215 and not w21328;
w21330 <= w21215 and w21328;
w21331 <= not w21329 and not w21330;
w21332 <= not w21214 and w21331;
w21333 <= w21214 and not w21331;
w21334 <= not w21332 and not w21333;
w21335 <= not w21203 and w21334;
w21336 <= w21203 and not w21334;
w21337 <= not w21335 and not w21336;
w21338 <= b(47) and w5520;
w21339 <= b(45) and w5802;
w21340 <= b(46) and w5515;
w21341 <= not w21339 and not w21340;
w21342 <= not w21338 and w21341;
w21343 <= w5523 and w7446;
w21344 <= w21342 and not w21343;
w21345 <= a(41) and not w21344;
w21346 <= a(41) and not w21345;
w21347 <= not w21344 and not w21345;
w21348 <= not w21346 and not w21347;
w21349 <= w21337 and not w21348;
w21350 <= w21337 and not w21349;
w21351 <= not w21348 and not w21349;
w21352 <= not w21350 and not w21351;
w21353 <= not w21051 and not w21064;
w21354 <= w21352 and w21353;
w21355 <= not w21352 and not w21353;
w21356 <= not w21354 and not w21355;
w21357 <= b(50) and w4778;
w21358 <= b(48) and w5020;
w21359 <= b(49) and w4773;
w21360 <= not w21358 and not w21359;
w21361 <= not w21357 and w21360;
w21362 <= w4781 and w8692;
w21363 <= w21361 and not w21362;
w21364 <= a(38) and not w21363;
w21365 <= a(38) and not w21364;
w21366 <= not w21363 and not w21364;
w21367 <= not w21365 and not w21366;
w21368 <= not w21356 and w21367;
w21369 <= w21356 and not w21367;
w21370 <= not w21368 and not w21369;
w21371 <= not w21202 and w21370;
w21372 <= not w21202 and not w21371;
w21373 <= w21370 and not w21371;
w21374 <= not w21372 and not w21373;
w21375 <= not w21201 and not w21374;
w21376 <= not w21201 and not w21375;
w21377 <= not w21374 and not w21375;
w21378 <= not w21376 and not w21377;
w21379 <= w21190 and not w21378;
w21380 <= w21190 and not w21379;
w21381 <= not w21378 and not w21379;
w21382 <= not w21380 and not w21381;
w21383 <= not w21175 and w21382;
w21384 <= w21175 and not w21382;
w21385 <= not w21383 and not w21384;
w21386 <= w21158 and not w21385;
w21387 <= w21158 and not w21386;
w21388 <= not w21385 and not w21386;
w21389 <= not w21387 and not w21388;
w21390 <= not w21143 and w21389;
w21391 <= w21143 and not w21389;
w21392 <= not w21390 and not w21391;
w21393 <= not w21131 and not w21392;
w21394 <= not w21131 and not w21393;
w21395 <= not w21392 and not w21393;
w21396 <= not w21394 and not w21395;
w21397 <= not w21130 and not w21396;
w21398 <= w21130 and not w21395;
w21399 <= not w21394 and w21398;
w21400 <= not w21397 and not w21399;
w21401 <= not w21393 and not w21397;
w21402 <= not w21143 and not w21389;
w21403 <= not w21140 and not w21402;
w21404 <= not w21157 and not w21386;
w21405 <= b(63) and w2282;
w21406 <= b(61) and w2428;
w21407 <= b(62) and w2277;
w21408 <= not w21406 and not w21407;
w21409 <= not w21405 and w21408;
w21410 <= w2285 and w13514;
w21411 <= w21409 and not w21410;
w21412 <= a(26) and not w21411;
w21413 <= a(26) and not w21412;
w21414 <= not w21411 and not w21412;
w21415 <= not w21413 and not w21414;
w21416 <= not w21404 and not w21415;
w21417 <= not w21404 and not w21416;
w21418 <= not w21415 and not w21416;
w21419 <= not w21417 and not w21418;
w21420 <= not w21175 and not w21382;
w21421 <= not w21172 and not w21420;
w21422 <= b(60) and w2793;
w21423 <= b(58) and w2986;
w21424 <= b(59) and w2788;
w21425 <= not w21423 and not w21424;
w21426 <= not w21422 and w21425;
w21427 <= w2796 and w11954;
w21428 <= w21426 and not w21427;
w21429 <= a(29) and not w21428;
w21430 <= a(29) and not w21429;
w21431 <= not w21428 and not w21429;
w21432 <= not w21430 and not w21431;
w21433 <= not w21421 and w21432;
w21434 <= w21421 and not w21432;
w21435 <= not w21433 and not w21434;
w21436 <= b(57) and w3381;
w21437 <= b(55) and w3586;
w21438 <= b(56) and w3376;
w21439 <= not w21437 and not w21438;
w21440 <= not w21436 and w21439;
w21441 <= w3384 and w11153;
w21442 <= w21440 and not w21441;
w21443 <= a(32) and not w21442;
w21444 <= a(32) and not w21443;
w21445 <= not w21442 and not w21443;
w21446 <= not w21444 and not w21445;
w21447 <= not w21189 and not w21379;
w21448 <= w21446 and w21447;
w21449 <= not w21446 and not w21447;
w21450 <= not w21448 and not w21449;
w21451 <= not w21371 and not w21375;
w21452 <= not w21355 and not w21369;
w21453 <= not w21329 and not w21332;
w21454 <= not w21314 and not w21325;
w21455 <= not w21311 and not w21454;
w21456 <= b(36) and w9082;
w21457 <= b(34) and w9475;
w21458 <= b(35) and w9077;
w21459 <= not w21457 and not w21458;
w21460 <= not w21456 and w21459;
w21461 <= w4665 and w9085;
w21462 <= w21460 and not w21461;
w21463 <= a(53) and not w21462;
w21464 <= a(53) and not w21463;
w21465 <= not w21462 and not w21463;
w21466 <= not w21464 and not w21465;
w21467 <= not w21250 and not w21264;
w21468 <= not w21233 and not w21247;
w21469 <= b(23) and w13646;
w21470 <= b(24) and not w13231;
w21471 <= not w21469 and not w21470;
w21472 <= not a(23) and not w21471;
w21473 <= a(23) and w21471;
w21474 <= not w21472 and not w21473;
w21475 <= not w21232 and w21474;
w21476 <= w21232 and not w21474;
w21477 <= not w21475 and not w21476;
w21478 <= b(27) and w12411;
w21479 <= b(25) and w12790;
w21480 <= b(26) and w12406;
w21481 <= not w21479 and not w21480;
w21482 <= not w21478 and w21481;
w21483 <= w2733 and w12414;
w21484 <= w21482 and not w21483;
w21485 <= a(62) and not w21484;
w21486 <= a(62) and not w21485;
w21487 <= not w21484 and not w21485;
w21488 <= not w21486 and not w21487;
w21489 <= w21477 and not w21488;
w21490 <= w21477 and not w21489;
w21491 <= not w21488 and not w21489;
w21492 <= not w21490 and not w21491;
w21493 <= not w21468 and w21492;
w21494 <= w21468 and not w21492;
w21495 <= not w21493 and not w21494;
w21496 <= b(30) and w11274;
w21497 <= b(28) and w11639;
w21498 <= b(29) and w11269;
w21499 <= not w21497 and not w21498;
w21500 <= not w21496 and w21499;
w21501 <= w3320 and w11277;
w21502 <= w21500 and not w21501;
w21503 <= a(59) and not w21502;
w21504 <= a(59) and not w21503;
w21505 <= not w21502 and not w21503;
w21506 <= not w21504 and not w21505;
w21507 <= not w21495 and not w21506;
w21508 <= w21495 and w21506;
w21509 <= not w21507 and not w21508;
w21510 <= w21467 and not w21509;
w21511 <= not w21467 and w21509;
w21512 <= not w21510 and not w21511;
w21513 <= b(33) and w10169;
w21514 <= b(31) and w10539;
w21515 <= b(32) and w10164;
w21516 <= not w21514 and not w21515;
w21517 <= not w21513 and w21516;
w21518 <= w3966 and w10172;
w21519 <= w21517 and not w21518;
w21520 <= a(56) and not w21519;
w21521 <= a(56) and not w21520;
w21522 <= not w21519 and not w21520;
w21523 <= not w21521 and not w21522;
w21524 <= not w21270 and not w21284;
w21525 <= not w21523 and not w21524;
w21526 <= w21523 and w21524;
w21527 <= not w21525 and not w21526;
w21528 <= w21512 and w21527;
w21529 <= not w21512 and not w21527;
w21530 <= not w21528 and not w21529;
w21531 <= not w21466 and w21530;
w21532 <= w21530 and not w21531;
w21533 <= not w21466 and not w21531;
w21534 <= not w21532 and not w21533;
w21535 <= not w21286 and not w21289;
w21536 <= w21534 and w21535;
w21537 <= not w21534 and not w21535;
w21538 <= not w21536 and not w21537;
w21539 <= b(39) and w8105;
w21540 <= b(37) and w8458;
w21541 <= b(38) and w8100;
w21542 <= not w21540 and not w21541;
w21543 <= not w21539 and w21542;
w21544 <= w5194 and w8108;
w21545 <= w21543 and not w21544;
w21546 <= a(50) and not w21545;
w21547 <= a(50) and not w21546;
w21548 <= not w21545 and not w21546;
w21549 <= not w21547 and not w21548;
w21550 <= w21538 and not w21549;
w21551 <= w21538 and not w21550;
w21552 <= not w21549 and not w21550;
w21553 <= not w21551 and not w21552;
w21554 <= not w21292 and not w21306;
w21555 <= w21553 and w21554;
w21556 <= not w21553 and not w21554;
w21557 <= not w21555 and not w21556;
w21558 <= b(42) and w7189;
w21559 <= b(40) and w7530;
w21560 <= b(41) and w7184;
w21561 <= not w21559 and not w21560;
w21562 <= not w21558 and w21561;
w21563 <= w6232 and w7192;
w21564 <= w21562 and not w21563;
w21565 <= a(47) and not w21564;
w21566 <= a(47) and not w21565;
w21567 <= not w21564 and not w21565;
w21568 <= not w21566 and not w21567;
w21569 <= w21557 and not w21568;
w21570 <= w21557 and not w21569;
w21571 <= not w21568 and not w21569;
w21572 <= not w21570 and not w21571;
w21573 <= not w21455 and w21572;
w21574 <= w21455 and not w21572;
w21575 <= not w21573 and not w21574;
w21576 <= b(45) and w6338;
w21577 <= b(43) and w6645;
w21578 <= b(44) and w6333;
w21579 <= not w21577 and not w21578;
w21580 <= not w21576 and w21579;
w21581 <= w6341 and w7104;
w21582 <= w21580 and not w21581;
w21583 <= a(44) and not w21582;
w21584 <= a(44) and not w21583;
w21585 <= not w21582 and not w21583;
w21586 <= not w21584 and not w21585;
w21587 <= not w21575 and not w21586;
w21588 <= w21575 and w21586;
w21589 <= not w21587 and not w21588;
w21590 <= w21453 and not w21589;
w21591 <= not w21453 and w21589;
w21592 <= not w21590 and not w21591;
w21593 <= b(48) and w5520;
w21594 <= b(46) and w5802;
w21595 <= b(47) and w5515;
w21596 <= not w21594 and not w21595;
w21597 <= not w21593 and w21596;
w21598 <= w5523 and w7752;
w21599 <= w21597 and not w21598;
w21600 <= a(41) and not w21599;
w21601 <= a(41) and not w21600;
w21602 <= not w21599 and not w21600;
w21603 <= not w21601 and not w21602;
w21604 <= w21592 and not w21603;
w21605 <= w21592 and not w21604;
w21606 <= not w21603 and not w21604;
w21607 <= not w21605 and not w21606;
w21608 <= not w21335 and not w21349;
w21609 <= w21607 and w21608;
w21610 <= not w21607 and not w21608;
w21611 <= not w21609 and not w21610;
w21612 <= b(51) and w4778;
w21613 <= b(49) and w5020;
w21614 <= b(50) and w4773;
w21615 <= not w21613 and not w21614;
w21616 <= not w21612 and w21615;
w21617 <= w4781 and w8719;
w21618 <= w21616 and not w21617;
w21619 <= a(38) and not w21618;
w21620 <= a(38) and not w21619;
w21621 <= not w21618 and not w21619;
w21622 <= not w21620 and not w21621;
w21623 <= w21611 and not w21622;
w21624 <= not w21611 and w21622;
w21625 <= not w21452 and not w21624;
w21626 <= not w21623 and w21625;
w21627 <= not w21452 and not w21626;
w21628 <= not w21623 and not w21626;
w21629 <= not w21624 and w21628;
w21630 <= not w21627 and not w21629;
w21631 <= b(54) and w4030;
w21632 <= b(52) and w4275;
w21633 <= b(53) and w4025;
w21634 <= not w21632 and not w21633;
w21635 <= not w21631 and w21634;
w21636 <= w4033 and w9741;
w21637 <= w21635 and not w21636;
w21638 <= a(35) and not w21637;
w21639 <= a(35) and not w21638;
w21640 <= not w21637 and not w21638;
w21641 <= not w21639 and not w21640;
w21642 <= w21630 and w21641;
w21643 <= not w21630 and not w21641;
w21644 <= not w21642 and not w21643;
w21645 <= not w21451 and w21644;
w21646 <= w21451 and not w21644;
w21647 <= not w21645 and not w21646;
w21648 <= w21450 and w21647;
w21649 <= not w21450 and not w21647;
w21650 <= not w21435 and not w21649;
w21651 <= not w21648 and w21650;
w21652 <= not w21435 and not w21651;
w21653 <= not w21649 and not w21651;
w21654 <= not w21648 and w21653;
w21655 <= not w21652 and not w21654;
w21656 <= not w21419 and w21655;
w21657 <= w21419 and not w21655;
w21658 <= not w21656 and not w21657;
w21659 <= not w21403 and not w21658;
w21660 <= not w21403 and not w21659;
w21661 <= not w21658 and not w21659;
w21662 <= not w21660 and not w21661;
w21663 <= not w21401 and not w21662;
w21664 <= w21401 and not w21661;
w21665 <= not w21660 and w21664;
w21666 <= not w21663 and not w21665;
w21667 <= not w21659 and not w21663;
w21668 <= not w21419 and not w21655;
w21669 <= not w21416 and not w21668;
w21670 <= b(61) and w2793;
w21671 <= b(59) and w2986;
w21672 <= b(60) and w2788;
w21673 <= not w21671 and not w21672;
w21674 <= not w21670 and w21673;
w21675 <= w2796 and w12712;
w21676 <= w21674 and not w21675;
w21677 <= a(29) and not w21676;
w21678 <= a(29) and not w21677;
w21679 <= not w21676 and not w21677;
w21680 <= not w21678 and not w21679;
w21681 <= not w21449 and not w21648;
w21682 <= not w21680 and not w21681;
w21683 <= not w21680 and not w21682;
w21684 <= not w21681 and not w21682;
w21685 <= not w21683 and not w21684;
w21686 <= not w21643 and not w21645;
w21687 <= b(58) and w3381;
w21688 <= b(56) and w3586;
w21689 <= b(57) and w3376;
w21690 <= not w21688 and not w21689;
w21691 <= not w21687 and w21690;
w21692 <= not w3384 and w21691;
w21693 <= not w11179 and w21691;
w21694 <= not w21692 and not w21693;
w21695 <= a(32) and not w21694;
w21696 <= not a(32) and w21694;
w21697 <= not w21695 and not w21696;
w21698 <= not w21686 and not w21697;
w21699 <= w21686 and w21697;
w21700 <= not w21698 and not w21699;
w21701 <= b(43) and w7189;
w21702 <= b(41) and w7530;
w21703 <= b(42) and w7184;
w21704 <= not w21702 and not w21703;
w21705 <= not w21701 and w21704;
w21706 <= w6258 and w7192;
w21707 <= w21705 and not w21706;
w21708 <= a(47) and not w21707;
w21709 <= a(47) and not w21708;
w21710 <= not w21707 and not w21708;
w21711 <= not w21709 and not w21710;
w21712 <= not w21550 and not w21556;
w21713 <= b(40) and w8105;
w21714 <= b(38) and w8458;
w21715 <= b(39) and w8100;
w21716 <= not w21714 and not w21715;
w21717 <= not w21713 and w21716;
w21718 <= w5698 and w8108;
w21719 <= w21717 and not w21718;
w21720 <= a(50) and not w21719;
w21721 <= a(50) and not w21720;
w21722 <= not w21719 and not w21720;
w21723 <= not w21721 and not w21722;
w21724 <= not w21531 and not w21537;
w21725 <= not w21468 and not w21492;
w21726 <= not w21489 and not w21725;
w21727 <= b(24) and w13646;
w21728 <= b(25) and not w13231;
w21729 <= not w21727 and not w21728;
w21730 <= not w21472 and not w21475;
w21731 <= not w21729 and w21730;
w21732 <= w21729 and not w21730;
w21733 <= not w21731 and not w21732;
w21734 <= b(28) and w12411;
w21735 <= b(26) and w12790;
w21736 <= b(27) and w12406;
w21737 <= not w21735 and not w21736;
w21738 <= not w21734 and w21737;
w21739 <= not w12414 and w21738;
w21740 <= not w2932 and w21738;
w21741 <= not w21739 and not w21740;
w21742 <= a(62) and not w21741;
w21743 <= not a(62) and w21741;
w21744 <= not w21742 and not w21743;
w21745 <= w21733 and not w21744;
w21746 <= not w21733 and w21744;
w21747 <= not w21745 and not w21746;
w21748 <= not w21726 and w21747;
w21749 <= w21726 and not w21747;
w21750 <= not w21748 and not w21749;
w21751 <= b(31) and w11274;
w21752 <= b(29) and w11639;
w21753 <= b(30) and w11269;
w21754 <= not w21752 and not w21753;
w21755 <= not w21751 and w21754;
w21756 <= w3539 and w11277;
w21757 <= w21755 and not w21756;
w21758 <= a(59) and not w21757;
w21759 <= a(59) and not w21758;
w21760 <= not w21757 and not w21758;
w21761 <= not w21759 and not w21760;
w21762 <= w21750 and not w21761;
w21763 <= w21750 and not w21762;
w21764 <= not w21761 and not w21762;
w21765 <= not w21763 and not w21764;
w21766 <= not w21507 and not w21511;
w21767 <= w21765 and w21766;
w21768 <= not w21765 and not w21766;
w21769 <= not w21767 and not w21768;
w21770 <= b(34) and w10169;
w21771 <= b(32) and w10539;
w21772 <= b(33) and w10164;
w21773 <= not w21771 and not w21772;
w21774 <= not w21770 and w21773;
w21775 <= w4209 and w10172;
w21776 <= w21774 and not w21775;
w21777 <= a(56) and not w21776;
w21778 <= a(56) and not w21777;
w21779 <= not w21776 and not w21777;
w21780 <= not w21778 and not w21779;
w21781 <= w21769 and not w21780;
w21782 <= w21769 and not w21781;
w21783 <= not w21780 and not w21781;
w21784 <= not w21782 and not w21783;
w21785 <= not w21525 and not w21528;
w21786 <= w21784 and w21785;
w21787 <= not w21784 and not w21785;
w21788 <= not w21786 and not w21787;
w21789 <= b(37) and w9082;
w21790 <= b(35) and w9475;
w21791 <= b(36) and w9077;
w21792 <= not w21790 and not w21791;
w21793 <= not w21789 and w21792;
w21794 <= w4924 and w9085;
w21795 <= w21793 and not w21794;
w21796 <= a(53) and not w21795;
w21797 <= a(53) and not w21796;
w21798 <= not w21795 and not w21796;
w21799 <= not w21797 and not w21798;
w21800 <= not w21788 and w21799;
w21801 <= w21788 and not w21799;
w21802 <= not w21800 and not w21801;
w21803 <= not w21724 and w21802;
w21804 <= not w21724 and not w21803;
w21805 <= w21802 and not w21803;
w21806 <= not w21804 and not w21805;
w21807 <= not w21723 and not w21806;
w21808 <= w21723 and not w21805;
w21809 <= not w21804 and w21808;
w21810 <= not w21807 and not w21809;
w21811 <= not w21712 and w21810;
w21812 <= w21712 and not w21810;
w21813 <= not w21811 and not w21812;
w21814 <= not w21711 and w21813;
w21815 <= w21813 and not w21814;
w21816 <= not w21711 and not w21814;
w21817 <= not w21815 and not w21816;
w21818 <= not w21455 and not w21572;
w21819 <= not w21569 and not w21818;
w21820 <= w21817 and w21819;
w21821 <= not w21817 and not w21819;
w21822 <= not w21820 and not w21821;
w21823 <= b(46) and w6338;
w21824 <= b(44) and w6645;
w21825 <= b(45) and w6333;
w21826 <= not w21824 and not w21825;
w21827 <= not w21823 and w21826;
w21828 <= w6341 and w7420;
w21829 <= w21827 and not w21828;
w21830 <= a(44) and not w21829;
w21831 <= a(44) and not w21830;
w21832 <= not w21829 and not w21830;
w21833 <= not w21831 and not w21832;
w21834 <= w21822 and not w21833;
w21835 <= w21822 and not w21834;
w21836 <= not w21833 and not w21834;
w21837 <= not w21835 and not w21836;
w21838 <= not w21587 and not w21591;
w21839 <= w21837 and w21838;
w21840 <= not w21837 and not w21838;
w21841 <= not w21839 and not w21840;
w21842 <= b(49) and w5520;
w21843 <= b(47) and w5802;
w21844 <= b(48) and w5515;
w21845 <= not w21843 and not w21844;
w21846 <= not w21842 and w21845;
w21847 <= w5523 and w8368;
w21848 <= w21846 and not w21847;
w21849 <= a(41) and not w21848;
w21850 <= a(41) and not w21849;
w21851 <= not w21848 and not w21849;
w21852 <= not w21850 and not w21851;
w21853 <= w21841 and not w21852;
w21854 <= w21841 and not w21853;
w21855 <= not w21852 and not w21853;
w21856 <= not w21854 and not w21855;
w21857 <= not w21604 and not w21610;
w21858 <= w21856 and w21857;
w21859 <= not w21856 and not w21857;
w21860 <= not w21858 and not w21859;
w21861 <= b(52) and w4778;
w21862 <= b(50) and w5020;
w21863 <= b(51) and w4773;
w21864 <= not w21862 and not w21863;
w21865 <= not w21861 and w21864;
w21866 <= w4781 and w9371;
w21867 <= w21865 and not w21866;
w21868 <= a(38) and not w21867;
w21869 <= a(38) and not w21868;
w21870 <= not w21867 and not w21868;
w21871 <= not w21869 and not w21870;
w21872 <= w21860 and not w21871;
w21873 <= w21860 and not w21872;
w21874 <= not w21871 and not w21872;
w21875 <= not w21873 and not w21874;
w21876 <= not w21628 and w21875;
w21877 <= w21628 and not w21875;
w21878 <= not w21876 and not w21877;
w21879 <= b(55) and w4030;
w21880 <= b(53) and w4275;
w21881 <= b(54) and w4025;
w21882 <= not w21880 and not w21881;
w21883 <= not w21879 and w21882;
w21884 <= w4033 and w10427;
w21885 <= w21883 and not w21884;
w21886 <= a(35) and not w21885;
w21887 <= a(35) and not w21886;
w21888 <= not w21885 and not w21886;
w21889 <= not w21887 and not w21888;
w21890 <= not w21878 and not w21889;
w21891 <= w21878 and w21889;
w21892 <= not w21890 and not w21891;
w21893 <= w21700 and w21892;
w21894 <= not w21700 and not w21892;
w21895 <= not w21893 and not w21894;
w21896 <= not w21685 and w21895;
w21897 <= not w21685 and not w21896;
w21898 <= w21895 and not w21896;
w21899 <= not w21897 and not w21898;
w21900 <= not w21421 and not w21432;
w21901 <= not w21651 and not w21900;
w21902 <= b(62) and w2428;
w21903 <= b(63) and w2277;
w21904 <= not w21902 and not w21903;
w21905 <= not w2285 and w21904;
w21906 <= w13543 and w21904;
w21907 <= not w21905 and not w21906;
w21908 <= a(26) and not w21907;
w21909 <= not a(26) and w21907;
w21910 <= not w21908 and not w21909;
w21911 <= not w21901 and not w21910;
w21912 <= not w21901 and not w21911;
w21913 <= not w21910 and not w21911;
w21914 <= not w21912 and not w21913;
w21915 <= not w21899 and not w21914;
w21916 <= w21899 and not w21913;
w21917 <= not w21912 and w21916;
w21918 <= not w21915 and not w21917;
w21919 <= not w21669 and w21918;
w21920 <= not w21669 and not w21919;
w21921 <= w21918 and not w21919;
w21922 <= not w21920 and not w21921;
w21923 <= not w21667 and not w21922;
w21924 <= w21667 and not w21921;
w21925 <= not w21920 and w21924;
w21926 <= not w21923 and not w21925;
w21927 <= not w21919 and not w21923;
w21928 <= not w21911 and not w21915;
w21929 <= not w21682 and not w21896;
w21930 <= b(63) and w2428;
w21931 <= w2285 and w13540;
w21932 <= not w21930 and not w21931;
w21933 <= a(26) and not w21932;
w21934 <= a(26) and not w21933;
w21935 <= not w21932 and not w21933;
w21936 <= not w21934 and not w21935;
w21937 <= not w21929 and not w21936;
w21938 <= not w21929 and not w21937;
w21939 <= not w21936 and not w21937;
w21940 <= not w21938 and not w21939;
w21941 <= b(62) and w2793;
w21942 <= b(60) and w2986;
w21943 <= b(61) and w2788;
w21944 <= not w21942 and not w21943;
w21945 <= not w21941 and w21944;
w21946 <= w2796 and w13113;
w21947 <= w21945 and not w21946;
w21948 <= a(29) and not w21947;
w21949 <= a(29) and not w21948;
w21950 <= not w21947 and not w21948;
w21951 <= not w21949 and not w21950;
w21952 <= not w21698 and not w21893;
w21953 <= w21951 and w21952;
w21954 <= not w21951 and not w21952;
w21955 <= not w21953 and not w21954;
w21956 <= b(59) and w3381;
w21957 <= b(57) and w3586;
w21958 <= b(58) and w3376;
w21959 <= not w21957 and not w21958;
w21960 <= not w21956 and w21959;
w21961 <= w3384 and w11922;
w21962 <= w21960 and not w21961;
w21963 <= a(32) and not w21962;
w21964 <= a(32) and not w21963;
w21965 <= not w21962 and not w21963;
w21966 <= not w21964 and not w21965;
w21967 <= not w21628 and not w21875;
w21968 <= not w21890 and not w21967;
w21969 <= w21966 and w21968;
w21970 <= not w21966 and not w21968;
w21971 <= not w21969 and not w21970;
w21972 <= b(56) and w4030;
w21973 <= b(54) and w4275;
w21974 <= b(55) and w4025;
w21975 <= not w21973 and not w21974;
w21976 <= not w21972 and w21975;
w21977 <= w4033 and w10451;
w21978 <= w21976 and not w21977;
w21979 <= a(35) and not w21978;
w21980 <= a(35) and not w21979;
w21981 <= not w21978 and not w21979;
w21982 <= not w21980 and not w21981;
w21983 <= not w21859 and not w21872;
w21984 <= b(53) and w4778;
w21985 <= b(51) and w5020;
w21986 <= b(52) and w4773;
w21987 <= not w21985 and not w21986;
w21988 <= not w21984 and w21987;
w21989 <= w4781 and w9715;
w21990 <= w21988 and not w21989;
w21991 <= a(38) and not w21990;
w21992 <= a(38) and not w21991;
w21993 <= not w21990 and not w21991;
w21994 <= not w21992 and not w21993;
w21995 <= not w21840 and not w21853;
w21996 <= not w21811 and not w21814;
w21997 <= b(44) and w7189;
w21998 <= b(42) and w7530;
w21999 <= b(43) and w7184;
w22000 <= not w21998 and not w21999;
w22001 <= not w21997 and w22000;
w22002 <= w6815 and w7192;
w22003 <= w22001 and not w22002;
w22004 <= a(47) and not w22003;
w22005 <= a(47) and not w22004;
w22006 <= not w22003 and not w22004;
w22007 <= not w22005 and not w22006;
w22008 <= not w21803 and not w21807;
w22009 <= not w21768 and not w21781;
w22010 <= b(35) and w10169;
w22011 <= b(33) and w10539;
w22012 <= b(34) and w10164;
w22013 <= not w22011 and not w22012;
w22014 <= not w22010 and w22013;
w22015 <= w4439 and w10172;
w22016 <= w22014 and not w22015;
w22017 <= a(56) and not w22016;
w22018 <= a(56) and not w22017;
w22019 <= not w22016 and not w22017;
w22020 <= not w22018 and not w22019;
w22021 <= not w21748 and not w21762;
w22022 <= b(32) and w11274;
w22023 <= b(30) and w11639;
w22024 <= b(31) and w11269;
w22025 <= not w22023 and not w22024;
w22026 <= not w22022 and w22025;
w22027 <= w3756 and w11277;
w22028 <= w22026 and not w22027;
w22029 <= a(59) and not w22028;
w22030 <= a(59) and not w22029;
w22031 <= not w22028 and not w22029;
w22032 <= not w22030 and not w22031;
w22033 <= not w21732 and not w21745;
w22034 <= b(25) and w13646;
w22035 <= b(26) and not w13231;
w22036 <= not w22034 and not w22035;
w22037 <= not w21729 and w22036;
w22038 <= w21729 and not w22036;
w22039 <= not w22037 and not w22038;
w22040 <= b(29) and w12411;
w22041 <= b(27) and w12790;
w22042 <= b(28) and w12406;
w22043 <= not w22041 and not w22042;
w22044 <= not w22040 and w22043;
w22045 <= not w12414 and w22044;
w22046 <= not w3126 and w22044;
w22047 <= not w22045 and not w22046;
w22048 <= a(62) and not w22047;
w22049 <= not a(62) and w22047;
w22050 <= not w22048 and not w22049;
w22051 <= w22039 and not w22050;
w22052 <= not w22039 and w22050;
w22053 <= not w22051 and not w22052;
w22054 <= not w22033 and w22053;
w22055 <= w22033 and not w22053;
w22056 <= not w22054 and not w22055;
w22057 <= not w22032 and w22056;
w22058 <= w22032 and not w22056;
w22059 <= not w22057 and not w22058;
w22060 <= not w22021 and w22059;
w22061 <= w22021 and not w22059;
w22062 <= not w22060 and not w22061;
w22063 <= not w22020 and w22062;
w22064 <= w22020 and not w22062;
w22065 <= not w22063 and not w22064;
w22066 <= not w22009 and w22065;
w22067 <= w22009 and not w22065;
w22068 <= not w22066 and not w22067;
w22069 <= b(38) and w9082;
w22070 <= b(36) and w9475;
w22071 <= b(37) and w9077;
w22072 <= not w22070 and not w22071;
w22073 <= not w22069 and w22072;
w22074 <= w4948 and w9085;
w22075 <= w22073 and not w22074;
w22076 <= a(53) and not w22075;
w22077 <= a(53) and not w22076;
w22078 <= not w22075 and not w22076;
w22079 <= not w22077 and not w22078;
w22080 <= w22068 and not w22079;
w22081 <= w22068 and not w22080;
w22082 <= not w22079 and not w22080;
w22083 <= not w22081 and not w22082;
w22084 <= not w21787 and not w21801;
w22085 <= not w22083 and not w22084;
w22086 <= not w22083 and not w22085;
w22087 <= not w22084 and not w22085;
w22088 <= not w22086 and not w22087;
w22089 <= b(41) and w8105;
w22090 <= b(39) and w8458;
w22091 <= b(40) and w8100;
w22092 <= not w22090 and not w22091;
w22093 <= not w22089 and w22092;
w22094 <= w5962 and w8108;
w22095 <= w22093 and not w22094;
w22096 <= a(50) and not w22095;
w22097 <= a(50) and not w22096;
w22098 <= not w22095 and not w22096;
w22099 <= not w22097 and not w22098;
w22100 <= not w22088 and w22099;
w22101 <= w22088 and not w22099;
w22102 <= not w22100 and not w22101;
w22103 <= not w22008 and not w22102;
w22104 <= w22008 and w22102;
w22105 <= not w22103 and not w22104;
w22106 <= not w22007 and w22105;
w22107 <= w22007 and not w22105;
w22108 <= not w22106 and not w22107;
w22109 <= not w21996 and w22108;
w22110 <= w21996 and not w22108;
w22111 <= not w22109 and not w22110;
w22112 <= b(47) and w6338;
w22113 <= b(45) and w6645;
w22114 <= b(46) and w6333;
w22115 <= not w22113 and not w22114;
w22116 <= not w22112 and w22115;
w22117 <= w6341 and w7446;
w22118 <= w22116 and not w22117;
w22119 <= a(44) and not w22118;
w22120 <= a(44) and not w22119;
w22121 <= not w22118 and not w22119;
w22122 <= not w22120 and not w22121;
w22123 <= w22111 and not w22122;
w22124 <= w22111 and not w22123;
w22125 <= not w22122 and not w22123;
w22126 <= not w22124 and not w22125;
w22127 <= not w21821 and not w21834;
w22128 <= w22126 and w22127;
w22129 <= not w22126 and not w22127;
w22130 <= not w22128 and not w22129;
w22131 <= b(50) and w5520;
w22132 <= b(48) and w5802;
w22133 <= b(49) and w5515;
w22134 <= not w22132 and not w22133;
w22135 <= not w22131 and w22134;
w22136 <= w5523 and w8692;
w22137 <= w22135 and not w22136;
w22138 <= a(41) and not w22137;
w22139 <= a(41) and not w22138;
w22140 <= not w22137 and not w22138;
w22141 <= not w22139 and not w22140;
w22142 <= not w22130 and w22141;
w22143 <= w22130 and not w22141;
w22144 <= not w22142 and not w22143;
w22145 <= not w21995 and w22144;
w22146 <= not w21995 and not w22145;
w22147 <= w22144 and not w22145;
w22148 <= not w22146 and not w22147;
w22149 <= not w21994 and not w22148;
w22150 <= w21994 and not w22147;
w22151 <= not w22146 and w22150;
w22152 <= not w22149 and not w22151;
w22153 <= not w21983 and w22152;
w22154 <= w21983 and not w22152;
w22155 <= not w22153 and not w22154;
w22156 <= not w21982 and w22155;
w22157 <= not w21982 and not w22156;
w22158 <= w22155 and not w22156;
w22159 <= not w22157 and not w22158;
w22160 <= w21971 and not w22159;
w22161 <= w21971 and not w22160;
w22162 <= not w22159 and not w22160;
w22163 <= not w22161 and not w22162;
w22164 <= not w21955 and w22163;
w22165 <= w21955 and not w22163;
w22166 <= not w22164 and not w22165;
w22167 <= not w21940 and w22166;
w22168 <= w21940 and not w22166;
w22169 <= not w22167 and not w22168;
w22170 <= not w21928 and w22169;
w22171 <= w21928 and not w22169;
w22172 <= not w22170 and not w22171;
w22173 <= not w21927 and w22172;
w22174 <= w21927 and not w22172;
w22175 <= not w22173 and not w22174;
w22176 <= not w21937 and not w22167;
w22177 <= not w21954 and not w22165;
w22178 <= b(63) and w2793;
w22179 <= b(61) and w2986;
w22180 <= b(62) and w2788;
w22181 <= not w22179 and not w22180;
w22182 <= not w22178 and w22181;
w22183 <= w2796 and w13514;
w22184 <= w22182 and not w22183;
w22185 <= a(29) and not w22184;
w22186 <= a(29) and not w22185;
w22187 <= not w22184 and not w22185;
w22188 <= not w22186 and not w22187;
w22189 <= not w22177 and not w22188;
w22190 <= not w22177 and not w22189;
w22191 <= not w22188 and not w22189;
w22192 <= not w22190 and not w22191;
w22193 <= b(57) and w4030;
w22194 <= b(55) and w4275;
w22195 <= b(56) and w4025;
w22196 <= not w22194 and not w22195;
w22197 <= not w22193 and w22196;
w22198 <= w4033 and w11153;
w22199 <= w22197 and not w22198;
w22200 <= a(35) and not w22199;
w22201 <= a(35) and not w22200;
w22202 <= not w22199 and not w22200;
w22203 <= not w22201 and not w22202;
w22204 <= not w22145 and not w22149;
w22205 <= not w22129 and not w22143;
w22206 <= not w22103 and not w22106;
w22207 <= not w22088 and not w22099;
w22208 <= not w22085 and not w22207;
w22209 <= b(33) and w11274;
w22210 <= b(31) and w11639;
w22211 <= b(32) and w11269;
w22212 <= not w22210 and not w22211;
w22213 <= not w22209 and w22212;
w22214 <= w3966 and w11277;
w22215 <= w22213 and not w22214;
w22216 <= a(59) and not w22215;
w22217 <= a(59) and not w22216;
w22218 <= not w22215 and not w22216;
w22219 <= not w22217 and not w22218;
w22220 <= not w22054 and not w22057;
w22221 <= w22219 and w22220;
w22222 <= not w22219 and not w22220;
w22223 <= not w22221 and not w22222;
w22224 <= not w22037 and not w22051;
w22225 <= b(26) and w13646;
w22226 <= b(27) and not w13231;
w22227 <= not w22225 and not w22226;
w22228 <= not a(26) and not w22227;
w22229 <= a(26) and w22227;
w22230 <= not w22228 and not w22229;
w22231 <= not w22036 and w22230;
w22232 <= w22036 and not w22230;
w22233 <= not w22231 and not w22232;
w22234 <= not w22224 and w22233;
w22235 <= w22224 and not w22233;
w22236 <= not w22234 and not w22235;
w22237 <= b(30) and w12411;
w22238 <= b(28) and w12790;
w22239 <= b(29) and w12406;
w22240 <= not w22238 and not w22239;
w22241 <= not w22237 and w22240;
w22242 <= w3320 and w12414;
w22243 <= w22241 and not w22242;
w22244 <= a(62) and not w22243;
w22245 <= a(62) and not w22244;
w22246 <= not w22243 and not w22244;
w22247 <= not w22245 and not w22246;
w22248 <= w22236 and not w22247;
w22249 <= w22236 and not w22248;
w22250 <= not w22247 and not w22248;
w22251 <= not w22249 and not w22250;
w22252 <= not w22223 and w22251;
w22253 <= w22223 and not w22251;
w22254 <= not w22252 and not w22253;
w22255 <= b(36) and w10169;
w22256 <= b(34) and w10539;
w22257 <= b(35) and w10164;
w22258 <= not w22256 and not w22257;
w22259 <= not w22255 and w22258;
w22260 <= w4665 and w10172;
w22261 <= w22259 and not w22260;
w22262 <= a(56) and not w22261;
w22263 <= a(56) and not w22262;
w22264 <= not w22261 and not w22262;
w22265 <= not w22263 and not w22264;
w22266 <= w22254 and not w22265;
w22267 <= w22254 and not w22266;
w22268 <= not w22265 and not w22266;
w22269 <= not w22267 and not w22268;
w22270 <= not w22060 and not w22063;
w22271 <= w22269 and w22270;
w22272 <= not w22269 and not w22270;
w22273 <= not w22271 and not w22272;
w22274 <= b(39) and w9082;
w22275 <= b(37) and w9475;
w22276 <= b(38) and w9077;
w22277 <= not w22275 and not w22276;
w22278 <= not w22274 and w22277;
w22279 <= w5194 and w9085;
w22280 <= w22278 and not w22279;
w22281 <= a(53) and not w22280;
w22282 <= a(53) and not w22281;
w22283 <= not w22280 and not w22281;
w22284 <= not w22282 and not w22283;
w22285 <= w22273 and not w22284;
w22286 <= w22273 and not w22285;
w22287 <= not w22284 and not w22285;
w22288 <= not w22286 and not w22287;
w22289 <= not w22066 and not w22080;
w22290 <= w22288 and w22289;
w22291 <= not w22288 and not w22289;
w22292 <= not w22290 and not w22291;
w22293 <= b(42) and w8105;
w22294 <= b(40) and w8458;
w22295 <= b(41) and w8100;
w22296 <= not w22294 and not w22295;
w22297 <= not w22293 and w22296;
w22298 <= w6232 and w8108;
w22299 <= w22297 and not w22298;
w22300 <= a(50) and not w22299;
w22301 <= a(50) and not w22300;
w22302 <= not w22299 and not w22300;
w22303 <= not w22301 and not w22302;
w22304 <= w22292 and not w22303;
w22305 <= w22292 and not w22304;
w22306 <= not w22303 and not w22304;
w22307 <= not w22305 and not w22306;
w22308 <= not w22208 and w22307;
w22309 <= w22208 and not w22307;
w22310 <= not w22308 and not w22309;
w22311 <= b(45) and w7189;
w22312 <= b(43) and w7530;
w22313 <= b(44) and w7184;
w22314 <= not w22312 and not w22313;
w22315 <= not w22311 and w22314;
w22316 <= w7104 and w7192;
w22317 <= w22315 and not w22316;
w22318 <= a(47) and not w22317;
w22319 <= a(47) and not w22318;
w22320 <= not w22317 and not w22318;
w22321 <= not w22319 and not w22320;
w22322 <= not w22310 and not w22321;
w22323 <= w22310 and w22321;
w22324 <= not w22322 and not w22323;
w22325 <= w22206 and not w22324;
w22326 <= not w22206 and w22324;
w22327 <= not w22325 and not w22326;
w22328 <= b(48) and w6338;
w22329 <= b(46) and w6645;
w22330 <= b(47) and w6333;
w22331 <= not w22329 and not w22330;
w22332 <= not w22328 and w22331;
w22333 <= w6341 and w7752;
w22334 <= w22332 and not w22333;
w22335 <= a(44) and not w22334;
w22336 <= a(44) and not w22335;
w22337 <= not w22334 and not w22335;
w22338 <= not w22336 and not w22337;
w22339 <= w22327 and not w22338;
w22340 <= w22327 and not w22339;
w22341 <= not w22338 and not w22339;
w22342 <= not w22340 and not w22341;
w22343 <= not w22109 and not w22123;
w22344 <= w22342 and w22343;
w22345 <= not w22342 and not w22343;
w22346 <= not w22344 and not w22345;
w22347 <= b(51) and w5520;
w22348 <= b(49) and w5802;
w22349 <= b(50) and w5515;
w22350 <= not w22348 and not w22349;
w22351 <= not w22347 and w22350;
w22352 <= w5523 and w8719;
w22353 <= w22351 and not w22352;
w22354 <= a(41) and not w22353;
w22355 <= a(41) and not w22354;
w22356 <= not w22353 and not w22354;
w22357 <= not w22355 and not w22356;
w22358 <= w22346 and not w22357;
w22359 <= not w22346 and w22357;
w22360 <= not w22205 and not w22359;
w22361 <= not w22358 and w22360;
w22362 <= not w22205 and not w22361;
w22363 <= not w22358 and not w22361;
w22364 <= not w22359 and w22363;
w22365 <= not w22362 and not w22364;
w22366 <= b(54) and w4778;
w22367 <= b(52) and w5020;
w22368 <= b(53) and w4773;
w22369 <= not w22367 and not w22368;
w22370 <= not w22366 and w22369;
w22371 <= w4781 and w9741;
w22372 <= w22370 and not w22371;
w22373 <= a(38) and not w22372;
w22374 <= a(38) and not w22373;
w22375 <= not w22372 and not w22373;
w22376 <= not w22374 and not w22375;
w22377 <= w22365 and w22376;
w22378 <= not w22365 and not w22376;
w22379 <= not w22377 and not w22378;
w22380 <= not w22204 and w22379;
w22381 <= w22204 and not w22379;
w22382 <= not w22380 and not w22381;
w22383 <= not w22203 and w22382;
w22384 <= w22382 and not w22383;
w22385 <= not w22203 and not w22383;
w22386 <= not w22384 and not w22385;
w22387 <= not w22153 and not w22156;
w22388 <= w22386 and w22387;
w22389 <= not w22386 and not w22387;
w22390 <= not w22388 and not w22389;
w22391 <= b(60) and w3381;
w22392 <= b(58) and w3586;
w22393 <= b(59) and w3376;
w22394 <= not w22392 and not w22393;
w22395 <= not w22391 and w22394;
w22396 <= w3384 and w11954;
w22397 <= w22395 and not w22396;
w22398 <= a(32) and not w22397;
w22399 <= a(32) and not w22398;
w22400 <= not w22397 and not w22398;
w22401 <= not w22399 and not w22400;
w22402 <= not w21970 and not w22160;
w22403 <= w22401 and w22402;
w22404 <= not w22401 and not w22402;
w22405 <= not w22403 and not w22404;
w22406 <= w22390 and not w22405;
w22407 <= not w22390 and w22405;
w22408 <= not w22406 and not w22407;
w22409 <= not w22192 and not w22408;
w22410 <= w22192 and w22408;
w22411 <= not w22409 and not w22410;
w22412 <= w22176 and not w22411;
w22413 <= not w22176 and w22411;
w22414 <= not w22412 and not w22413;
w22415 <= not w22170 and not w22173;
w22416 <= w22414 and not w22415;
w22417 <= not w22414 and w22415;
w22418 <= not w22416 and not w22417;
w22419 <= w22390 and w22405;
w22420 <= not w22404 and not w22419;
w22421 <= b(62) and w2986;
w22422 <= b(63) and w2788;
w22423 <= not w22421 and not w22422;
w22424 <= not w2796 and w22423;
w22425 <= w13543 and w22423;
w22426 <= not w22424 and not w22425;
w22427 <= a(29) and not w22426;
w22428 <= not a(29) and w22426;
w22429 <= not w22427 and not w22428;
w22430 <= not w22420 and not w22429;
w22431 <= w22420 and w22429;
w22432 <= not w22430 and not w22431;
w22433 <= b(61) and w3381;
w22434 <= b(59) and w3586;
w22435 <= b(60) and w3376;
w22436 <= not w22434 and not w22435;
w22437 <= not w22433 and w22436;
w22438 <= w3384 and w12712;
w22439 <= w22437 and not w22438;
w22440 <= a(32) and not w22439;
w22441 <= a(32) and not w22440;
w22442 <= not w22439 and not w22440;
w22443 <= not w22441 and not w22442;
w22444 <= not w22383 and not w22389;
w22445 <= w22443 and w22444;
w22446 <= not w22443 and not w22444;
w22447 <= not w22445 and not w22446;
w22448 <= b(58) and w4030;
w22449 <= b(56) and w4275;
w22450 <= b(57) and w4025;
w22451 <= not w22449 and not w22450;
w22452 <= not w22448 and w22451;
w22453 <= w4033 and w11179;
w22454 <= w22452 and not w22453;
w22455 <= a(35) and not w22454;
w22456 <= a(35) and not w22455;
w22457 <= not w22454 and not w22455;
w22458 <= not w22456 and not w22457;
w22459 <= not w22378 and not w22380;
w22460 <= b(43) and w8105;
w22461 <= b(41) and w8458;
w22462 <= b(42) and w8100;
w22463 <= not w22461 and not w22462;
w22464 <= not w22460 and w22463;
w22465 <= w6258 and w8108;
w22466 <= w22464 and not w22465;
w22467 <= a(50) and not w22466;
w22468 <= a(50) and not w22467;
w22469 <= not w22466 and not w22467;
w22470 <= not w22468 and not w22469;
w22471 <= not w22285 and not w22291;
w22472 <= b(40) and w9082;
w22473 <= b(38) and w9475;
w22474 <= b(39) and w9077;
w22475 <= not w22473 and not w22474;
w22476 <= not w22472 and w22475;
w22477 <= w5698 and w9085;
w22478 <= w22476 and not w22477;
w22479 <= a(53) and not w22478;
w22480 <= a(53) and not w22479;
w22481 <= not w22478 and not w22479;
w22482 <= not w22480 and not w22481;
w22483 <= not w22266 and not w22272;
w22484 <= b(34) and w11274;
w22485 <= b(32) and w11639;
w22486 <= b(33) and w11269;
w22487 <= not w22485 and not w22486;
w22488 <= not w22484 and w22487;
w22489 <= w4209 and w11277;
w22490 <= w22488 and not w22489;
w22491 <= a(59) and not w22490;
w22492 <= a(59) and not w22491;
w22493 <= not w22490 and not w22491;
w22494 <= not w22492 and not w22493;
w22495 <= b(27) and w13646;
w22496 <= b(28) and not w13231;
w22497 <= not w22495 and not w22496;
w22498 <= not w22228 and not w22231;
w22499 <= not w22497 and w22498;
w22500 <= w22497 and not w22498;
w22501 <= not w22499 and not w22500;
w22502 <= b(31) and w12411;
w22503 <= b(29) and w12790;
w22504 <= b(30) and w12406;
w22505 <= not w22503 and not w22504;
w22506 <= not w22502 and w22505;
w22507 <= w3539 and w12414;
w22508 <= w22506 and not w22507;
w22509 <= a(62) and not w22508;
w22510 <= a(62) and not w22509;
w22511 <= not w22508 and not w22509;
w22512 <= not w22510 and not w22511;
w22513 <= not w22501 and w22512;
w22514 <= w22501 and not w22512;
w22515 <= not w22513 and not w22514;
w22516 <= not w22234 and not w22248;
w22517 <= w22515 and not w22516;
w22518 <= not w22515 and w22516;
w22519 <= not w22517 and not w22518;
w22520 <= not w22494 and w22519;
w22521 <= w22519 and not w22520;
w22522 <= not w22494 and not w22520;
w22523 <= not w22521 and not w22522;
w22524 <= not w22222 and not w22253;
w22525 <= not w22523 and not w22524;
w22526 <= not w22523 and not w22525;
w22527 <= not w22524 and not w22525;
w22528 <= not w22526 and not w22527;
w22529 <= b(37) and w10169;
w22530 <= b(35) and w10539;
w22531 <= b(36) and w10164;
w22532 <= not w22530 and not w22531;
w22533 <= not w22529 and w22532;
w22534 <= w4924 and w10172;
w22535 <= w22533 and not w22534;
w22536 <= a(56) and not w22535;
w22537 <= a(56) and not w22536;
w22538 <= not w22535 and not w22536;
w22539 <= not w22537 and not w22538;
w22540 <= not w22528 and w22539;
w22541 <= w22528 and not w22539;
w22542 <= not w22540 and not w22541;
w22543 <= not w22483 and not w22542;
w22544 <= not w22483 and not w22543;
w22545 <= not w22542 and not w22543;
w22546 <= not w22544 and not w22545;
w22547 <= not w22482 and not w22546;
w22548 <= w22482 and not w22545;
w22549 <= not w22544 and w22548;
w22550 <= not w22547 and not w22549;
w22551 <= not w22471 and w22550;
w22552 <= w22471 and not w22550;
w22553 <= not w22551 and not w22552;
w22554 <= not w22470 and w22553;
w22555 <= w22553 and not w22554;
w22556 <= not w22470 and not w22554;
w22557 <= not w22555 and not w22556;
w22558 <= not w22208 and not w22307;
w22559 <= not w22304 and not w22558;
w22560 <= w22557 and w22559;
w22561 <= not w22557 and not w22559;
w22562 <= not w22560 and not w22561;
w22563 <= b(46) and w7189;
w22564 <= b(44) and w7530;
w22565 <= b(45) and w7184;
w22566 <= not w22564 and not w22565;
w22567 <= not w22563 and w22566;
w22568 <= w7192 and w7420;
w22569 <= w22567 and not w22568;
w22570 <= a(47) and not w22569;
w22571 <= a(47) and not w22570;
w22572 <= not w22569 and not w22570;
w22573 <= not w22571 and not w22572;
w22574 <= w22562 and not w22573;
w22575 <= w22562 and not w22574;
w22576 <= not w22573 and not w22574;
w22577 <= not w22575 and not w22576;
w22578 <= not w22322 and not w22326;
w22579 <= w22577 and w22578;
w22580 <= not w22577 and not w22578;
w22581 <= not w22579 and not w22580;
w22582 <= b(49) and w6338;
w22583 <= b(47) and w6645;
w22584 <= b(48) and w6333;
w22585 <= not w22583 and not w22584;
w22586 <= not w22582 and w22585;
w22587 <= w6341 and w8368;
w22588 <= w22586 and not w22587;
w22589 <= a(44) and not w22588;
w22590 <= a(44) and not w22589;
w22591 <= not w22588 and not w22589;
w22592 <= not w22590 and not w22591;
w22593 <= w22581 and not w22592;
w22594 <= w22581 and not w22593;
w22595 <= not w22592 and not w22593;
w22596 <= not w22594 and not w22595;
w22597 <= not w22339 and not w22345;
w22598 <= w22596 and w22597;
w22599 <= not w22596 and not w22597;
w22600 <= not w22598 and not w22599;
w22601 <= b(52) and w5520;
w22602 <= b(50) and w5802;
w22603 <= b(51) and w5515;
w22604 <= not w22602 and not w22603;
w22605 <= not w22601 and w22604;
w22606 <= w5523 and w9371;
w22607 <= w22605 and not w22606;
w22608 <= a(41) and not w22607;
w22609 <= a(41) and not w22608;
w22610 <= not w22607 and not w22608;
w22611 <= not w22609 and not w22610;
w22612 <= w22600 and not w22611;
w22613 <= w22600 and not w22612;
w22614 <= not w22611 and not w22612;
w22615 <= not w22613 and not w22614;
w22616 <= not w22363 and w22615;
w22617 <= w22363 and not w22615;
w22618 <= not w22616 and not w22617;
w22619 <= b(55) and w4778;
w22620 <= b(53) and w5020;
w22621 <= b(54) and w4773;
w22622 <= not w22620 and not w22621;
w22623 <= not w22619 and w22622;
w22624 <= w4781 and w10427;
w22625 <= w22623 and not w22624;
w22626 <= a(38) and not w22625;
w22627 <= a(38) and not w22626;
w22628 <= not w22625 and not w22626;
w22629 <= not w22627 and not w22628;
w22630 <= not w22618 and not w22629;
w22631 <= w22618 and w22629;
w22632 <= not w22630 and not w22631;
w22633 <= not w22459 and w22632;
w22634 <= w22459 and not w22632;
w22635 <= not w22633 and not w22634;
w22636 <= not w22458 and w22635;
w22637 <= w22635 and not w22636;
w22638 <= not w22458 and not w22636;
w22639 <= not w22637 and not w22638;
w22640 <= w22447 and not w22639;
w22641 <= not w22447 and w22639;
w22642 <= w22432 and not w22641;
w22643 <= not w22640 and w22642;
w22644 <= w22432 and not w22643;
w22645 <= not w22641 and not w22643;
w22646 <= not w22640 and w22645;
w22647 <= not w22644 and not w22646;
w22648 <= not w22189 and not w22409;
w22649 <= w22647 and w22648;
w22650 <= not w22647 and not w22648;
w22651 <= not w22649 and not w22650;
w22652 <= not w22413 and not w22416;
w22653 <= w22651 and not w22652;
w22654 <= not w22651 and w22652;
w22655 <= not w22653 and not w22654;
w22656 <= not w22650 and not w22653;
w22657 <= not w22430 and not w22643;
w22658 <= not w22446 and not w22640;
w22659 <= b(63) and w2986;
w22660 <= w2796 and w13540;
w22661 <= not w22659 and not w22660;
w22662 <= a(29) and not w22661;
w22663 <= a(29) and not w22662;
w22664 <= not w22661 and not w22662;
w22665 <= not w22663 and not w22664;
w22666 <= not w22658 and not w22665;
w22667 <= not w22658 and not w22666;
w22668 <= not w22665 and not w22666;
w22669 <= not w22667 and not w22668;
w22670 <= b(62) and w3381;
w22671 <= b(60) and w3586;
w22672 <= b(61) and w3376;
w22673 <= not w22671 and not w22672;
w22674 <= not w22670 and w22673;
w22675 <= w3384 and w13113;
w22676 <= w22674 and not w22675;
w22677 <= a(32) and not w22676;
w22678 <= a(32) and not w22677;
w22679 <= not w22676 and not w22677;
w22680 <= not w22678 and not w22679;
w22681 <= not w22633 and not w22636;
w22682 <= w22680 and w22681;
w22683 <= not w22680 and not w22681;
w22684 <= not w22682 and not w22683;
w22685 <= not w22363 and not w22615;
w22686 <= not w22630 and not w22685;
w22687 <= b(56) and w4778;
w22688 <= b(54) and w5020;
w22689 <= b(55) and w4773;
w22690 <= not w22688 and not w22689;
w22691 <= not w22687 and w22690;
w22692 <= w4781 and w10451;
w22693 <= w22691 and not w22692;
w22694 <= a(38) and not w22693;
w22695 <= a(38) and not w22694;
w22696 <= not w22693 and not w22694;
w22697 <= not w22695 and not w22696;
w22698 <= not w22599 and not w22612;
w22699 <= b(53) and w5520;
w22700 <= b(51) and w5802;
w22701 <= b(52) and w5515;
w22702 <= not w22700 and not w22701;
w22703 <= not w22699 and w22702;
w22704 <= w5523 and w9715;
w22705 <= w22703 and not w22704;
w22706 <= a(41) and not w22705;
w22707 <= a(41) and not w22706;
w22708 <= not w22705 and not w22706;
w22709 <= not w22707 and not w22708;
w22710 <= not w22580 and not w22593;
w22711 <= not w22551 and not w22554;
w22712 <= b(44) and w8105;
w22713 <= b(42) and w8458;
w22714 <= b(43) and w8100;
w22715 <= not w22713 and not w22714;
w22716 <= not w22712 and w22715;
w22717 <= w6815 and w8108;
w22718 <= w22716 and not w22717;
w22719 <= a(50) and not w22718;
w22720 <= a(50) and not w22719;
w22721 <= not w22718 and not w22719;
w22722 <= not w22720 and not w22721;
w22723 <= not w22543 and not w22547;
w22724 <= not w22517 and not w22520;
w22725 <= b(35) and w11274;
w22726 <= b(33) and w11639;
w22727 <= b(34) and w11269;
w22728 <= not w22726 and not w22727;
w22729 <= not w22725 and w22728;
w22730 <= w4439 and w11277;
w22731 <= w22729 and not w22730;
w22732 <= a(59) and not w22731;
w22733 <= a(59) and not w22732;
w22734 <= not w22731 and not w22732;
w22735 <= not w22733 and not w22734;
w22736 <= not w22500 and not w22514;
w22737 <= b(28) and w13646;
w22738 <= b(29) and not w13231;
w22739 <= not w22737 and not w22738;
w22740 <= w22497 and not w22739;
w22741 <= not w22497 and w22739;
w22742 <= not w22736 and not w22741;
w22743 <= not w22740 and w22742;
w22744 <= not w22736 and not w22743;
w22745 <= not w22741 and not w22743;
w22746 <= not w22740 and w22745;
w22747 <= not w22744 and not w22746;
w22748 <= b(32) and w12411;
w22749 <= b(30) and w12790;
w22750 <= b(31) and w12406;
w22751 <= not w22749 and not w22750;
w22752 <= not w22748 and w22751;
w22753 <= w3756 and w12414;
w22754 <= w22752 and not w22753;
w22755 <= a(62) and not w22754;
w22756 <= a(62) and not w22755;
w22757 <= not w22754 and not w22755;
w22758 <= not w22756 and not w22757;
w22759 <= not w22747 and w22758;
w22760 <= w22747 and not w22758;
w22761 <= not w22759 and not w22760;
w22762 <= not w22735 and not w22761;
w22763 <= w22735 and w22761;
w22764 <= not w22762 and not w22763;
w22765 <= not w22724 and w22764;
w22766 <= w22724 and not w22764;
w22767 <= not w22765 and not w22766;
w22768 <= b(38) and w10169;
w22769 <= b(36) and w10539;
w22770 <= b(37) and w10164;
w22771 <= not w22769 and not w22770;
w22772 <= not w22768 and w22771;
w22773 <= w4948 and w10172;
w22774 <= w22772 and not w22773;
w22775 <= a(56) and not w22774;
w22776 <= a(56) and not w22775;
w22777 <= not w22774 and not w22775;
w22778 <= not w22776 and not w22777;
w22779 <= w22767 and not w22778;
w22780 <= w22767 and not w22779;
w22781 <= not w22778 and not w22779;
w22782 <= not w22780 and not w22781;
w22783 <= not w22528 and not w22539;
w22784 <= not w22525 and not w22783;
w22785 <= not w22782 and not w22784;
w22786 <= not w22782 and not w22785;
w22787 <= not w22784 and not w22785;
w22788 <= not w22786 and not w22787;
w22789 <= b(41) and w9082;
w22790 <= b(39) and w9475;
w22791 <= b(40) and w9077;
w22792 <= not w22790 and not w22791;
w22793 <= not w22789 and w22792;
w22794 <= w5962 and w9085;
w22795 <= w22793 and not w22794;
w22796 <= a(53) and not w22795;
w22797 <= a(53) and not w22796;
w22798 <= not w22795 and not w22796;
w22799 <= not w22797 and not w22798;
w22800 <= not w22788 and w22799;
w22801 <= w22788 and not w22799;
w22802 <= not w22800 and not w22801;
w22803 <= not w22723 and not w22802;
w22804 <= w22723 and w22802;
w22805 <= not w22803 and not w22804;
w22806 <= not w22722 and w22805;
w22807 <= w22722 and not w22805;
w22808 <= not w22806 and not w22807;
w22809 <= not w22711 and w22808;
w22810 <= w22711 and not w22808;
w22811 <= not w22809 and not w22810;
w22812 <= b(47) and w7189;
w22813 <= b(45) and w7530;
w22814 <= b(46) and w7184;
w22815 <= not w22813 and not w22814;
w22816 <= not w22812 and w22815;
w22817 <= w7192 and w7446;
w22818 <= w22816 and not w22817;
w22819 <= a(47) and not w22818;
w22820 <= a(47) and not w22819;
w22821 <= not w22818 and not w22819;
w22822 <= not w22820 and not w22821;
w22823 <= w22811 and not w22822;
w22824 <= w22811 and not w22823;
w22825 <= not w22822 and not w22823;
w22826 <= not w22824 and not w22825;
w22827 <= not w22561 and not w22574;
w22828 <= w22826 and w22827;
w22829 <= not w22826 and not w22827;
w22830 <= not w22828 and not w22829;
w22831 <= b(50) and w6338;
w22832 <= b(48) and w6645;
w22833 <= b(49) and w6333;
w22834 <= not w22832 and not w22833;
w22835 <= not w22831 and w22834;
w22836 <= w6341 and w8692;
w22837 <= w22835 and not w22836;
w22838 <= a(44) and not w22837;
w22839 <= a(44) and not w22838;
w22840 <= not w22837 and not w22838;
w22841 <= not w22839 and not w22840;
w22842 <= not w22830 and w22841;
w22843 <= w22830 and not w22841;
w22844 <= not w22842 and not w22843;
w22845 <= not w22710 and w22844;
w22846 <= not w22710 and not w22845;
w22847 <= w22844 and not w22845;
w22848 <= not w22846 and not w22847;
w22849 <= not w22709 and not w22848;
w22850 <= w22709 and not w22847;
w22851 <= not w22846 and w22850;
w22852 <= not w22849 and not w22851;
w22853 <= not w22698 and w22852;
w22854 <= w22698 and not w22852;
w22855 <= not w22853 and not w22854;
w22856 <= not w22697 and w22855;
w22857 <= w22697 and not w22855;
w22858 <= not w22856 and not w22857;
w22859 <= not w22686 and w22858;
w22860 <= w22686 and not w22858;
w22861 <= not w22859 and not w22860;
w22862 <= b(59) and w4030;
w22863 <= b(57) and w4275;
w22864 <= b(58) and w4025;
w22865 <= not w22863 and not w22864;
w22866 <= not w22862 and w22865;
w22867 <= w4033 and w11922;
w22868 <= w22866 and not w22867;
w22869 <= a(35) and not w22868;
w22870 <= a(35) and not w22869;
w22871 <= not w22868 and not w22869;
w22872 <= not w22870 and not w22871;
w22873 <= w22861 and not w22872;
w22874 <= w22861 and not w22873;
w22875 <= not w22872 and not w22873;
w22876 <= not w22874 and not w22875;
w22877 <= not w22684 and w22876;
w22878 <= w22684 and not w22876;
w22879 <= not w22877 and not w22878;
w22880 <= not w22669 and w22879;
w22881 <= w22669 and not w22879;
w22882 <= not w22880 and not w22881;
w22883 <= not w22657 and w22882;
w22884 <= not w22657 and not w22883;
w22885 <= w22882 and not w22883;
w22886 <= not w22884 and not w22885;
w22887 <= not w22656 and not w22886;
w22888 <= w22656 and not w22885;
w22889 <= not w22884 and w22888;
w22890 <= not w22887 and not w22889;
w22891 <= not w22883 and not w22887;
w22892 <= not w22666 and not w22880;
w22893 <= b(57) and w4778;
w22894 <= b(55) and w5020;
w22895 <= b(56) and w4773;
w22896 <= not w22894 and not w22895;
w22897 <= not w22893 and w22896;
w22898 <= w4781 and w11153;
w22899 <= w22897 and not w22898;
w22900 <= a(38) and not w22899;
w22901 <= a(38) and not w22900;
w22902 <= not w22899 and not w22900;
w22903 <= not w22901 and not w22902;
w22904 <= not w22845 and not w22849;
w22905 <= not w22829 and not w22843;
w22906 <= not w22803 and not w22806;
w22907 <= not w22788 and not w22799;
w22908 <= not w22785 and not w22907;
w22909 <= b(39) and w10169;
w22910 <= b(37) and w10539;
w22911 <= b(38) and w10164;
w22912 <= not w22910 and not w22911;
w22913 <= not w22909 and w22912;
w22914 <= w5194 and w10172;
w22915 <= w22913 and not w22914;
w22916 <= a(56) and not w22915;
w22917 <= a(56) and not w22916;
w22918 <= not w22915 and not w22916;
w22919 <= not w22917 and not w22918;
w22920 <= not w22747 and not w22758;
w22921 <= not w22762 and not w22920;
w22922 <= b(29) and w13646;
w22923 <= b(30) and not w13231;
w22924 <= not w22922 and not w22923;
w22925 <= not a(29) and not w22924;
w22926 <= a(29) and w22924;
w22927 <= not w22925 and not w22926;
w22928 <= not w22739 and w22927;
w22929 <= not w22739 and not w22928;
w22930 <= w22927 and not w22928;
w22931 <= not w22929 and not w22930;
w22932 <= not w22745 and not w22931;
w22933 <= not w22745 and not w22932;
w22934 <= not w22931 and not w22932;
w22935 <= not w22933 and not w22934;
w22936 <= b(33) and w12411;
w22937 <= b(31) and w12790;
w22938 <= b(32) and w12406;
w22939 <= not w22937 and not w22938;
w22940 <= not w22936 and w22939;
w22941 <= w3966 and w12414;
w22942 <= w22940 and not w22941;
w22943 <= a(62) and not w22942;
w22944 <= a(62) and not w22943;
w22945 <= not w22942 and not w22943;
w22946 <= not w22944 and not w22945;
w22947 <= not w22935 and w22946;
w22948 <= w22935 and not w22946;
w22949 <= not w22947 and not w22948;
w22950 <= b(36) and w11274;
w22951 <= b(34) and w11639;
w22952 <= b(35) and w11269;
w22953 <= not w22951 and not w22952;
w22954 <= not w22950 and w22953;
w22955 <= w4665 and w11277;
w22956 <= w22954 and not w22955;
w22957 <= a(59) and not w22956;
w22958 <= a(59) and not w22957;
w22959 <= not w22956 and not w22957;
w22960 <= not w22958 and not w22959;
w22961 <= not w22949 and not w22960;
w22962 <= w22949 and w22960;
w22963 <= not w22961 and not w22962;
w22964 <= not w22921 and w22963;
w22965 <= w22921 and not w22963;
w22966 <= not w22964 and not w22965;
w22967 <= not w22919 and w22966;
w22968 <= w22966 and not w22967;
w22969 <= not w22919 and not w22967;
w22970 <= not w22968 and not w22969;
w22971 <= not w22765 and not w22779;
w22972 <= w22970 and w22971;
w22973 <= not w22970 and not w22971;
w22974 <= not w22972 and not w22973;
w22975 <= b(42) and w9082;
w22976 <= b(40) and w9475;
w22977 <= b(41) and w9077;
w22978 <= not w22976 and not w22977;
w22979 <= not w22975 and w22978;
w22980 <= w6232 and w9085;
w22981 <= w22979 and not w22980;
w22982 <= a(53) and not w22981;
w22983 <= a(53) and not w22982;
w22984 <= not w22981 and not w22982;
w22985 <= not w22983 and not w22984;
w22986 <= w22974 and not w22985;
w22987 <= w22974 and not w22986;
w22988 <= not w22985 and not w22986;
w22989 <= not w22987 and not w22988;
w22990 <= not w22908 and w22989;
w22991 <= w22908 and not w22989;
w22992 <= not w22990 and not w22991;
w22993 <= b(45) and w8105;
w22994 <= b(43) and w8458;
w22995 <= b(44) and w8100;
w22996 <= not w22994 and not w22995;
w22997 <= not w22993 and w22996;
w22998 <= w7104 and w8108;
w22999 <= w22997 and not w22998;
w23000 <= a(50) and not w22999;
w23001 <= a(50) and not w23000;
w23002 <= not w22999 and not w23000;
w23003 <= not w23001 and not w23002;
w23004 <= not w22992 and not w23003;
w23005 <= w22992 and w23003;
w23006 <= not w23004 and not w23005;
w23007 <= w22906 and not w23006;
w23008 <= not w22906 and w23006;
w23009 <= not w23007 and not w23008;
w23010 <= b(48) and w7189;
w23011 <= b(46) and w7530;
w23012 <= b(47) and w7184;
w23013 <= not w23011 and not w23012;
w23014 <= not w23010 and w23013;
w23015 <= w7192 and w7752;
w23016 <= w23014 and not w23015;
w23017 <= a(47) and not w23016;
w23018 <= a(47) and not w23017;
w23019 <= not w23016 and not w23017;
w23020 <= not w23018 and not w23019;
w23021 <= w23009 and not w23020;
w23022 <= w23009 and not w23021;
w23023 <= not w23020 and not w23021;
w23024 <= not w23022 and not w23023;
w23025 <= not w22809 and not w22823;
w23026 <= w23024 and w23025;
w23027 <= not w23024 and not w23025;
w23028 <= not w23026 and not w23027;
w23029 <= b(51) and w6338;
w23030 <= b(49) and w6645;
w23031 <= b(50) and w6333;
w23032 <= not w23030 and not w23031;
w23033 <= not w23029 and w23032;
w23034 <= w6341 and w8719;
w23035 <= w23033 and not w23034;
w23036 <= a(44) and not w23035;
w23037 <= a(44) and not w23036;
w23038 <= not w23035 and not w23036;
w23039 <= not w23037 and not w23038;
w23040 <= w23028 and not w23039;
w23041 <= not w23028 and w23039;
w23042 <= not w22905 and not w23041;
w23043 <= not w23040 and w23042;
w23044 <= not w22905 and not w23043;
w23045 <= not w23040 and not w23043;
w23046 <= not w23041 and w23045;
w23047 <= not w23044 and not w23046;
w23048 <= b(54) and w5520;
w23049 <= b(52) and w5802;
w23050 <= b(53) and w5515;
w23051 <= not w23049 and not w23050;
w23052 <= not w23048 and w23051;
w23053 <= w5523 and w9741;
w23054 <= w23052 and not w23053;
w23055 <= a(41) and not w23054;
w23056 <= a(41) and not w23055;
w23057 <= not w23054 and not w23055;
w23058 <= not w23056 and not w23057;
w23059 <= w23047 and w23058;
w23060 <= not w23047 and not w23058;
w23061 <= not w23059 and not w23060;
w23062 <= not w22904 and w23061;
w23063 <= w22904 and not w23061;
w23064 <= not w23062 and not w23063;
w23065 <= not w22903 and w23064;
w23066 <= w23064 and not w23065;
w23067 <= not w22903 and not w23065;
w23068 <= not w23066 and not w23067;
w23069 <= not w22853 and not w22856;
w23070 <= w23068 and w23069;
w23071 <= not w23068 and not w23069;
w23072 <= not w23070 and not w23071;
w23073 <= b(60) and w4030;
w23074 <= b(58) and w4275;
w23075 <= b(59) and w4025;
w23076 <= not w23074 and not w23075;
w23077 <= not w23073 and w23076;
w23078 <= w4033 and w11954;
w23079 <= w23077 and not w23078;
w23080 <= a(35) and not w23079;
w23081 <= a(35) and not w23080;
w23082 <= not w23079 and not w23080;
w23083 <= not w23081 and not w23082;
w23084 <= w23072 and not w23083;
w23085 <= w23072 and not w23084;
w23086 <= not w23083 and not w23084;
w23087 <= not w23085 and not w23086;
w23088 <= not w22859 and not w22873;
w23089 <= w23087 and w23088;
w23090 <= not w23087 and not w23088;
w23091 <= not w23089 and not w23090;
w23092 <= not w22683 and not w22878;
w23093 <= b(63) and w3381;
w23094 <= b(61) and w3586;
w23095 <= b(62) and w3376;
w23096 <= not w23094 and not w23095;
w23097 <= not w23093 and w23096;
w23098 <= w3384 and w13514;
w23099 <= w23097 and not w23098;
w23100 <= a(32) and not w23099;
w23101 <= a(32) and not w23100;
w23102 <= not w23099 and not w23100;
w23103 <= not w23101 and not w23102;
w23104 <= not w23092 and not w23103;
w23105 <= not w23092 and not w23104;
w23106 <= not w23103 and not w23104;
w23107 <= not w23105 and not w23106;
w23108 <= not w23091 and w23107;
w23109 <= w23091 and not w23107;
w23110 <= not w23108 and not w23109;
w23111 <= not w22892 and w23110;
w23112 <= w22892 and not w23110;
w23113 <= not w23111 and not w23112;
w23114 <= not w22891 and w23113;
w23115 <= w22891 and not w23113;
w23116 <= not w23114 and not w23115;
w23117 <= not w23084 and not w23090;
w23118 <= b(62) and w3586;
w23119 <= b(63) and w3376;
w23120 <= not w23118 and not w23119;
w23121 <= not w3384 and w23120;
w23122 <= w13543 and w23120;
w23123 <= not w23121 and not w23122;
w23124 <= a(32) and not w23123;
w23125 <= not a(32) and w23123;
w23126 <= not w23124 and not w23125;
w23127 <= not w23117 and not w23126;
w23128 <= w23117 and w23126;
w23129 <= not w23127 and not w23128;
w23130 <= b(58) and w4778;
w23131 <= b(56) and w5020;
w23132 <= b(57) and w4773;
w23133 <= not w23131 and not w23132;
w23134 <= not w23130 and w23133;
w23135 <= w4781 and w11179;
w23136 <= w23134 and not w23135;
w23137 <= a(38) and not w23136;
w23138 <= a(38) and not w23137;
w23139 <= not w23136 and not w23137;
w23140 <= not w23138 and not w23139;
w23141 <= not w23060 and not w23062;
w23142 <= b(43) and w9082;
w23143 <= b(41) and w9475;
w23144 <= b(42) and w9077;
w23145 <= not w23143 and not w23144;
w23146 <= not w23142 and w23145;
w23147 <= w6258 and w9085;
w23148 <= w23146 and not w23147;
w23149 <= a(53) and not w23148;
w23150 <= a(53) and not w23149;
w23151 <= not w23148 and not w23149;
w23152 <= not w23150 and not w23151;
w23153 <= not w22967 and not w22973;
w23154 <= b(40) and w10169;
w23155 <= b(38) and w10539;
w23156 <= b(39) and w10164;
w23157 <= not w23155 and not w23156;
w23158 <= not w23154 and w23157;
w23159 <= w5698 and w10172;
w23160 <= w23158 and not w23159;
w23161 <= a(56) and not w23160;
w23162 <= a(56) and not w23161;
w23163 <= not w23160 and not w23161;
w23164 <= not w23162 and not w23163;
w23165 <= not w22961 and not w22964;
w23166 <= b(37) and w11274;
w23167 <= b(35) and w11639;
w23168 <= b(36) and w11269;
w23169 <= not w23167 and not w23168;
w23170 <= not w23166 and w23169;
w23171 <= w4924 and w11277;
w23172 <= w23170 and not w23171;
w23173 <= a(59) and not w23172;
w23174 <= a(59) and not w23173;
w23175 <= not w23172 and not w23173;
w23176 <= not w23174 and not w23175;
w23177 <= not w22935 and not w22946;
w23178 <= not w22932 and not w23177;
w23179 <= b(30) and w13646;
w23180 <= b(31) and not w13231;
w23181 <= not w23179 and not w23180;
w23182 <= not w22925 and not w22928;
w23183 <= not w23181 and w23182;
w23184 <= w23181 and not w23182;
w23185 <= not w23183 and not w23184;
w23186 <= b(34) and w12411;
w23187 <= b(32) and w12790;
w23188 <= b(33) and w12406;
w23189 <= not w23187 and not w23188;
w23190 <= not w23186 and w23189;
w23191 <= w4209 and w12414;
w23192 <= w23190 and not w23191;
w23193 <= a(62) and not w23192;
w23194 <= a(62) and not w23193;
w23195 <= not w23192 and not w23193;
w23196 <= not w23194 and not w23195;
w23197 <= not w23185 and w23196;
w23198 <= w23185 and not w23196;
w23199 <= not w23197 and not w23198;
w23200 <= not w23178 and w23199;
w23201 <= not w23178 and not w23200;
w23202 <= w23199 and not w23200;
w23203 <= not w23201 and not w23202;
w23204 <= not w23176 and not w23203;
w23205 <= w23176 and not w23202;
w23206 <= not w23201 and w23205;
w23207 <= not w23204 and not w23206;
w23208 <= not w23165 and w23207;
w23209 <= not w23165 and not w23208;
w23210 <= w23207 and not w23208;
w23211 <= not w23209 and not w23210;
w23212 <= not w23164 and not w23211;
w23213 <= w23164 and not w23210;
w23214 <= not w23209 and w23213;
w23215 <= not w23212 and not w23214;
w23216 <= not w23153 and w23215;
w23217 <= w23153 and not w23215;
w23218 <= not w23216 and not w23217;
w23219 <= not w23152 and w23218;
w23220 <= w23218 and not w23219;
w23221 <= not w23152 and not w23219;
w23222 <= not w23220 and not w23221;
w23223 <= not w22908 and not w22989;
w23224 <= not w22986 and not w23223;
w23225 <= w23222 and w23224;
w23226 <= not w23222 and not w23224;
w23227 <= not w23225 and not w23226;
w23228 <= b(46) and w8105;
w23229 <= b(44) and w8458;
w23230 <= b(45) and w8100;
w23231 <= not w23229 and not w23230;
w23232 <= not w23228 and w23231;
w23233 <= w7420 and w8108;
w23234 <= w23232 and not w23233;
w23235 <= a(50) and not w23234;
w23236 <= a(50) and not w23235;
w23237 <= not w23234 and not w23235;
w23238 <= not w23236 and not w23237;
w23239 <= w23227 and not w23238;
w23240 <= w23227 and not w23239;
w23241 <= not w23238 and not w23239;
w23242 <= not w23240 and not w23241;
w23243 <= not w23004 and not w23008;
w23244 <= w23242 and w23243;
w23245 <= not w23242 and not w23243;
w23246 <= not w23244 and not w23245;
w23247 <= b(49) and w7189;
w23248 <= b(47) and w7530;
w23249 <= b(48) and w7184;
w23250 <= not w23248 and not w23249;
w23251 <= not w23247 and w23250;
w23252 <= w7192 and w8368;
w23253 <= w23251 and not w23252;
w23254 <= a(47) and not w23253;
w23255 <= a(47) and not w23254;
w23256 <= not w23253 and not w23254;
w23257 <= not w23255 and not w23256;
w23258 <= w23246 and not w23257;
w23259 <= w23246 and not w23258;
w23260 <= not w23257 and not w23258;
w23261 <= not w23259 and not w23260;
w23262 <= not w23021 and not w23027;
w23263 <= w23261 and w23262;
w23264 <= not w23261 and not w23262;
w23265 <= not w23263 and not w23264;
w23266 <= b(52) and w6338;
w23267 <= b(50) and w6645;
w23268 <= b(51) and w6333;
w23269 <= not w23267 and not w23268;
w23270 <= not w23266 and w23269;
w23271 <= w6341 and w9371;
w23272 <= w23270 and not w23271;
w23273 <= a(44) and not w23272;
w23274 <= a(44) and not w23273;
w23275 <= not w23272 and not w23273;
w23276 <= not w23274 and not w23275;
w23277 <= w23265 and not w23276;
w23278 <= w23265 and not w23277;
w23279 <= not w23276 and not w23277;
w23280 <= not w23278 and not w23279;
w23281 <= not w23045 and w23280;
w23282 <= w23045 and not w23280;
w23283 <= not w23281 and not w23282;
w23284 <= b(55) and w5520;
w23285 <= b(53) and w5802;
w23286 <= b(54) and w5515;
w23287 <= not w23285 and not w23286;
w23288 <= not w23284 and w23287;
w23289 <= w5523 and w10427;
w23290 <= w23288 and not w23289;
w23291 <= a(41) and not w23290;
w23292 <= a(41) and not w23291;
w23293 <= not w23290 and not w23291;
w23294 <= not w23292 and not w23293;
w23295 <= not w23283 and not w23294;
w23296 <= w23283 and w23294;
w23297 <= not w23295 and not w23296;
w23298 <= not w23141 and w23297;
w23299 <= w23141 and not w23297;
w23300 <= not w23298 and not w23299;
w23301 <= not w23140 and w23300;
w23302 <= w23300 and not w23301;
w23303 <= not w23140 and not w23301;
w23304 <= not w23302 and not w23303;
w23305 <= not w23065 and not w23071;
w23306 <= w23304 and w23305;
w23307 <= not w23304 and not w23305;
w23308 <= not w23306 and not w23307;
w23309 <= b(61) and w4030;
w23310 <= b(59) and w4275;
w23311 <= b(60) and w4025;
w23312 <= not w23310 and not w23311;
w23313 <= not w23309 and w23312;
w23314 <= w4033 and w12712;
w23315 <= w23313 and not w23314;
w23316 <= a(35) and not w23315;
w23317 <= a(35) and not w23316;
w23318 <= not w23315 and not w23316;
w23319 <= not w23317 and not w23318;
w23320 <= w23308 and not w23319;
w23321 <= not w23308 and w23319;
w23322 <= w23129 and not w23321;
w23323 <= not w23320 and w23322;
w23324 <= w23129 and not w23323;
w23325 <= not w23321 and not w23323;
w23326 <= not w23320 and w23325;
w23327 <= not w23324 and not w23326;
w23328 <= not w23104 and not w23109;
w23329 <= not w23327 and not w23328;
w23330 <= not w23327 and not w23329;
w23331 <= not w23328 and not w23329;
w23332 <= not w23330 and not w23331;
w23333 <= not w23111 and not w23114;
w23334 <= not w23332 and not w23333;
w23335 <= w23332 and w23333;
w23336 <= not w23334 and not w23335;
w23337 <= not w23329 and not w23334;
w23338 <= not w23127 and not w23323;
w23339 <= not w23307 and not w23320;
w23340 <= b(63) and w3586;
w23341 <= w3384 and w13540;
w23342 <= not w23340 and not w23341;
w23343 <= a(32) and not w23342;
w23344 <= a(32) and not w23343;
w23345 <= not w23342 and not w23343;
w23346 <= not w23344 and not w23345;
w23347 <= not w23339 and not w23346;
w23348 <= not w23339 and not w23347;
w23349 <= not w23346 and not w23347;
w23350 <= not w23348 and not w23349;
w23351 <= not w23045 and not w23280;
w23352 <= not w23295 and not w23351;
w23353 <= b(56) and w5520;
w23354 <= b(54) and w5802;
w23355 <= b(55) and w5515;
w23356 <= not w23354 and not w23355;
w23357 <= not w23353 and w23356;
w23358 <= w5523 and w10451;
w23359 <= w23357 and not w23358;
w23360 <= a(41) and not w23359;
w23361 <= a(41) and not w23360;
w23362 <= not w23359 and not w23360;
w23363 <= not w23361 and not w23362;
w23364 <= not w23264 and not w23277;
w23365 <= b(53) and w6338;
w23366 <= b(51) and w6645;
w23367 <= b(52) and w6333;
w23368 <= not w23366 and not w23367;
w23369 <= not w23365 and w23368;
w23370 <= w6341 and w9715;
w23371 <= w23369 and not w23370;
w23372 <= a(44) and not w23371;
w23373 <= a(44) and not w23372;
w23374 <= not w23371 and not w23372;
w23375 <= not w23373 and not w23374;
w23376 <= not w23245 and not w23258;
w23377 <= not w23216 and not w23219;
w23378 <= b(44) and w9082;
w23379 <= b(42) and w9475;
w23380 <= b(43) and w9077;
w23381 <= not w23379 and not w23380;
w23382 <= not w23378 and w23381;
w23383 <= w6815 and w9085;
w23384 <= w23382 and not w23383;
w23385 <= a(53) and not w23384;
w23386 <= a(53) and not w23385;
w23387 <= not w23384 and not w23385;
w23388 <= not w23386 and not w23387;
w23389 <= not w23208 and not w23212;
w23390 <= b(41) and w10169;
w23391 <= b(39) and w10539;
w23392 <= b(40) and w10164;
w23393 <= not w23391 and not w23392;
w23394 <= not w23390 and w23393;
w23395 <= w5962 and w10172;
w23396 <= w23394 and not w23395;
w23397 <= a(56) and not w23396;
w23398 <= a(56) and not w23397;
w23399 <= not w23396 and not w23397;
w23400 <= not w23398 and not w23399;
w23401 <= not w23200 and not w23204;
w23402 <= not w23184 and not w23198;
w23403 <= b(31) and w13646;
w23404 <= b(32) and not w13231;
w23405 <= not w23403 and not w23404;
w23406 <= not w23181 and w23405;
w23407 <= w23181 and not w23405;
w23408 <= not w23402 and not w23407;
w23409 <= not w23406 and w23408;
w23410 <= not w23402 and not w23409;
w23411 <= not w23406 and not w23409;
w23412 <= not w23407 and w23411;
w23413 <= not w23410 and not w23412;
w23414 <= b(35) and w12411;
w23415 <= b(33) and w12790;
w23416 <= b(34) and w12406;
w23417 <= not w23415 and not w23416;
w23418 <= not w23414 and w23417;
w23419 <= w4439 and w12414;
w23420 <= w23418 and not w23419;
w23421 <= a(62) and not w23420;
w23422 <= a(62) and not w23421;
w23423 <= not w23420 and not w23421;
w23424 <= not w23422 and not w23423;
w23425 <= not w23413 and not w23424;
w23426 <= not w23413 and not w23425;
w23427 <= not w23424 and not w23425;
w23428 <= not w23426 and not w23427;
w23429 <= b(38) and w11274;
w23430 <= b(36) and w11639;
w23431 <= b(37) and w11269;
w23432 <= not w23430 and not w23431;
w23433 <= not w23429 and w23432;
w23434 <= w4948 and w11277;
w23435 <= w23433 and not w23434;
w23436 <= a(59) and not w23435;
w23437 <= a(59) and not w23436;
w23438 <= not w23435 and not w23436;
w23439 <= not w23437 and not w23438;
w23440 <= not w23428 and w23439;
w23441 <= w23428 and not w23439;
w23442 <= not w23440 and not w23441;
w23443 <= not w23401 and not w23442;
w23444 <= w23401 and w23442;
w23445 <= not w23443 and not w23444;
w23446 <= not w23400 and w23445;
w23447 <= w23400 and not w23445;
w23448 <= not w23446 and not w23447;
w23449 <= not w23389 and w23448;
w23450 <= w23389 and not w23448;
w23451 <= not w23449 and not w23450;
w23452 <= not w23388 and w23451;
w23453 <= w23388 and not w23451;
w23454 <= not w23452 and not w23453;
w23455 <= not w23377 and w23454;
w23456 <= w23377 and not w23454;
w23457 <= not w23455 and not w23456;
w23458 <= b(47) and w8105;
w23459 <= b(45) and w8458;
w23460 <= b(46) and w8100;
w23461 <= not w23459 and not w23460;
w23462 <= not w23458 and w23461;
w23463 <= w7446 and w8108;
w23464 <= w23462 and not w23463;
w23465 <= a(50) and not w23464;
w23466 <= a(50) and not w23465;
w23467 <= not w23464 and not w23465;
w23468 <= not w23466 and not w23467;
w23469 <= w23457 and not w23468;
w23470 <= w23457 and not w23469;
w23471 <= not w23468 and not w23469;
w23472 <= not w23470 and not w23471;
w23473 <= not w23226 and not w23239;
w23474 <= w23472 and w23473;
w23475 <= not w23472 and not w23473;
w23476 <= not w23474 and not w23475;
w23477 <= b(50) and w7189;
w23478 <= b(48) and w7530;
w23479 <= b(49) and w7184;
w23480 <= not w23478 and not w23479;
w23481 <= not w23477 and w23480;
w23482 <= w7192 and w8692;
w23483 <= w23481 and not w23482;
w23484 <= a(47) and not w23483;
w23485 <= a(47) and not w23484;
w23486 <= not w23483 and not w23484;
w23487 <= not w23485 and not w23486;
w23488 <= not w23476 and w23487;
w23489 <= w23476 and not w23487;
w23490 <= not w23488 and not w23489;
w23491 <= not w23376 and w23490;
w23492 <= not w23376 and not w23491;
w23493 <= w23490 and not w23491;
w23494 <= not w23492 and not w23493;
w23495 <= not w23375 and not w23494;
w23496 <= w23375 and not w23493;
w23497 <= not w23492 and w23496;
w23498 <= not w23495 and not w23497;
w23499 <= not w23364 and w23498;
w23500 <= w23364 and not w23498;
w23501 <= not w23499 and not w23500;
w23502 <= not w23363 and w23501;
w23503 <= w23363 and not w23501;
w23504 <= not w23502 and not w23503;
w23505 <= not w23352 and w23504;
w23506 <= w23352 and not w23504;
w23507 <= not w23505 and not w23506;
w23508 <= b(59) and w4778;
w23509 <= b(57) and w5020;
w23510 <= b(58) and w4773;
w23511 <= not w23509 and not w23510;
w23512 <= not w23508 and w23511;
w23513 <= w4781 and w11922;
w23514 <= w23512 and not w23513;
w23515 <= a(38) and not w23514;
w23516 <= a(38) and not w23515;
w23517 <= not w23514 and not w23515;
w23518 <= not w23516 and not w23517;
w23519 <= w23507 and not w23518;
w23520 <= w23507 and not w23519;
w23521 <= not w23518 and not w23519;
w23522 <= not w23520 and not w23521;
w23523 <= not w23298 and not w23301;
w23524 <= w23522 and w23523;
w23525 <= not w23522 and not w23523;
w23526 <= not w23524 and not w23525;
w23527 <= b(62) and w4030;
w23528 <= b(60) and w4275;
w23529 <= b(61) and w4025;
w23530 <= not w23528 and not w23529;
w23531 <= not w23527 and w23530;
w23532 <= w4033 and w13113;
w23533 <= w23531 and not w23532;
w23534 <= a(35) and not w23533;
w23535 <= a(35) and not w23534;
w23536 <= not w23533 and not w23534;
w23537 <= not w23535 and not w23536;
w23538 <= w23526 and not w23537;
w23539 <= w23526 and not w23538;
w23540 <= not w23537 and not w23538;
w23541 <= not w23539 and not w23540;
w23542 <= not w23350 and w23541;
w23543 <= w23350 and not w23541;
w23544 <= not w23542 and not w23543;
w23545 <= not w23338 and not w23544;
w23546 <= not w23338 and not w23545;
w23547 <= not w23544 and not w23545;
w23548 <= not w23546 and not w23547;
w23549 <= not w23337 and not w23548;
w23550 <= w23337 and not w23547;
w23551 <= not w23546 and w23550;
w23552 <= not w23549 and not w23551;
w23553 <= not w23545 and not w23549;
w23554 <= not w23350 and not w23541;
w23555 <= not w23347 and not w23554;
w23556 <= b(57) and w5520;
w23557 <= b(55) and w5802;
w23558 <= b(56) and w5515;
w23559 <= not w23557 and not w23558;
w23560 <= not w23556 and w23559;
w23561 <= w5523 and w11153;
w23562 <= w23560 and not w23561;
w23563 <= a(41) and not w23562;
w23564 <= a(41) and not w23563;
w23565 <= not w23562 and not w23563;
w23566 <= not w23564 and not w23565;
w23567 <= not w23491 and not w23495;
w23568 <= not w23475 and not w23489;
w23569 <= b(42) and w10169;
w23570 <= b(40) and w10539;
w23571 <= b(41) and w10164;
w23572 <= not w23570 and not w23571;
w23573 <= not w23569 and w23572;
w23574 <= w6232 and w10172;
w23575 <= w23573 and not w23574;
w23576 <= a(56) and not w23575;
w23577 <= a(56) and not w23576;
w23578 <= not w23575 and not w23576;
w23579 <= not w23577 and not w23578;
w23580 <= not w23428 and not w23439;
w23581 <= not w23425 and not w23580;
w23582 <= b(32) and w13646;
w23583 <= b(33) and not w13231;
w23584 <= not w23582 and not w23583;
w23585 <= not a(32) and not w23584;
w23586 <= a(32) and w23584;
w23587 <= not w23585 and not w23586;
w23588 <= not w23405 and w23587;
w23589 <= not w23405 and not w23588;
w23590 <= w23587 and not w23588;
w23591 <= not w23589 and not w23590;
w23592 <= not w23411 and not w23591;
w23593 <= not w23411 and not w23592;
w23594 <= not w23591 and not w23592;
w23595 <= not w23593 and not w23594;
w23596 <= b(36) and w12411;
w23597 <= b(34) and w12790;
w23598 <= b(35) and w12406;
w23599 <= not w23597 and not w23598;
w23600 <= not w23596 and w23599;
w23601 <= w4665 and w12414;
w23602 <= w23600 and not w23601;
w23603 <= a(62) and not w23602;
w23604 <= a(62) and not w23603;
w23605 <= not w23602 and not w23603;
w23606 <= not w23604 and not w23605;
w23607 <= not w23595 and w23606;
w23608 <= w23595 and not w23606;
w23609 <= not w23607 and not w23608;
w23610 <= b(39) and w11274;
w23611 <= b(37) and w11639;
w23612 <= b(38) and w11269;
w23613 <= not w23611 and not w23612;
w23614 <= not w23610 and w23613;
w23615 <= w5194 and w11277;
w23616 <= w23614 and not w23615;
w23617 <= a(59) and not w23616;
w23618 <= a(59) and not w23617;
w23619 <= not w23616 and not w23617;
w23620 <= not w23618 and not w23619;
w23621 <= not w23609 and not w23620;
w23622 <= w23609 and w23620;
w23623 <= not w23621 and not w23622;
w23624 <= not w23581 and w23623;
w23625 <= w23581 and not w23623;
w23626 <= not w23624 and not w23625;
w23627 <= not w23579 and w23626;
w23628 <= w23626 and not w23627;
w23629 <= not w23579 and not w23627;
w23630 <= not w23628 and not w23629;
w23631 <= not w23443 and not w23446;
w23632 <= w23630 and w23631;
w23633 <= not w23630 and not w23631;
w23634 <= not w23632 and not w23633;
w23635 <= b(45) and w9082;
w23636 <= b(43) and w9475;
w23637 <= b(44) and w9077;
w23638 <= not w23636 and not w23637;
w23639 <= not w23635 and w23638;
w23640 <= w7104 and w9085;
w23641 <= w23639 and not w23640;
w23642 <= a(53) and not w23641;
w23643 <= a(53) and not w23642;
w23644 <= not w23641 and not w23642;
w23645 <= not w23643 and not w23644;
w23646 <= w23634 and not w23645;
w23647 <= w23634 and not w23646;
w23648 <= not w23645 and not w23646;
w23649 <= not w23647 and not w23648;
w23650 <= not w23449 and not w23452;
w23651 <= w23649 and w23650;
w23652 <= not w23649 and not w23650;
w23653 <= not w23651 and not w23652;
w23654 <= b(48) and w8105;
w23655 <= b(46) and w8458;
w23656 <= b(47) and w8100;
w23657 <= not w23655 and not w23656;
w23658 <= not w23654 and w23657;
w23659 <= w7752 and w8108;
w23660 <= w23658 and not w23659;
w23661 <= a(50) and not w23660;
w23662 <= a(50) and not w23661;
w23663 <= not w23660 and not w23661;
w23664 <= not w23662 and not w23663;
w23665 <= w23653 and not w23664;
w23666 <= w23653 and not w23665;
w23667 <= not w23664 and not w23665;
w23668 <= not w23666 and not w23667;
w23669 <= not w23455 and not w23469;
w23670 <= w23668 and w23669;
w23671 <= not w23668 and not w23669;
w23672 <= not w23670 and not w23671;
w23673 <= b(51) and w7189;
w23674 <= b(49) and w7530;
w23675 <= b(50) and w7184;
w23676 <= not w23674 and not w23675;
w23677 <= not w23673 and w23676;
w23678 <= w7192 and w8719;
w23679 <= w23677 and not w23678;
w23680 <= a(47) and not w23679;
w23681 <= a(47) and not w23680;
w23682 <= not w23679 and not w23680;
w23683 <= not w23681 and not w23682;
w23684 <= w23672 and not w23683;
w23685 <= not w23672 and w23683;
w23686 <= not w23568 and not w23685;
w23687 <= not w23684 and w23686;
w23688 <= not w23568 and not w23687;
w23689 <= not w23684 and not w23687;
w23690 <= not w23685 and w23689;
w23691 <= not w23688 and not w23690;
w23692 <= b(54) and w6338;
w23693 <= b(52) and w6645;
w23694 <= b(53) and w6333;
w23695 <= not w23693 and not w23694;
w23696 <= not w23692 and w23695;
w23697 <= w6341 and w9741;
w23698 <= w23696 and not w23697;
w23699 <= a(44) and not w23698;
w23700 <= a(44) and not w23699;
w23701 <= not w23698 and not w23699;
w23702 <= not w23700 and not w23701;
w23703 <= w23691 and w23702;
w23704 <= not w23691 and not w23702;
w23705 <= not w23703 and not w23704;
w23706 <= not w23567 and w23705;
w23707 <= w23567 and not w23705;
w23708 <= not w23706 and not w23707;
w23709 <= not w23566 and w23708;
w23710 <= w23708 and not w23709;
w23711 <= not w23566 and not w23709;
w23712 <= not w23710 and not w23711;
w23713 <= not w23499 and not w23502;
w23714 <= w23712 and w23713;
w23715 <= not w23712 and not w23713;
w23716 <= not w23714 and not w23715;
w23717 <= b(60) and w4778;
w23718 <= b(58) and w5020;
w23719 <= b(59) and w4773;
w23720 <= not w23718 and not w23719;
w23721 <= not w23717 and w23720;
w23722 <= w4781 and w11954;
w23723 <= w23721 and not w23722;
w23724 <= a(38) and not w23723;
w23725 <= a(38) and not w23724;
w23726 <= not w23723 and not w23724;
w23727 <= not w23725 and not w23726;
w23728 <= w23716 and not w23727;
w23729 <= w23716 and not w23728;
w23730 <= not w23727 and not w23728;
w23731 <= not w23729 and not w23730;
w23732 <= not w23505 and not w23519;
w23733 <= w23731 and w23732;
w23734 <= not w23731 and not w23732;
w23735 <= not w23733 and not w23734;
w23736 <= not w23525 and not w23538;
w23737 <= b(63) and w4030;
w23738 <= b(61) and w4275;
w23739 <= b(62) and w4025;
w23740 <= not w23738 and not w23739;
w23741 <= not w23737 and w23740;
w23742 <= w4033 and w13514;
w23743 <= w23741 and not w23742;
w23744 <= a(35) and not w23743;
w23745 <= a(35) and not w23744;
w23746 <= not w23743 and not w23744;
w23747 <= not w23745 and not w23746;
w23748 <= not w23736 and not w23747;
w23749 <= not w23736 and not w23748;
w23750 <= not w23747 and not w23748;
w23751 <= not w23749 and not w23750;
w23752 <= not w23735 and w23751;
w23753 <= w23735 and not w23751;
w23754 <= not w23752 and not w23753;
w23755 <= not w23555 and w23754;
w23756 <= w23555 and not w23754;
w23757 <= not w23755 and not w23756;
w23758 <= not w23553 and w23757;
w23759 <= w23553 and not w23757;
w23760 <= not w23758 and not w23759;
w23761 <= not w23728 and not w23734;
w23762 <= b(62) and w4275;
w23763 <= b(63) and w4025;
w23764 <= not w23762 and not w23763;
w23765 <= not w4033 and w23764;
w23766 <= w13543 and w23764;
w23767 <= not w23765 and not w23766;
w23768 <= a(35) and not w23767;
w23769 <= not a(35) and w23767;
w23770 <= not w23768 and not w23769;
w23771 <= not w23761 and not w23770;
w23772 <= w23761 and w23770;
w23773 <= not w23771 and not w23772;
w23774 <= b(58) and w5520;
w23775 <= b(56) and w5802;
w23776 <= b(57) and w5515;
w23777 <= not w23775 and not w23776;
w23778 <= not w23774 and w23777;
w23779 <= w5523 and w11179;
w23780 <= w23778 and not w23779;
w23781 <= a(41) and not w23780;
w23782 <= a(41) and not w23781;
w23783 <= not w23780 and not w23781;
w23784 <= not w23782 and not w23783;
w23785 <= not w23704 and not w23706;
w23786 <= b(43) and w10169;
w23787 <= b(41) and w10539;
w23788 <= b(42) and w10164;
w23789 <= not w23787 and not w23788;
w23790 <= not w23786 and w23789;
w23791 <= w6258 and w10172;
w23792 <= w23790 and not w23791;
w23793 <= a(56) and not w23792;
w23794 <= a(56) and not w23793;
w23795 <= not w23792 and not w23793;
w23796 <= not w23794 and not w23795;
w23797 <= not w23621 and not w23624;
w23798 <= b(40) and w11274;
w23799 <= b(38) and w11639;
w23800 <= b(39) and w11269;
w23801 <= not w23799 and not w23800;
w23802 <= not w23798 and w23801;
w23803 <= w5698 and w11277;
w23804 <= w23802 and not w23803;
w23805 <= a(59) and not w23804;
w23806 <= a(59) and not w23805;
w23807 <= not w23804 and not w23805;
w23808 <= not w23806 and not w23807;
w23809 <= not w23595 and not w23606;
w23810 <= not w23592 and not w23809;
w23811 <= b(33) and w13646;
w23812 <= b(34) and not w13231;
w23813 <= not w23811 and not w23812;
w23814 <= not w23585 and not w23588;
w23815 <= not w23813 and w23814;
w23816 <= w23813 and not w23814;
w23817 <= not w23815 and not w23816;
w23818 <= b(37) and w12411;
w23819 <= b(35) and w12790;
w23820 <= b(36) and w12406;
w23821 <= not w23819 and not w23820;
w23822 <= not w23818 and w23821;
w23823 <= w4924 and w12414;
w23824 <= w23822 and not w23823;
w23825 <= a(62) and not w23824;
w23826 <= a(62) and not w23825;
w23827 <= not w23824 and not w23825;
w23828 <= not w23826 and not w23827;
w23829 <= not w23817 and w23828;
w23830 <= w23817 and not w23828;
w23831 <= not w23829 and not w23830;
w23832 <= not w23810 and w23831;
w23833 <= not w23810 and not w23832;
w23834 <= w23831 and not w23832;
w23835 <= not w23833 and not w23834;
w23836 <= not w23808 and not w23835;
w23837 <= w23808 and not w23834;
w23838 <= not w23833 and w23837;
w23839 <= not w23836 and not w23838;
w23840 <= not w23797 and w23839;
w23841 <= w23797 and not w23839;
w23842 <= not w23840 and not w23841;
w23843 <= not w23796 and w23842;
w23844 <= w23842 and not w23843;
w23845 <= not w23796 and not w23843;
w23846 <= not w23844 and not w23845;
w23847 <= not w23627 and not w23633;
w23848 <= w23846 and w23847;
w23849 <= not w23846 and not w23847;
w23850 <= not w23848 and not w23849;
w23851 <= b(46) and w9082;
w23852 <= b(44) and w9475;
w23853 <= b(45) and w9077;
w23854 <= not w23852 and not w23853;
w23855 <= not w23851 and w23854;
w23856 <= w7420 and w9085;
w23857 <= w23855 and not w23856;
w23858 <= a(53) and not w23857;
w23859 <= a(53) and not w23858;
w23860 <= not w23857 and not w23858;
w23861 <= not w23859 and not w23860;
w23862 <= w23850 and not w23861;
w23863 <= w23850 and not w23862;
w23864 <= not w23861 and not w23862;
w23865 <= not w23863 and not w23864;
w23866 <= not w23646 and not w23652;
w23867 <= w23865 and w23866;
w23868 <= not w23865 and not w23866;
w23869 <= not w23867 and not w23868;
w23870 <= b(49) and w8105;
w23871 <= b(47) and w8458;
w23872 <= b(48) and w8100;
w23873 <= not w23871 and not w23872;
w23874 <= not w23870 and w23873;
w23875 <= w8108 and w8368;
w23876 <= w23874 and not w23875;
w23877 <= a(50) and not w23876;
w23878 <= a(50) and not w23877;
w23879 <= not w23876 and not w23877;
w23880 <= not w23878 and not w23879;
w23881 <= w23869 and not w23880;
w23882 <= w23869 and not w23881;
w23883 <= not w23880 and not w23881;
w23884 <= not w23882 and not w23883;
w23885 <= not w23665 and not w23671;
w23886 <= w23884 and w23885;
w23887 <= not w23884 and not w23885;
w23888 <= not w23886 and not w23887;
w23889 <= b(52) and w7189;
w23890 <= b(50) and w7530;
w23891 <= b(51) and w7184;
w23892 <= not w23890 and not w23891;
w23893 <= not w23889 and w23892;
w23894 <= w7192 and w9371;
w23895 <= w23893 and not w23894;
w23896 <= a(47) and not w23895;
w23897 <= a(47) and not w23896;
w23898 <= not w23895 and not w23896;
w23899 <= not w23897 and not w23898;
w23900 <= w23888 and not w23899;
w23901 <= w23888 and not w23900;
w23902 <= not w23899 and not w23900;
w23903 <= not w23901 and not w23902;
w23904 <= not w23689 and w23903;
w23905 <= w23689 and not w23903;
w23906 <= not w23904 and not w23905;
w23907 <= b(55) and w6338;
w23908 <= b(53) and w6645;
w23909 <= b(54) and w6333;
w23910 <= not w23908 and not w23909;
w23911 <= not w23907 and w23910;
w23912 <= w6341 and w10427;
w23913 <= w23911 and not w23912;
w23914 <= a(44) and not w23913;
w23915 <= a(44) and not w23914;
w23916 <= not w23913 and not w23914;
w23917 <= not w23915 and not w23916;
w23918 <= not w23906 and not w23917;
w23919 <= w23906 and w23917;
w23920 <= not w23918 and not w23919;
w23921 <= not w23785 and w23920;
w23922 <= w23785 and not w23920;
w23923 <= not w23921 and not w23922;
w23924 <= not w23784 and w23923;
w23925 <= w23923 and not w23924;
w23926 <= not w23784 and not w23924;
w23927 <= not w23925 and not w23926;
w23928 <= not w23709 and not w23715;
w23929 <= w23927 and w23928;
w23930 <= not w23927 and not w23928;
w23931 <= not w23929 and not w23930;
w23932 <= b(61) and w4778;
w23933 <= b(59) and w5020;
w23934 <= b(60) and w4773;
w23935 <= not w23933 and not w23934;
w23936 <= not w23932 and w23935;
w23937 <= w4781 and w12712;
w23938 <= w23936 and not w23937;
w23939 <= a(38) and not w23938;
w23940 <= a(38) and not w23939;
w23941 <= not w23938 and not w23939;
w23942 <= not w23940 and not w23941;
w23943 <= w23931 and not w23942;
w23944 <= not w23931 and w23942;
w23945 <= w23773 and not w23944;
w23946 <= not w23943 and w23945;
w23947 <= w23773 and not w23946;
w23948 <= not w23944 and not w23946;
w23949 <= not w23943 and w23948;
w23950 <= not w23947 and not w23949;
w23951 <= not w23748 and not w23753;
w23952 <= not w23950 and not w23951;
w23953 <= not w23950 and not w23952;
w23954 <= not w23951 and not w23952;
w23955 <= not w23953 and not w23954;
w23956 <= not w23755 and not w23758;
w23957 <= not w23955 and not w23956;
w23958 <= w23955 and w23956;
w23959 <= not w23957 and not w23958;
w23960 <= not w23952 and not w23957;
w23961 <= not w23771 and not w23946;
w23962 <= not w23930 and not w23943;
w23963 <= b(63) and w4275;
w23964 <= w4033 and w13540;
w23965 <= not w23963 and not w23964;
w23966 <= a(35) and not w23965;
w23967 <= a(35) and not w23966;
w23968 <= not w23965 and not w23966;
w23969 <= not w23967 and not w23968;
w23970 <= not w23962 and not w23969;
w23971 <= not w23962 and not w23970;
w23972 <= not w23969 and not w23970;
w23973 <= not w23971 and not w23972;
w23974 <= not w23689 and not w23903;
w23975 <= not w23918 and not w23974;
w23976 <= b(56) and w6338;
w23977 <= b(54) and w6645;
w23978 <= b(55) and w6333;
w23979 <= not w23977 and not w23978;
w23980 <= not w23976 and w23979;
w23981 <= w6341 and w10451;
w23982 <= w23980 and not w23981;
w23983 <= a(44) and not w23982;
w23984 <= a(44) and not w23983;
w23985 <= not w23982 and not w23983;
w23986 <= not w23984 and not w23985;
w23987 <= not w23887 and not w23900;
w23988 <= b(53) and w7189;
w23989 <= b(51) and w7530;
w23990 <= b(52) and w7184;
w23991 <= not w23989 and not w23990;
w23992 <= not w23988 and w23991;
w23993 <= w7192 and w9715;
w23994 <= w23992 and not w23993;
w23995 <= a(47) and not w23994;
w23996 <= a(47) and not w23995;
w23997 <= not w23994 and not w23995;
w23998 <= not w23996 and not w23997;
w23999 <= not w23868 and not w23881;
w24000 <= not w23840 and not w23843;
w24001 <= b(44) and w10169;
w24002 <= b(42) and w10539;
w24003 <= b(43) and w10164;
w24004 <= not w24002 and not w24003;
w24005 <= not w24001 and w24004;
w24006 <= w6815 and w10172;
w24007 <= w24005 and not w24006;
w24008 <= a(56) and not w24007;
w24009 <= a(56) and not w24008;
w24010 <= not w24007 and not w24008;
w24011 <= not w24009 and not w24010;
w24012 <= not w23832 and not w23836;
w24013 <= not w23816 and not w23830;
w24014 <= b(34) and w13646;
w24015 <= b(35) and not w13231;
w24016 <= not w24014 and not w24015;
w24017 <= not w23813 and w24016;
w24018 <= w23813 and not w24016;
w24019 <= not w24013 and not w24018;
w24020 <= not w24017 and w24019;
w24021 <= not w24013 and not w24020;
w24022 <= not w24017 and not w24020;
w24023 <= not w24018 and w24022;
w24024 <= not w24021 and not w24023;
w24025 <= b(38) and w12411;
w24026 <= b(36) and w12790;
w24027 <= b(37) and w12406;
w24028 <= not w24026 and not w24027;
w24029 <= not w24025 and w24028;
w24030 <= w4948 and w12414;
w24031 <= w24029 and not w24030;
w24032 <= a(62) and not w24031;
w24033 <= a(62) and not w24032;
w24034 <= not w24031 and not w24032;
w24035 <= not w24033 and not w24034;
w24036 <= not w24024 and not w24035;
w24037 <= not w24024 and not w24036;
w24038 <= not w24035 and not w24036;
w24039 <= not w24037 and not w24038;
w24040 <= b(41) and w11274;
w24041 <= b(39) and w11639;
w24042 <= b(40) and w11269;
w24043 <= not w24041 and not w24042;
w24044 <= not w24040 and w24043;
w24045 <= w5962 and w11277;
w24046 <= w24044 and not w24045;
w24047 <= a(59) and not w24046;
w24048 <= a(59) and not w24047;
w24049 <= not w24046 and not w24047;
w24050 <= not w24048 and not w24049;
w24051 <= not w24039 and w24050;
w24052 <= w24039 and not w24050;
w24053 <= not w24051 and not w24052;
w24054 <= not w24012 and not w24053;
w24055 <= w24012 and w24053;
w24056 <= not w24054 and not w24055;
w24057 <= not w24011 and w24056;
w24058 <= w24011 and not w24056;
w24059 <= not w24057 and not w24058;
w24060 <= not w24000 and w24059;
w24061 <= w24000 and not w24059;
w24062 <= not w24060 and not w24061;
w24063 <= b(47) and w9082;
w24064 <= b(45) and w9475;
w24065 <= b(46) and w9077;
w24066 <= not w24064 and not w24065;
w24067 <= not w24063 and w24066;
w24068 <= w7446 and w9085;
w24069 <= w24067 and not w24068;
w24070 <= a(53) and not w24069;
w24071 <= a(53) and not w24070;
w24072 <= not w24069 and not w24070;
w24073 <= not w24071 and not w24072;
w24074 <= w24062 and not w24073;
w24075 <= w24062 and not w24074;
w24076 <= not w24073 and not w24074;
w24077 <= not w24075 and not w24076;
w24078 <= not w23849 and not w23862;
w24079 <= w24077 and w24078;
w24080 <= not w24077 and not w24078;
w24081 <= not w24079 and not w24080;
w24082 <= b(50) and w8105;
w24083 <= b(48) and w8458;
w24084 <= b(49) and w8100;
w24085 <= not w24083 and not w24084;
w24086 <= not w24082 and w24085;
w24087 <= w8108 and w8692;
w24088 <= w24086 and not w24087;
w24089 <= a(50) and not w24088;
w24090 <= a(50) and not w24089;
w24091 <= not w24088 and not w24089;
w24092 <= not w24090 and not w24091;
w24093 <= not w24081 and w24092;
w24094 <= w24081 and not w24092;
w24095 <= not w24093 and not w24094;
w24096 <= not w23999 and w24095;
w24097 <= not w23999 and not w24096;
w24098 <= w24095 and not w24096;
w24099 <= not w24097 and not w24098;
w24100 <= not w23998 and not w24099;
w24101 <= w23998 and not w24098;
w24102 <= not w24097 and w24101;
w24103 <= not w24100 and not w24102;
w24104 <= not w23987 and w24103;
w24105 <= w23987 and not w24103;
w24106 <= not w24104 and not w24105;
w24107 <= not w23986 and w24106;
w24108 <= w23986 and not w24106;
w24109 <= not w24107 and not w24108;
w24110 <= not w23975 and w24109;
w24111 <= w23975 and not w24109;
w24112 <= not w24110 and not w24111;
w24113 <= b(59) and w5520;
w24114 <= b(57) and w5802;
w24115 <= b(58) and w5515;
w24116 <= not w24114 and not w24115;
w24117 <= not w24113 and w24116;
w24118 <= w5523 and w11922;
w24119 <= w24117 and not w24118;
w24120 <= a(41) and not w24119;
w24121 <= a(41) and not w24120;
w24122 <= not w24119 and not w24120;
w24123 <= not w24121 and not w24122;
w24124 <= w24112 and not w24123;
w24125 <= w24112 and not w24124;
w24126 <= not w24123 and not w24124;
w24127 <= not w24125 and not w24126;
w24128 <= not w23921 and not w23924;
w24129 <= w24127 and w24128;
w24130 <= not w24127 and not w24128;
w24131 <= not w24129 and not w24130;
w24132 <= b(62) and w4778;
w24133 <= b(60) and w5020;
w24134 <= b(61) and w4773;
w24135 <= not w24133 and not w24134;
w24136 <= not w24132 and w24135;
w24137 <= w4781 and w13113;
w24138 <= w24136 and not w24137;
w24139 <= a(38) and not w24138;
w24140 <= a(38) and not w24139;
w24141 <= not w24138 and not w24139;
w24142 <= not w24140 and not w24141;
w24143 <= w24131 and not w24142;
w24144 <= w24131 and not w24143;
w24145 <= not w24142 and not w24143;
w24146 <= not w24144 and not w24145;
w24147 <= not w23973 and w24146;
w24148 <= w23973 and not w24146;
w24149 <= not w24147 and not w24148;
w24150 <= not w23961 and not w24149;
w24151 <= w23961 and w24149;
w24152 <= not w24150 and not w24151;
w24153 <= not w23960 and w24152;
w24154 <= w23960 and not w24152;
w24155 <= not w24153 and not w24154;
w24156 <= not w24150 and not w24153;
w24157 <= not w24096 and not w24100;
w24158 <= b(54) and w7189;
w24159 <= b(52) and w7530;
w24160 <= b(53) and w7184;
w24161 <= not w24159 and not w24160;
w24162 <= not w24158 and w24161;
w24163 <= w7192 and w9741;
w24164 <= w24162 and not w24163;
w24165 <= a(47) and not w24164;
w24166 <= a(47) and not w24165;
w24167 <= not w24164 and not w24165;
w24168 <= not w24166 and not w24167;
w24169 <= not w24080 and not w24094;
w24170 <= b(35) and w13646;
w24171 <= b(36) and not w13231;
w24172 <= not w24170 and not w24171;
w24173 <= a(35) and not w24016;
w24174 <= not a(35) and w24016;
w24175 <= not w24173 and not w24174;
w24176 <= not w24172 and not w24175;
w24177 <= w24172 and w24175;
w24178 <= not w24176 and not w24177;
w24179 <= not w24022 and w24178;
w24180 <= w24022 and not w24178;
w24181 <= not w24179 and not w24180;
w24182 <= b(39) and w12411;
w24183 <= b(37) and w12790;
w24184 <= b(38) and w12406;
w24185 <= not w24183 and not w24184;
w24186 <= not w24182 and w24185;
w24187 <= w5194 and w12414;
w24188 <= w24186 and not w24187;
w24189 <= a(62) and not w24188;
w24190 <= a(62) and not w24189;
w24191 <= not w24188 and not w24189;
w24192 <= not w24190 and not w24191;
w24193 <= not w24181 and w24192;
w24194 <= w24181 and not w24192;
w24195 <= not w24193 and not w24194;
w24196 <= b(42) and w11274;
w24197 <= b(40) and w11639;
w24198 <= b(41) and w11269;
w24199 <= not w24197 and not w24198;
w24200 <= not w24196 and w24199;
w24201 <= w6232 and w11277;
w24202 <= w24200 and not w24201;
w24203 <= a(59) and not w24202;
w24204 <= a(59) and not w24203;
w24205 <= not w24202 and not w24203;
w24206 <= not w24204 and not w24205;
w24207 <= w24195 and not w24206;
w24208 <= w24195 and not w24207;
w24209 <= not w24206 and not w24207;
w24210 <= not w24208 and not w24209;
w24211 <= not w24039 and not w24050;
w24212 <= not w24036 and not w24211;
w24213 <= not w24210 and not w24212;
w24214 <= not w24210 and not w24213;
w24215 <= not w24212 and not w24213;
w24216 <= not w24214 and not w24215;
w24217 <= b(45) and w10169;
w24218 <= b(43) and w10539;
w24219 <= b(44) and w10164;
w24220 <= not w24218 and not w24219;
w24221 <= not w24217 and w24220;
w24222 <= w7104 and w10172;
w24223 <= w24221 and not w24222;
w24224 <= a(56) and not w24223;
w24225 <= a(56) and not w24224;
w24226 <= not w24223 and not w24224;
w24227 <= not w24225 and not w24226;
w24228 <= not w24216 and not w24227;
w24229 <= not w24216 and not w24228;
w24230 <= not w24227 and not w24228;
w24231 <= not w24229 and not w24230;
w24232 <= not w24054 and not w24057;
w24233 <= w24231 and w24232;
w24234 <= not w24231 and not w24232;
w24235 <= not w24233 and not w24234;
w24236 <= b(48) and w9082;
w24237 <= b(46) and w9475;
w24238 <= b(47) and w9077;
w24239 <= not w24237 and not w24238;
w24240 <= not w24236 and w24239;
w24241 <= w7752 and w9085;
w24242 <= w24240 and not w24241;
w24243 <= a(53) and not w24242;
w24244 <= a(53) and not w24243;
w24245 <= not w24242 and not w24243;
w24246 <= not w24244 and not w24245;
w24247 <= w24235 and not w24246;
w24248 <= w24235 and not w24247;
w24249 <= not w24246 and not w24247;
w24250 <= not w24248 and not w24249;
w24251 <= not w24060 and not w24074;
w24252 <= w24250 and w24251;
w24253 <= not w24250 and not w24251;
w24254 <= not w24252 and not w24253;
w24255 <= b(51) and w8105;
w24256 <= b(49) and w8458;
w24257 <= b(50) and w8100;
w24258 <= not w24256 and not w24257;
w24259 <= not w24255 and w24258;
w24260 <= w8108 and w8719;
w24261 <= w24259 and not w24260;
w24262 <= a(50) and not w24261;
w24263 <= a(50) and not w24262;
w24264 <= not w24261 and not w24262;
w24265 <= not w24263 and not w24264;
w24266 <= not w24254 and w24265;
w24267 <= w24254 and not w24265;
w24268 <= not w24266 and not w24267;
w24269 <= not w24169 and w24268;
w24270 <= w24169 and not w24268;
w24271 <= not w24269 and not w24270;
w24272 <= not w24168 and w24271;
w24273 <= w24168 and not w24271;
w24274 <= not w24272 and not w24273;
w24275 <= not w24157 and w24274;
w24276 <= w24157 and not w24274;
w24277 <= not w24275 and not w24276;
w24278 <= b(57) and w6338;
w24279 <= b(55) and w6645;
w24280 <= b(56) and w6333;
w24281 <= not w24279 and not w24280;
w24282 <= not w24278 and w24281;
w24283 <= w6341 and w11153;
w24284 <= w24282 and not w24283;
w24285 <= a(44) and not w24284;
w24286 <= a(44) and not w24285;
w24287 <= not w24284 and not w24285;
w24288 <= not w24286 and not w24287;
w24289 <= w24277 and not w24288;
w24290 <= w24277 and not w24289;
w24291 <= not w24288 and not w24289;
w24292 <= not w24290 and not w24291;
w24293 <= not w24104 and not w24107;
w24294 <= w24292 and w24293;
w24295 <= not w24292 and not w24293;
w24296 <= not w24294 and not w24295;
w24297 <= b(60) and w5520;
w24298 <= b(58) and w5802;
w24299 <= b(59) and w5515;
w24300 <= not w24298 and not w24299;
w24301 <= not w24297 and w24300;
w24302 <= w5523 and w11954;
w24303 <= w24301 and not w24302;
w24304 <= a(41) and not w24303;
w24305 <= a(41) and not w24304;
w24306 <= not w24303 and not w24304;
w24307 <= not w24305 and not w24306;
w24308 <= w24296 and not w24307;
w24309 <= w24296 and not w24308;
w24310 <= not w24307 and not w24308;
w24311 <= not w24309 and not w24310;
w24312 <= not w24110 and not w24124;
w24313 <= w24311 and w24312;
w24314 <= not w24311 and not w24312;
w24315 <= not w24313 and not w24314;
w24316 <= b(63) and w4778;
w24317 <= b(61) and w5020;
w24318 <= b(62) and w4773;
w24319 <= not w24317 and not w24318;
w24320 <= not w24316 and w24319;
w24321 <= w4781 and w13514;
w24322 <= w24320 and not w24321;
w24323 <= a(38) and not w24322;
w24324 <= a(38) and not w24323;
w24325 <= not w24322 and not w24323;
w24326 <= not w24324 and not w24325;
w24327 <= w24315 and not w24326;
w24328 <= w24315 and not w24327;
w24329 <= not w24326 and not w24327;
w24330 <= not w24328 and not w24329;
w24331 <= not w24130 and not w24143;
w24332 <= w24330 and w24331;
w24333 <= not w24330 and not w24331;
w24334 <= not w24332 and not w24333;
w24335 <= not w23973 and not w24146;
w24336 <= not w23970 and not w24335;
w24337 <= w24334 and not w24336;
w24338 <= not w24334 and w24336;
w24339 <= not w24337 and not w24338;
w24340 <= not w24156 and w24339;
w24341 <= w24156 and not w24339;
w24342 <= not w24340 and not w24341;
w24343 <= not w24308 and not w24314;
w24344 <= b(62) and w5020;
w24345 <= b(63) and w4773;
w24346 <= not w24344 and not w24345;
w24347 <= not w4781 and w24346;
w24348 <= w13543 and w24346;
w24349 <= not w24347 and not w24348;
w24350 <= a(38) and not w24349;
w24351 <= not a(38) and w24349;
w24352 <= not w24350 and not w24351;
w24353 <= not w24343 and not w24352;
w24354 <= w24343 and w24352;
w24355 <= not w24353 and not w24354;
w24356 <= b(40) and w12411;
w24357 <= b(38) and w12790;
w24358 <= b(39) and w12406;
w24359 <= not w24357 and not w24358;
w24360 <= not w24356 and w24359;
w24361 <= w5698 and w12414;
w24362 <= w24360 and not w24361;
w24363 <= a(62) and not w24362;
w24364 <= a(62) and not w24363;
w24365 <= not w24362 and not w24363;
w24366 <= not w24364 and not w24365;
w24367 <= b(36) and w13646;
w24368 <= b(37) and not w13231;
w24369 <= not w24367 and not w24368;
w24370 <= not a(35) and not w24016;
w24371 <= not w24176 and not w24370;
w24372 <= w24369 and not w24371;
w24373 <= w24369 and not w24372;
w24374 <= not w24371 and not w24372;
w24375 <= not w24373 and not w24374;
w24376 <= not w24366 and not w24375;
w24377 <= not w24366 and not w24376;
w24378 <= not w24375 and not w24376;
w24379 <= not w24377 and not w24378;
w24380 <= not w24179 and not w24194;
w24381 <= w24379 and w24380;
w24382 <= not w24379 and not w24380;
w24383 <= not w24381 and not w24382;
w24384 <= b(43) and w11274;
w24385 <= b(41) and w11639;
w24386 <= b(42) and w11269;
w24387 <= not w24385 and not w24386;
w24388 <= not w24384 and w24387;
w24389 <= w6258 and w11277;
w24390 <= w24388 and not w24389;
w24391 <= a(59) and not w24390;
w24392 <= a(59) and not w24391;
w24393 <= not w24390 and not w24391;
w24394 <= not w24392 and not w24393;
w24395 <= w24383 and not w24394;
w24396 <= w24383 and not w24395;
w24397 <= not w24394 and not w24395;
w24398 <= not w24396 and not w24397;
w24399 <= not w24207 and not w24213;
w24400 <= w24398 and w24399;
w24401 <= not w24398 and not w24399;
w24402 <= not w24400 and not w24401;
w24403 <= b(46) and w10169;
w24404 <= b(44) and w10539;
w24405 <= b(45) and w10164;
w24406 <= not w24404 and not w24405;
w24407 <= not w24403 and w24406;
w24408 <= w7420 and w10172;
w24409 <= w24407 and not w24408;
w24410 <= a(56) and not w24409;
w24411 <= a(56) and not w24410;
w24412 <= not w24409 and not w24410;
w24413 <= not w24411 and not w24412;
w24414 <= w24402 and not w24413;
w24415 <= w24402 and not w24414;
w24416 <= not w24413 and not w24414;
w24417 <= not w24415 and not w24416;
w24418 <= not w24228 and not w24234;
w24419 <= w24417 and w24418;
w24420 <= not w24417 and not w24418;
w24421 <= not w24419 and not w24420;
w24422 <= b(49) and w9082;
w24423 <= b(47) and w9475;
w24424 <= b(48) and w9077;
w24425 <= not w24423 and not w24424;
w24426 <= not w24422 and w24425;
w24427 <= w8368 and w9085;
w24428 <= w24426 and not w24427;
w24429 <= a(53) and not w24428;
w24430 <= a(53) and not w24429;
w24431 <= not w24428 and not w24429;
w24432 <= not w24430 and not w24431;
w24433 <= w24421 and not w24432;
w24434 <= w24421 and not w24433;
w24435 <= not w24432 and not w24433;
w24436 <= not w24434 and not w24435;
w24437 <= not w24247 and not w24253;
w24438 <= w24436 and w24437;
w24439 <= not w24436 and not w24437;
w24440 <= not w24438 and not w24439;
w24441 <= b(52) and w8105;
w24442 <= b(50) and w8458;
w24443 <= b(51) and w8100;
w24444 <= not w24442 and not w24443;
w24445 <= not w24441 and w24444;
w24446 <= w8108 and w9371;
w24447 <= w24445 and not w24446;
w24448 <= a(50) and not w24447;
w24449 <= a(50) and not w24448;
w24450 <= not w24447 and not w24448;
w24451 <= not w24449 and not w24450;
w24452 <= w24440 and not w24451;
w24453 <= w24440 and not w24452;
w24454 <= not w24451 and not w24452;
w24455 <= not w24453 and not w24454;
w24456 <= not w24267 and not w24269;
w24457 <= not w24455 and not w24456;
w24458 <= not w24455 and not w24457;
w24459 <= not w24456 and not w24457;
w24460 <= not w24458 and not w24459;
w24461 <= b(55) and w7189;
w24462 <= b(53) and w7530;
w24463 <= b(54) and w7184;
w24464 <= not w24462 and not w24463;
w24465 <= not w24461 and w24464;
w24466 <= w7192 and w10427;
w24467 <= w24465 and not w24466;
w24468 <= a(47) and not w24467;
w24469 <= a(47) and not w24468;
w24470 <= not w24467 and not w24468;
w24471 <= not w24469 and not w24470;
w24472 <= not w24460 and not w24471;
w24473 <= not w24460 and not w24472;
w24474 <= not w24471 and not w24472;
w24475 <= not w24473 and not w24474;
w24476 <= not w24272 and not w24275;
w24477 <= w24475 and w24476;
w24478 <= not w24475 and not w24476;
w24479 <= not w24477 and not w24478;
w24480 <= b(58) and w6338;
w24481 <= b(56) and w6645;
w24482 <= b(57) and w6333;
w24483 <= not w24481 and not w24482;
w24484 <= not w24480 and w24483;
w24485 <= w6341 and w11179;
w24486 <= w24484 and not w24485;
w24487 <= a(44) and not w24486;
w24488 <= a(44) and not w24487;
w24489 <= not w24486 and not w24487;
w24490 <= not w24488 and not w24489;
w24491 <= w24479 and not w24490;
w24492 <= w24479 and not w24491;
w24493 <= not w24490 and not w24491;
w24494 <= not w24492 and not w24493;
w24495 <= not w24289 and not w24295;
w24496 <= w24494 and w24495;
w24497 <= not w24494 and not w24495;
w24498 <= not w24496 and not w24497;
w24499 <= b(61) and w5520;
w24500 <= b(59) and w5802;
w24501 <= b(60) and w5515;
w24502 <= not w24500 and not w24501;
w24503 <= not w24499 and w24502;
w24504 <= w5523 and w12712;
w24505 <= w24503 and not w24504;
w24506 <= a(41) and not w24505;
w24507 <= a(41) and not w24506;
w24508 <= not w24505 and not w24506;
w24509 <= not w24507 and not w24508;
w24510 <= w24498 and not w24509;
w24511 <= not w24498 and w24509;
w24512 <= w24355 and not w24511;
w24513 <= not w24510 and w24512;
w24514 <= w24355 and not w24513;
w24515 <= not w24511 and not w24513;
w24516 <= not w24510 and w24515;
w24517 <= not w24514 and not w24516;
w24518 <= not w24327 and not w24333;
w24519 <= w24517 and w24518;
w24520 <= not w24517 and not w24518;
w24521 <= not w24519 and not w24520;
w24522 <= not w24337 and not w24340;
w24523 <= w24521 and not w24522;
w24524 <= not w24521 and w24522;
w24525 <= not w24523 and not w24524;
w24526 <= not w24520 and not w24523;
w24527 <= not w24353 and not w24513;
w24528 <= not w24497 and not w24510;
w24529 <= b(63) and w5020;
w24530 <= w4781 and w13540;
w24531 <= not w24529 and not w24530;
w24532 <= a(38) and not w24531;
w24533 <= a(38) and not w24532;
w24534 <= not w24531 and not w24532;
w24535 <= not w24533 and not w24534;
w24536 <= not w24528 and not w24535;
w24537 <= not w24528 and not w24536;
w24538 <= not w24535 and not w24536;
w24539 <= not w24537 and not w24538;
w24540 <= not w24457 and not w24472;
w24541 <= b(56) and w7189;
w24542 <= b(54) and w7530;
w24543 <= b(55) and w7184;
w24544 <= not w24542 and not w24543;
w24545 <= not w24541 and w24544;
w24546 <= w7192 and w10451;
w24547 <= w24545 and not w24546;
w24548 <= a(47) and not w24547;
w24549 <= a(47) and not w24548;
w24550 <= not w24547 and not w24548;
w24551 <= not w24549 and not w24550;
w24552 <= not w24439 and not w24452;
w24553 <= b(53) and w8105;
w24554 <= b(51) and w8458;
w24555 <= b(52) and w8100;
w24556 <= not w24554 and not w24555;
w24557 <= not w24553 and w24556;
w24558 <= w8108 and w9715;
w24559 <= w24557 and not w24558;
w24560 <= a(50) and not w24559;
w24561 <= a(50) and not w24560;
w24562 <= not w24559 and not w24560;
w24563 <= not w24561 and not w24562;
w24564 <= not w24420 and not w24433;
w24565 <= not w24372 and not w24376;
w24566 <= b(37) and w13646;
w24567 <= b(38) and not w13231;
w24568 <= not w24566 and not w24567;
w24569 <= w24369 and not w24568;
w24570 <= w24369 and not w24569;
w24571 <= not w24568 and not w24569;
w24572 <= not w24570 and not w24571;
w24573 <= not w24565 and not w24572;
w24574 <= not w24565 and not w24573;
w24575 <= not w24572 and not w24573;
w24576 <= not w24574 and not w24575;
w24577 <= b(41) and w12411;
w24578 <= b(39) and w12790;
w24579 <= b(40) and w12406;
w24580 <= not w24578 and not w24579;
w24581 <= not w24577 and w24580;
w24582 <= w5962 and w12414;
w24583 <= w24581 and not w24582;
w24584 <= a(62) and not w24583;
w24585 <= a(62) and not w24584;
w24586 <= not w24583 and not w24584;
w24587 <= not w24585 and not w24586;
w24588 <= not w24576 and not w24587;
w24589 <= not w24576 and not w24588;
w24590 <= not w24587 and not w24588;
w24591 <= not w24589 and not w24590;
w24592 <= b(44) and w11274;
w24593 <= b(42) and w11639;
w24594 <= b(43) and w11269;
w24595 <= not w24593 and not w24594;
w24596 <= not w24592 and w24595;
w24597 <= w6815 and w11277;
w24598 <= w24596 and not w24597;
w24599 <= a(59) and not w24598;
w24600 <= a(59) and not w24599;
w24601 <= not w24598 and not w24599;
w24602 <= not w24600 and not w24601;
w24603 <= not w24591 and w24602;
w24604 <= w24591 and not w24602;
w24605 <= not w24603 and not w24604;
w24606 <= not w24382 and not w24395;
w24607 <= w24605 and w24606;
w24608 <= not w24605 and not w24606;
w24609 <= not w24607 and not w24608;
w24610 <= b(47) and w10169;
w24611 <= b(45) and w10539;
w24612 <= b(46) and w10164;
w24613 <= not w24611 and not w24612;
w24614 <= not w24610 and w24613;
w24615 <= w7446 and w10172;
w24616 <= w24614 and not w24615;
w24617 <= a(56) and not w24616;
w24618 <= a(56) and not w24617;
w24619 <= not w24616 and not w24617;
w24620 <= not w24618 and not w24619;
w24621 <= w24609 and not w24620;
w24622 <= w24609 and not w24621;
w24623 <= not w24620 and not w24621;
w24624 <= not w24622 and not w24623;
w24625 <= not w24401 and not w24414;
w24626 <= w24624 and w24625;
w24627 <= not w24624 and not w24625;
w24628 <= not w24626 and not w24627;
w24629 <= b(50) and w9082;
w24630 <= b(48) and w9475;
w24631 <= b(49) and w9077;
w24632 <= not w24630 and not w24631;
w24633 <= not w24629 and w24632;
w24634 <= w8692 and w9085;
w24635 <= w24633 and not w24634;
w24636 <= a(53) and not w24635;
w24637 <= a(53) and not w24636;
w24638 <= not w24635 and not w24636;
w24639 <= not w24637 and not w24638;
w24640 <= not w24628 and w24639;
w24641 <= w24628 and not w24639;
w24642 <= not w24640 and not w24641;
w24643 <= not w24564 and w24642;
w24644 <= not w24564 and not w24643;
w24645 <= w24642 and not w24643;
w24646 <= not w24644 and not w24645;
w24647 <= not w24563 and not w24646;
w24648 <= w24563 and not w24645;
w24649 <= not w24644 and w24648;
w24650 <= not w24647 and not w24649;
w24651 <= not w24552 and w24650;
w24652 <= w24552 and not w24650;
w24653 <= not w24651 and not w24652;
w24654 <= not w24551 and w24653;
w24655 <= w24551 and not w24653;
w24656 <= not w24654 and not w24655;
w24657 <= not w24540 and w24656;
w24658 <= w24540 and not w24656;
w24659 <= not w24657 and not w24658;
w24660 <= b(59) and w6338;
w24661 <= b(57) and w6645;
w24662 <= b(58) and w6333;
w24663 <= not w24661 and not w24662;
w24664 <= not w24660 and w24663;
w24665 <= w6341 and w11922;
w24666 <= w24664 and not w24665;
w24667 <= a(44) and not w24666;
w24668 <= a(44) and not w24667;
w24669 <= not w24666 and not w24667;
w24670 <= not w24668 and not w24669;
w24671 <= w24659 and not w24670;
w24672 <= w24659 and not w24671;
w24673 <= not w24670 and not w24671;
w24674 <= not w24672 and not w24673;
w24675 <= not w24478 and not w24491;
w24676 <= w24674 and w24675;
w24677 <= not w24674 and not w24675;
w24678 <= not w24676 and not w24677;
w24679 <= b(62) and w5520;
w24680 <= b(60) and w5802;
w24681 <= b(61) and w5515;
w24682 <= not w24680 and not w24681;
w24683 <= not w24679 and w24682;
w24684 <= w5523 and w13113;
w24685 <= w24683 and not w24684;
w24686 <= a(41) and not w24685;
w24687 <= a(41) and not w24686;
w24688 <= not w24685 and not w24686;
w24689 <= not w24687 and not w24688;
w24690 <= w24678 and not w24689;
w24691 <= w24678 and not w24690;
w24692 <= not w24689 and not w24690;
w24693 <= not w24691 and not w24692;
w24694 <= not w24539 and w24693;
w24695 <= w24539 and not w24693;
w24696 <= not w24694 and not w24695;
w24697 <= not w24527 and not w24696;
w24698 <= w24527 and w24696;
w24699 <= not w24697 and not w24698;
w24700 <= not w24526 and w24699;
w24701 <= w24526 and not w24699;
w24702 <= not w24700 and not w24701;
w24703 <= not w24697 and not w24700;
w24704 <= not w24643 and not w24647;
w24705 <= b(54) and w8105;
w24706 <= b(52) and w8458;
w24707 <= b(53) and w8100;
w24708 <= not w24706 and not w24707;
w24709 <= not w24705 and w24708;
w24710 <= w8108 and w9741;
w24711 <= w24709 and not w24710;
w24712 <= a(50) and not w24711;
w24713 <= a(50) and not w24712;
w24714 <= not w24711 and not w24712;
w24715 <= not w24713 and not w24714;
w24716 <= not w24627 and not w24641;
w24717 <= not w24569 and not w24573;
w24718 <= b(38) and w13646;
w24719 <= b(39) and not w13231;
w24720 <= not w24718 and not w24719;
w24721 <= a(38) and not w24369;
w24722 <= not a(38) and w24369;
w24723 <= not w24721 and not w24722;
w24724 <= not w24720 and not w24723;
w24725 <= w24720 and w24723;
w24726 <= not w24724 and not w24725;
w24727 <= not w24717 and w24726;
w24728 <= w24717 and not w24726;
w24729 <= not w24727 and not w24728;
w24730 <= b(42) and w12411;
w24731 <= b(40) and w12790;
w24732 <= b(41) and w12406;
w24733 <= not w24731 and not w24732;
w24734 <= not w24730 and w24733;
w24735 <= w6232 and w12414;
w24736 <= w24734 and not w24735;
w24737 <= a(62) and not w24736;
w24738 <= a(62) and not w24737;
w24739 <= not w24736 and not w24737;
w24740 <= not w24738 and not w24739;
w24741 <= w24729 and not w24740;
w24742 <= w24729 and not w24741;
w24743 <= not w24740 and not w24741;
w24744 <= not w24742 and not w24743;
w24745 <= b(45) and w11274;
w24746 <= b(43) and w11639;
w24747 <= b(44) and w11269;
w24748 <= not w24746 and not w24747;
w24749 <= not w24745 and w24748;
w24750 <= w7104 and w11277;
w24751 <= w24749 and not w24750;
w24752 <= a(59) and not w24751;
w24753 <= a(59) and not w24752;
w24754 <= not w24751 and not w24752;
w24755 <= not w24753 and not w24754;
w24756 <= not w24744 and not w24755;
w24757 <= not w24744 and not w24756;
w24758 <= not w24755 and not w24756;
w24759 <= not w24757 and not w24758;
w24760 <= not w24591 and not w24602;
w24761 <= not w24588 and not w24760;
w24762 <= not w24759 and not w24761;
w24763 <= not w24759 and not w24762;
w24764 <= not w24761 and not w24762;
w24765 <= not w24763 and not w24764;
w24766 <= b(48) and w10169;
w24767 <= b(46) and w10539;
w24768 <= b(47) and w10164;
w24769 <= not w24767 and not w24768;
w24770 <= not w24766 and w24769;
w24771 <= w7752 and w10172;
w24772 <= w24770 and not w24771;
w24773 <= a(56) and not w24772;
w24774 <= a(56) and not w24773;
w24775 <= not w24772 and not w24773;
w24776 <= not w24774 and not w24775;
w24777 <= not w24765 and not w24776;
w24778 <= not w24765 and not w24777;
w24779 <= not w24776 and not w24777;
w24780 <= not w24778 and not w24779;
w24781 <= not w24608 and not w24621;
w24782 <= w24780 and w24781;
w24783 <= not w24780 and not w24781;
w24784 <= not w24782 and not w24783;
w24785 <= b(51) and w9082;
w24786 <= b(49) and w9475;
w24787 <= b(50) and w9077;
w24788 <= not w24786 and not w24787;
w24789 <= not w24785 and w24788;
w24790 <= w8719 and w9085;
w24791 <= w24789 and not w24790;
w24792 <= a(53) and not w24791;
w24793 <= a(53) and not w24792;
w24794 <= not w24791 and not w24792;
w24795 <= not w24793 and not w24794;
w24796 <= not w24784 and w24795;
w24797 <= w24784 and not w24795;
w24798 <= not w24796 and not w24797;
w24799 <= not w24716 and w24798;
w24800 <= w24716 and not w24798;
w24801 <= not w24799 and not w24800;
w24802 <= not w24715 and w24801;
w24803 <= w24715 and not w24801;
w24804 <= not w24802 and not w24803;
w24805 <= not w24704 and w24804;
w24806 <= w24704 and not w24804;
w24807 <= not w24805 and not w24806;
w24808 <= b(57) and w7189;
w24809 <= b(55) and w7530;
w24810 <= b(56) and w7184;
w24811 <= not w24809 and not w24810;
w24812 <= not w24808 and w24811;
w24813 <= w7192 and w11153;
w24814 <= w24812 and not w24813;
w24815 <= a(47) and not w24814;
w24816 <= a(47) and not w24815;
w24817 <= not w24814 and not w24815;
w24818 <= not w24816 and not w24817;
w24819 <= w24807 and not w24818;
w24820 <= w24807 and not w24819;
w24821 <= not w24818 and not w24819;
w24822 <= not w24820 and not w24821;
w24823 <= not w24651 and not w24654;
w24824 <= w24822 and w24823;
w24825 <= not w24822 and not w24823;
w24826 <= not w24824 and not w24825;
w24827 <= b(60) and w6338;
w24828 <= b(58) and w6645;
w24829 <= b(59) and w6333;
w24830 <= not w24828 and not w24829;
w24831 <= not w24827 and w24830;
w24832 <= w6341 and w11954;
w24833 <= w24831 and not w24832;
w24834 <= a(44) and not w24833;
w24835 <= a(44) and not w24834;
w24836 <= not w24833 and not w24834;
w24837 <= not w24835 and not w24836;
w24838 <= w24826 and not w24837;
w24839 <= w24826 and not w24838;
w24840 <= not w24837 and not w24838;
w24841 <= not w24839 and not w24840;
w24842 <= not w24657 and not w24671;
w24843 <= w24841 and w24842;
w24844 <= not w24841 and not w24842;
w24845 <= not w24843 and not w24844;
w24846 <= b(63) and w5520;
w24847 <= b(61) and w5802;
w24848 <= b(62) and w5515;
w24849 <= not w24847 and not w24848;
w24850 <= not w24846 and w24849;
w24851 <= w5523 and w13514;
w24852 <= w24850 and not w24851;
w24853 <= a(41) and not w24852;
w24854 <= a(41) and not w24853;
w24855 <= not w24852 and not w24853;
w24856 <= not w24854 and not w24855;
w24857 <= w24845 and not w24856;
w24858 <= w24845 and not w24857;
w24859 <= not w24856 and not w24857;
w24860 <= not w24858 and not w24859;
w24861 <= not w24677 and not w24690;
w24862 <= w24860 and w24861;
w24863 <= not w24860 and not w24861;
w24864 <= not w24862 and not w24863;
w24865 <= not w24539 and not w24693;
w24866 <= not w24536 and not w24865;
w24867 <= w24864 and not w24866;
w24868 <= not w24864 and w24866;
w24869 <= not w24867 and not w24868;
w24870 <= not w24703 and w24869;
w24871 <= w24703 and not w24869;
w24872 <= not w24870 and not w24871;
w24873 <= not w24838 and not w24844;
w24874 <= b(62) and w5802;
w24875 <= b(63) and w5515;
w24876 <= not w24874 and not w24875;
w24877 <= not w5523 and w24876;
w24878 <= w13543 and w24876;
w24879 <= not w24877 and not w24878;
w24880 <= a(41) and not w24879;
w24881 <= not a(41) and w24879;
w24882 <= not w24880 and not w24881;
w24883 <= not w24873 and not w24882;
w24884 <= w24873 and w24882;
w24885 <= not w24883 and not w24884;
w24886 <= not w24727 and not w24741;
w24887 <= b(39) and w13646;
w24888 <= b(40) and not w13231;
w24889 <= not w24887 and not w24888;
w24890 <= not a(38) and not w24369;
w24891 <= not w24724 and not w24890;
w24892 <= w24889 and not w24891;
w24893 <= not w24889 and w24891;
w24894 <= not w24892 and not w24893;
w24895 <= b(43) and w12411;
w24896 <= b(41) and w12790;
w24897 <= b(42) and w12406;
w24898 <= not w24896 and not w24897;
w24899 <= not w24895 and w24898;
w24900 <= not w12414 and w24899;
w24901 <= not w6258 and w24899;
w24902 <= not w24900 and not w24901;
w24903 <= a(62) and not w24902;
w24904 <= not a(62) and w24902;
w24905 <= not w24903 and not w24904;
w24906 <= w24894 and not w24905;
w24907 <= not w24894 and w24905;
w24908 <= not w24906 and not w24907;
w24909 <= not w24886 and w24908;
w24910 <= w24886 and not w24908;
w24911 <= not w24909 and not w24910;
w24912 <= b(46) and w11274;
w24913 <= b(44) and w11639;
w24914 <= b(45) and w11269;
w24915 <= not w24913 and not w24914;
w24916 <= not w24912 and w24915;
w24917 <= w7420 and w11277;
w24918 <= w24916 and not w24917;
w24919 <= a(59) and not w24918;
w24920 <= a(59) and not w24919;
w24921 <= not w24918 and not w24919;
w24922 <= not w24920 and not w24921;
w24923 <= w24911 and not w24922;
w24924 <= w24911 and not w24923;
w24925 <= not w24922 and not w24923;
w24926 <= not w24924 and not w24925;
w24927 <= not w24756 and not w24762;
w24928 <= w24926 and w24927;
w24929 <= not w24926 and not w24927;
w24930 <= not w24928 and not w24929;
w24931 <= b(49) and w10169;
w24932 <= b(47) and w10539;
w24933 <= b(48) and w10164;
w24934 <= not w24932 and not w24933;
w24935 <= not w24931 and w24934;
w24936 <= w8368 and w10172;
w24937 <= w24935 and not w24936;
w24938 <= a(56) and not w24937;
w24939 <= a(56) and not w24938;
w24940 <= not w24937 and not w24938;
w24941 <= not w24939 and not w24940;
w24942 <= w24930 and not w24941;
w24943 <= w24930 and not w24942;
w24944 <= not w24941 and not w24942;
w24945 <= not w24943 and not w24944;
w24946 <= not w24777 and not w24783;
w24947 <= w24945 and w24946;
w24948 <= not w24945 and not w24946;
w24949 <= not w24947 and not w24948;
w24950 <= b(52) and w9082;
w24951 <= b(50) and w9475;
w24952 <= b(51) and w9077;
w24953 <= not w24951 and not w24952;
w24954 <= not w24950 and w24953;
w24955 <= w9085 and w9371;
w24956 <= w24954 and not w24955;
w24957 <= a(53) and not w24956;
w24958 <= a(53) and not w24957;
w24959 <= not w24956 and not w24957;
w24960 <= not w24958 and not w24959;
w24961 <= w24949 and not w24960;
w24962 <= w24949 and not w24961;
w24963 <= not w24960 and not w24961;
w24964 <= not w24962 and not w24963;
w24965 <= not w24797 and not w24799;
w24966 <= not w24964 and not w24965;
w24967 <= not w24964 and not w24966;
w24968 <= not w24965 and not w24966;
w24969 <= not w24967 and not w24968;
w24970 <= b(55) and w8105;
w24971 <= b(53) and w8458;
w24972 <= b(54) and w8100;
w24973 <= not w24971 and not w24972;
w24974 <= not w24970 and w24973;
w24975 <= w8108 and w10427;
w24976 <= w24974 and not w24975;
w24977 <= a(50) and not w24976;
w24978 <= a(50) and not w24977;
w24979 <= not w24976 and not w24977;
w24980 <= not w24978 and not w24979;
w24981 <= not w24969 and not w24980;
w24982 <= not w24969 and not w24981;
w24983 <= not w24980 and not w24981;
w24984 <= not w24982 and not w24983;
w24985 <= not w24802 and not w24805;
w24986 <= w24984 and w24985;
w24987 <= not w24984 and not w24985;
w24988 <= not w24986 and not w24987;
w24989 <= b(58) and w7189;
w24990 <= b(56) and w7530;
w24991 <= b(57) and w7184;
w24992 <= not w24990 and not w24991;
w24993 <= not w24989 and w24992;
w24994 <= w7192 and w11179;
w24995 <= w24993 and not w24994;
w24996 <= a(47) and not w24995;
w24997 <= a(47) and not w24996;
w24998 <= not w24995 and not w24996;
w24999 <= not w24997 and not w24998;
w25000 <= w24988 and not w24999;
w25001 <= w24988 and not w25000;
w25002 <= not w24999 and not w25000;
w25003 <= not w25001 and not w25002;
w25004 <= not w24819 and not w24825;
w25005 <= w25003 and w25004;
w25006 <= not w25003 and not w25004;
w25007 <= not w25005 and not w25006;
w25008 <= b(61) and w6338;
w25009 <= b(59) and w6645;
w25010 <= b(60) and w6333;
w25011 <= not w25009 and not w25010;
w25012 <= not w25008 and w25011;
w25013 <= w6341 and w12712;
w25014 <= w25012 and not w25013;
w25015 <= a(44) and not w25014;
w25016 <= a(44) and not w25015;
w25017 <= not w25014 and not w25015;
w25018 <= not w25016 and not w25017;
w25019 <= w25007 and not w25018;
w25020 <= not w25007 and w25018;
w25021 <= w24885 and not w25020;
w25022 <= not w25019 and w25021;
w25023 <= w24885 and not w25022;
w25024 <= not w25020 and not w25022;
w25025 <= not w25019 and w25024;
w25026 <= not w25023 and not w25025;
w25027 <= not w24857 and not w24863;
w25028 <= w25026 and w25027;
w25029 <= not w25026 and not w25027;
w25030 <= not w25028 and not w25029;
w25031 <= not w24867 and not w24870;
w25032 <= w25030 and not w25031;
w25033 <= not w25030 and w25031;
w25034 <= not w25032 and not w25033;
w25035 <= not w25029 and not w25032;
w25036 <= not w24883 and not w25022;
w25037 <= not w25006 and not w25019;
w25038 <= b(63) and w5802;
w25039 <= w5523 and w13540;
w25040 <= not w25038 and not w25039;
w25041 <= a(41) and not w25040;
w25042 <= a(41) and not w25041;
w25043 <= not w25040 and not w25041;
w25044 <= not w25042 and not w25043;
w25045 <= not w25037 and not w25044;
w25046 <= not w25037 and not w25045;
w25047 <= not w25044 and not w25045;
w25048 <= not w25046 and not w25047;
w25049 <= b(59) and w7189;
w25050 <= b(57) and w7530;
w25051 <= b(58) and w7184;
w25052 <= not w25050 and not w25051;
w25053 <= not w25049 and w25052;
w25054 <= w7192 and w11922;
w25055 <= w25053 and not w25054;
w25056 <= a(47) and not w25055;
w25057 <= a(47) and not w25056;
w25058 <= not w25055 and not w25056;
w25059 <= not w25057 and not w25058;
w25060 <= not w24966 and not w24981;
w25061 <= b(56) and w8105;
w25062 <= b(54) and w8458;
w25063 <= b(55) and w8100;
w25064 <= not w25062 and not w25063;
w25065 <= not w25061 and w25064;
w25066 <= w8108 and w10451;
w25067 <= w25065 and not w25066;
w25068 <= a(50) and not w25067;
w25069 <= a(50) and not w25068;
w25070 <= not w25067 and not w25068;
w25071 <= not w25069 and not w25070;
w25072 <= not w24948 and not w24961;
w25073 <= b(53) and w9082;
w25074 <= b(51) and w9475;
w25075 <= b(52) and w9077;
w25076 <= not w25074 and not w25075;
w25077 <= not w25073 and w25076;
w25078 <= w9085 and w9715;
w25079 <= w25077 and not w25078;
w25080 <= a(53) and not w25079;
w25081 <= a(53) and not w25080;
w25082 <= not w25079 and not w25080;
w25083 <= not w25081 and not w25082;
w25084 <= not w24929 and not w24942;
w25085 <= not w24909 and not w24923;
w25086 <= not w24892 and not w24906;
w25087 <= b(40) and w13646;
w25088 <= b(41) and not w13231;
w25089 <= not w25087 and not w25088;
w25090 <= w24889 and not w25089;
w25091 <= w24889 and not w25090;
w25092 <= not w25089 and not w25090;
w25093 <= not w25091 and not w25092;
w25094 <= not w25086 and not w25093;
w25095 <= not w25086 and not w25094;
w25096 <= not w25093 and not w25094;
w25097 <= not w25095 and not w25096;
w25098 <= b(44) and w12411;
w25099 <= b(42) and w12790;
w25100 <= b(43) and w12406;
w25101 <= not w25099 and not w25100;
w25102 <= not w25098 and w25101;
w25103 <= w6815 and w12414;
w25104 <= w25102 and not w25103;
w25105 <= a(62) and not w25104;
w25106 <= a(62) and not w25105;
w25107 <= not w25104 and not w25105;
w25108 <= not w25106 and not w25107;
w25109 <= not w25097 and w25108;
w25110 <= w25097 and not w25108;
w25111 <= not w25109 and not w25110;
w25112 <= b(47) and w11274;
w25113 <= b(45) and w11639;
w25114 <= b(46) and w11269;
w25115 <= not w25113 and not w25114;
w25116 <= not w25112 and w25115;
w25117 <= w7446 and w11277;
w25118 <= w25116 and not w25117;
w25119 <= a(59) and not w25118;
w25120 <= a(59) and not w25119;
w25121 <= not w25118 and not w25119;
w25122 <= not w25120 and not w25121;
w25123 <= not w25111 and not w25122;
w25124 <= w25111 and w25122;
w25125 <= not w25123 and not w25124;
w25126 <= w25085 and not w25125;
w25127 <= not w25085 and w25125;
w25128 <= not w25126 and not w25127;
w25129 <= b(50) and w10169;
w25130 <= b(48) and w10539;
w25131 <= b(49) and w10164;
w25132 <= not w25130 and not w25131;
w25133 <= not w25129 and w25132;
w25134 <= w8692 and w10172;
w25135 <= w25133 and not w25134;
w25136 <= a(56) and not w25135;
w25137 <= a(56) and not w25136;
w25138 <= not w25135 and not w25136;
w25139 <= not w25137 and not w25138;
w25140 <= not w25128 and w25139;
w25141 <= w25128 and not w25139;
w25142 <= not w25140 and not w25141;
w25143 <= not w25084 and w25142;
w25144 <= not w25084 and not w25143;
w25145 <= w25142 and not w25143;
w25146 <= not w25144 and not w25145;
w25147 <= not w25083 and not w25146;
w25148 <= w25083 and not w25145;
w25149 <= not w25144 and w25148;
w25150 <= not w25147 and not w25149;
w25151 <= not w25072 and w25150;
w25152 <= not w25072 and not w25151;
w25153 <= w25150 and not w25151;
w25154 <= not w25152 and not w25153;
w25155 <= not w25071 and not w25154;
w25156 <= w25071 and not w25153;
w25157 <= not w25152 and w25156;
w25158 <= not w25155 and not w25157;
w25159 <= not w25060 and w25158;
w25160 <= w25060 and not w25158;
w25161 <= not w25159 and not w25160;
w25162 <= not w25059 and w25161;
w25163 <= w25161 and not w25162;
w25164 <= not w25059 and not w25162;
w25165 <= not w25163 and not w25164;
w25166 <= not w24987 and not w25000;
w25167 <= w25165 and w25166;
w25168 <= not w25165 and not w25166;
w25169 <= not w25167 and not w25168;
w25170 <= b(62) and w6338;
w25171 <= b(60) and w6645;
w25172 <= b(61) and w6333;
w25173 <= not w25171 and not w25172;
w25174 <= not w25170 and w25173;
w25175 <= w6341 and w13113;
w25176 <= w25174 and not w25175;
w25177 <= a(44) and not w25176;
w25178 <= a(44) and not w25177;
w25179 <= not w25176 and not w25177;
w25180 <= not w25178 and not w25179;
w25181 <= w25169 and not w25180;
w25182 <= w25169 and not w25181;
w25183 <= not w25180 and not w25181;
w25184 <= not w25182 and not w25183;
w25185 <= not w25048 and w25184;
w25186 <= w25048 and not w25184;
w25187 <= not w25185 and not w25186;
w25188 <= not w25036 and not w25187;
w25189 <= w25036 and w25187;
w25190 <= not w25188 and not w25189;
w25191 <= not w25035 and w25190;
w25192 <= w25035 and not w25190;
w25193 <= not w25191 and not w25192;
w25194 <= not w25188 and not w25191;
w25195 <= b(60) and w7189;
w25196 <= b(58) and w7530;
w25197 <= b(59) and w7184;
w25198 <= not w25196 and not w25197;
w25199 <= not w25195 and w25198;
w25200 <= w7192 and w11954;
w25201 <= w25199 and not w25200;
w25202 <= a(47) and not w25201;
w25203 <= a(47) and not w25202;
w25204 <= not w25201 and not w25202;
w25205 <= not w25203 and not w25204;
w25206 <= not w25151 and not w25155;
w25207 <= b(57) and w8105;
w25208 <= b(55) and w8458;
w25209 <= b(56) and w8100;
w25210 <= not w25208 and not w25209;
w25211 <= not w25207 and w25210;
w25212 <= w8108 and w11153;
w25213 <= w25211 and not w25212;
w25214 <= a(50) and not w25213;
w25215 <= a(50) and not w25214;
w25216 <= not w25213 and not w25214;
w25217 <= not w25215 and not w25216;
w25218 <= not w25143 and not w25147;
w25219 <= not w25127 and not w25141;
w25220 <= b(51) and w10169;
w25221 <= b(49) and w10539;
w25222 <= b(50) and w10164;
w25223 <= not w25221 and not w25222;
w25224 <= not w25220 and w25223;
w25225 <= w8719 and w10172;
w25226 <= w25224 and not w25225;
w25227 <= a(56) and not w25226;
w25228 <= a(56) and not w25227;
w25229 <= not w25226 and not w25227;
w25230 <= not w25228 and not w25229;
w25231 <= a(41) and not w24889;
w25232 <= not a(41) and w24889;
w25233 <= not w25231 and not w25232;
w25234 <= b(41) and w13646;
w25235 <= b(42) and not w13231;
w25236 <= not w25234 and not w25235;
w25237 <= w25233 and w25236;
w25238 <= not w25233 and not w25236;
w25239 <= not w25237 and not w25238;
w25240 <= b(45) and w12411;
w25241 <= b(43) and w12790;
w25242 <= b(44) and w12406;
w25243 <= not w25241 and not w25242;
w25244 <= not w25240 and w25243;
w25245 <= w7104 and w12414;
w25246 <= w25244 and not w25245;
w25247 <= a(62) and not w25246;
w25248 <= a(62) and not w25247;
w25249 <= not w25246 and not w25247;
w25250 <= not w25248 and not w25249;
w25251 <= w25239 and not w25250;
w25252 <= w25239 and not w25251;
w25253 <= not w25250 and not w25251;
w25254 <= not w25252 and not w25253;
w25255 <= not w25090 and not w25094;
w25256 <= w25254 and w25255;
w25257 <= not w25254 and not w25255;
w25258 <= not w25256 and not w25257;
w25259 <= b(48) and w11274;
w25260 <= b(46) and w11639;
w25261 <= b(47) and w11269;
w25262 <= not w25260 and not w25261;
w25263 <= not w25259 and w25262;
w25264 <= w7752 and w11277;
w25265 <= w25263 and not w25264;
w25266 <= a(59) and not w25265;
w25267 <= a(59) and not w25266;
w25268 <= not w25265 and not w25266;
w25269 <= not w25267 and not w25268;
w25270 <= w25258 and not w25269;
w25271 <= w25258 and not w25270;
w25272 <= not w25269 and not w25270;
w25273 <= not w25271 and not w25272;
w25274 <= not w25097 and not w25108;
w25275 <= not w25123 and not w25274;
w25276 <= not w25273 and not w25275;
w25277 <= w25273 and w25275;
w25278 <= not w25276 and not w25277;
w25279 <= not w25230 and w25278;
w25280 <= not w25230 and not w25279;
w25281 <= w25278 and not w25279;
w25282 <= not w25280 and not w25281;
w25283 <= not w25219 and not w25282;
w25284 <= not w25219 and not w25283;
w25285 <= not w25282 and not w25283;
w25286 <= not w25284 and not w25285;
w25287 <= b(54) and w9082;
w25288 <= b(52) and w9475;
w25289 <= b(53) and w9077;
w25290 <= not w25288 and not w25289;
w25291 <= not w25287 and w25290;
w25292 <= w9085 and w9741;
w25293 <= w25291 and not w25292;
w25294 <= a(53) and not w25293;
w25295 <= a(53) and not w25294;
w25296 <= not w25293 and not w25294;
w25297 <= not w25295 and not w25296;
w25298 <= w25286 and w25297;
w25299 <= not w25286 and not w25297;
w25300 <= not w25298 and not w25299;
w25301 <= not w25218 and w25300;
w25302 <= w25218 and not w25300;
w25303 <= not w25301 and not w25302;
w25304 <= w25217 and not w25303;
w25305 <= not w25217 and w25303;
w25306 <= not w25304 and not w25305;
w25307 <= not w25206 and w25306;
w25308 <= w25206 and not w25306;
w25309 <= not w25307 and not w25308;
w25310 <= not w25205 and w25309;
w25311 <= w25309 and not w25310;
w25312 <= not w25205 and not w25310;
w25313 <= not w25311 and not w25312;
w25314 <= not w25159 and not w25162;
w25315 <= w25313 and w25314;
w25316 <= not w25313 and not w25314;
w25317 <= not w25315 and not w25316;
w25318 <= b(63) and w6338;
w25319 <= b(61) and w6645;
w25320 <= b(62) and w6333;
w25321 <= not w25319 and not w25320;
w25322 <= not w25318 and w25321;
w25323 <= w6341 and w13514;
w25324 <= w25322 and not w25323;
w25325 <= a(44) and not w25324;
w25326 <= a(44) and not w25325;
w25327 <= not w25324 and not w25325;
w25328 <= not w25326 and not w25327;
w25329 <= w25317 and not w25328;
w25330 <= w25317 and not w25329;
w25331 <= not w25328 and not w25329;
w25332 <= not w25330 and not w25331;
w25333 <= not w25168 and not w25181;
w25334 <= w25332 and w25333;
w25335 <= not w25332 and not w25333;
w25336 <= not w25334 and not w25335;
w25337 <= not w25048 and not w25184;
w25338 <= not w25045 and not w25337;
w25339 <= w25336 and not w25338;
w25340 <= not w25336 and w25338;
w25341 <= not w25339 and not w25340;
w25342 <= not w25194 and w25341;
w25343 <= w25194 and not w25341;
w25344 <= not w25342 and not w25343;
w25345 <= not w25310 and not w25316;
w25346 <= b(62) and w6645;
w25347 <= b(63) and w6333;
w25348 <= not w25346 and not w25347;
w25349 <= not w6341 and w25348;
w25350 <= w13543 and w25348;
w25351 <= not w25349 and not w25350;
w25352 <= a(44) and not w25351;
w25353 <= not a(44) and w25351;
w25354 <= not w25352 and not w25353;
w25355 <= not w25345 and not w25354;
w25356 <= w25345 and w25354;
w25357 <= not w25355 and not w25356;
w25358 <= b(61) and w7189;
w25359 <= b(59) and w7530;
w25360 <= b(60) and w7184;
w25361 <= not w25359 and not w25360;
w25362 <= not w25358 and w25361;
w25363 <= w7192 and w12712;
w25364 <= w25362 and not w25363;
w25365 <= a(47) and not w25364;
w25366 <= a(47) and not w25365;
w25367 <= not w25364 and not w25365;
w25368 <= not w25366 and not w25367;
w25369 <= not w25305 and not w25307;
w25370 <= not w25299 and not w25301;
w25371 <= not w25251 and not w25257;
w25372 <= b(42) and w13646;
w25373 <= b(43) and not w13231;
w25374 <= not w25372 and not w25373;
w25375 <= not a(41) and not w24889;
w25376 <= not w25238 and not w25375;
w25377 <= w25374 and not w25376;
w25378 <= w25374 and not w25377;
w25379 <= not w25376 and not w25377;
w25380 <= not w25378 and not w25379;
w25381 <= b(46) and w12411;
w25382 <= b(44) and w12790;
w25383 <= b(45) and w12406;
w25384 <= not w25382 and not w25383;
w25385 <= not w25381 and w25384;
w25386 <= not w12414 and w25385;
w25387 <= not w7420 and w25385;
w25388 <= not w25386 and not w25387;
w25389 <= a(62) and not w25388;
w25390 <= not a(62) and w25388;
w25391 <= not w25389 and not w25390;
w25392 <= not w25380 and not w25391;
w25393 <= w25380 and w25391;
w25394 <= not w25392 and not w25393;
w25395 <= not w25371 and w25394;
w25396 <= w25371 and not w25394;
w25397 <= not w25395 and not w25396;
w25398 <= b(49) and w11274;
w25399 <= b(47) and w11639;
w25400 <= b(48) and w11269;
w25401 <= not w25399 and not w25400;
w25402 <= not w25398 and w25401;
w25403 <= w8368 and w11277;
w25404 <= w25402 and not w25403;
w25405 <= a(59) and not w25404;
w25406 <= a(59) and not w25405;
w25407 <= not w25404 and not w25405;
w25408 <= not w25406 and not w25407;
w25409 <= w25397 and not w25408;
w25410 <= w25397 and not w25409;
w25411 <= not w25408 and not w25409;
w25412 <= not w25410 and not w25411;
w25413 <= not w25270 and not w25276;
w25414 <= w25412 and w25413;
w25415 <= not w25412 and not w25413;
w25416 <= not w25414 and not w25415;
w25417 <= b(52) and w10169;
w25418 <= b(50) and w10539;
w25419 <= b(51) and w10164;
w25420 <= not w25418 and not w25419;
w25421 <= not w25417 and w25420;
w25422 <= w9371 and w10172;
w25423 <= w25421 and not w25422;
w25424 <= a(56) and not w25423;
w25425 <= a(56) and not w25424;
w25426 <= not w25423 and not w25424;
w25427 <= not w25425 and not w25426;
w25428 <= w25416 and not w25427;
w25429 <= w25416 and not w25428;
w25430 <= not w25427 and not w25428;
w25431 <= not w25429 and not w25430;
w25432 <= not w25279 and not w25283;
w25433 <= w25431 and w25432;
w25434 <= not w25431 and not w25432;
w25435 <= not w25433 and not w25434;
w25436 <= b(55) and w9082;
w25437 <= b(53) and w9475;
w25438 <= b(54) and w9077;
w25439 <= not w25437 and not w25438;
w25440 <= not w25436 and w25439;
w25441 <= w9085 and w10427;
w25442 <= w25440 and not w25441;
w25443 <= a(53) and not w25442;
w25444 <= a(53) and not w25443;
w25445 <= not w25442 and not w25443;
w25446 <= not w25444 and not w25445;
w25447 <= w25435 and not w25446;
w25448 <= w25435 and not w25447;
w25449 <= not w25446 and not w25447;
w25450 <= not w25448 and not w25449;
w25451 <= not w25370 and w25450;
w25452 <= w25370 and not w25450;
w25453 <= not w25451 and not w25452;
w25454 <= b(58) and w8105;
w25455 <= b(56) and w8458;
w25456 <= b(57) and w8100;
w25457 <= not w25455 and not w25456;
w25458 <= not w25454 and w25457;
w25459 <= w8108 and w11179;
w25460 <= w25458 and not w25459;
w25461 <= a(50) and not w25460;
w25462 <= a(50) and not w25461;
w25463 <= not w25460 and not w25461;
w25464 <= not w25462 and not w25463;
w25465 <= w25453 and w25464;
w25466 <= not w25453 and not w25464;
w25467 <= not w25465 and not w25466;
w25468 <= not w25369 and w25467;
w25469 <= not w25369 and not w25468;
w25470 <= w25467 and not w25468;
w25471 <= not w25469 and not w25470;
w25472 <= not w25368 and not w25471;
w25473 <= not w25368 and not w25472;
w25474 <= not w25471 and not w25472;
w25475 <= not w25473 and not w25474;
w25476 <= w25357 and not w25475;
w25477 <= w25357 and not w25476;
w25478 <= not w25475 and not w25476;
w25479 <= not w25477 and not w25478;
w25480 <= not w25329 and not w25335;
w25481 <= w25479 and w25480;
w25482 <= not w25479 and not w25480;
w25483 <= not w25481 and not w25482;
w25484 <= not w25339 and not w25342;
w25485 <= w25483 and not w25484;
w25486 <= not w25483 and w25484;
w25487 <= not w25485 and not w25486;
w25488 <= not w25482 and not w25485;
w25489 <= not w25355 and not w25476;
w25490 <= not w25468 and not w25472;
w25491 <= b(63) and w6645;
w25492 <= w6341 and w13540;
w25493 <= not w25491 and not w25492;
w25494 <= a(44) and not w25493;
w25495 <= a(44) and not w25494;
w25496 <= not w25493 and not w25494;
w25497 <= not w25495 and not w25496;
w25498 <= not w25490 and not w25497;
w25499 <= not w25490 and not w25498;
w25500 <= not w25497 and not w25498;
w25501 <= not w25499 and not w25500;
w25502 <= b(59) and w8105;
w25503 <= b(57) and w8458;
w25504 <= b(58) and w8100;
w25505 <= not w25503 and not w25504;
w25506 <= not w25502 and w25505;
w25507 <= w8108 and w11922;
w25508 <= w25506 and not w25507;
w25509 <= a(50) and not w25508;
w25510 <= a(50) and not w25509;
w25511 <= not w25508 and not w25509;
w25512 <= not w25510 and not w25511;
w25513 <= not w25434 and not w25447;
w25514 <= b(56) and w9082;
w25515 <= b(54) and w9475;
w25516 <= b(55) and w9077;
w25517 <= not w25515 and not w25516;
w25518 <= not w25514 and w25517;
w25519 <= w9085 and w10451;
w25520 <= w25518 and not w25519;
w25521 <= a(53) and not w25520;
w25522 <= a(53) and not w25521;
w25523 <= not w25520 and not w25521;
w25524 <= not w25522 and not w25523;
w25525 <= not w25415 and not w25428;
w25526 <= b(53) and w10169;
w25527 <= b(51) and w10539;
w25528 <= b(52) and w10164;
w25529 <= not w25527 and not w25528;
w25530 <= not w25526 and w25529;
w25531 <= w9715 and w10172;
w25532 <= w25530 and not w25531;
w25533 <= a(56) and not w25532;
w25534 <= a(56) and not w25533;
w25535 <= not w25532 and not w25533;
w25536 <= not w25534 and not w25535;
w25537 <= not w25395 and not w25409;
w25538 <= b(50) and w11274;
w25539 <= b(48) and w11639;
w25540 <= b(49) and w11269;
w25541 <= not w25539 and not w25540;
w25542 <= not w25538 and w25541;
w25543 <= w8692 and w11277;
w25544 <= w25542 and not w25543;
w25545 <= a(59) and not w25544;
w25546 <= a(59) and not w25545;
w25547 <= not w25544 and not w25545;
w25548 <= not w25546 and not w25547;
w25549 <= not w25377 and not w25392;
w25550 <= b(43) and w13646;
w25551 <= b(44) and not w13231;
w25552 <= not w25550 and not w25551;
w25553 <= w25374 and not w25552;
w25554 <= not w25374 and w25552;
w25555 <= not w25553 and not w25554;
w25556 <= b(47) and w12411;
w25557 <= b(45) and w12790;
w25558 <= b(46) and w12406;
w25559 <= not w25557 and not w25558;
w25560 <= not w25556 and w25559;
w25561 <= not w12414 and w25560;
w25562 <= not w7446 and w25560;
w25563 <= not w25561 and not w25562;
w25564 <= a(62) and not w25563;
w25565 <= not a(62) and w25563;
w25566 <= not w25564 and not w25565;
w25567 <= w25555 and not w25566;
w25568 <= not w25555 and w25566;
w25569 <= not w25567 and not w25568;
w25570 <= not w25549 and w25569;
w25571 <= not w25549 and not w25570;
w25572 <= w25569 and not w25570;
w25573 <= not w25571 and not w25572;
w25574 <= not w25548 and not w25573;
w25575 <= w25548 and not w25572;
w25576 <= not w25571 and w25575;
w25577 <= not w25574 and not w25576;
w25578 <= not w25537 and w25577;
w25579 <= not w25537 and not w25578;
w25580 <= w25577 and not w25578;
w25581 <= not w25579 and not w25580;
w25582 <= not w25536 and not w25581;
w25583 <= w25536 and not w25580;
w25584 <= not w25579 and w25583;
w25585 <= not w25582 and not w25584;
w25586 <= not w25525 and w25585;
w25587 <= not w25525 and not w25586;
w25588 <= w25585 and not w25586;
w25589 <= not w25587 and not w25588;
w25590 <= not w25524 and not w25589;
w25591 <= w25524 and not w25588;
w25592 <= not w25587 and w25591;
w25593 <= not w25590 and not w25592;
w25594 <= not w25513 and w25593;
w25595 <= w25513 and not w25593;
w25596 <= not w25594 and not w25595;
w25597 <= not w25512 and w25596;
w25598 <= w25596 and not w25597;
w25599 <= not w25512 and not w25597;
w25600 <= not w25598 and not w25599;
w25601 <= not w25370 and not w25450;
w25602 <= not w25466 and not w25601;
w25603 <= not w25600 and not w25602;
w25604 <= not w25600 and not w25603;
w25605 <= not w25602 and not w25603;
w25606 <= not w25604 and not w25605;
w25607 <= b(62) and w7189;
w25608 <= b(60) and w7530;
w25609 <= b(61) and w7184;
w25610 <= not w25608 and not w25609;
w25611 <= not w25607 and w25610;
w25612 <= w7192 and w13113;
w25613 <= w25611 and not w25612;
w25614 <= a(47) and not w25613;
w25615 <= a(47) and not w25614;
w25616 <= not w25613 and not w25614;
w25617 <= not w25615 and not w25616;
w25618 <= not w25606 and not w25617;
w25619 <= not w25606 and not w25618;
w25620 <= not w25617 and not w25618;
w25621 <= not w25619 and not w25620;
w25622 <= not w25501 and w25621;
w25623 <= w25501 and not w25621;
w25624 <= not w25622 and not w25623;
w25625 <= not w25489 and not w25624;
w25626 <= w25489 and w25624;
w25627 <= not w25625 and not w25626;
w25628 <= not w25488 and w25627;
w25629 <= w25488 and not w25627;
w25630 <= not w25628 and not w25629;
w25631 <= not w25625 and not w25628;
w25632 <= b(63) and w7189;
w25633 <= b(61) and w7530;
w25634 <= b(62) and w7184;
w25635 <= not w25633 and not w25634;
w25636 <= not w25632 and w25635;
w25637 <= w7192 and w13514;
w25638 <= w25636 and not w25637;
w25639 <= a(47) and not w25638;
w25640 <= a(47) and not w25639;
w25641 <= not w25638 and not w25639;
w25642 <= not w25640 and not w25641;
w25643 <= not w25594 and not w25597;
w25644 <= b(60) and w8105;
w25645 <= b(58) and w8458;
w25646 <= b(59) and w8100;
w25647 <= not w25645 and not w25646;
w25648 <= not w25644 and w25647;
w25649 <= w8108 and w11954;
w25650 <= w25648 and not w25649;
w25651 <= a(50) and not w25650;
w25652 <= a(50) and not w25651;
w25653 <= not w25650 and not w25651;
w25654 <= not w25652 and not w25653;
w25655 <= not w25586 and not w25590;
w25656 <= b(57) and w9082;
w25657 <= b(55) and w9475;
w25658 <= b(56) and w9077;
w25659 <= not w25657 and not w25658;
w25660 <= not w25656 and w25659;
w25661 <= w9085 and w11153;
w25662 <= w25660 and not w25661;
w25663 <= a(53) and not w25662;
w25664 <= a(53) and not w25663;
w25665 <= not w25662 and not w25663;
w25666 <= not w25664 and not w25665;
w25667 <= not w25578 and not w25582;
w25668 <= b(54) and w10169;
w25669 <= b(52) and w10539;
w25670 <= b(53) and w10164;
w25671 <= not w25669 and not w25670;
w25672 <= not w25668 and w25671;
w25673 <= w9741 and w10172;
w25674 <= w25672 and not w25673;
w25675 <= a(56) and not w25674;
w25676 <= a(56) and not w25675;
w25677 <= not w25674 and not w25675;
w25678 <= not w25676 and not w25677;
w25679 <= not w25570 and not w25574;
w25680 <= not w25553 and not w25567;
w25681 <= b(44) and w13646;
w25682 <= b(45) and not w13231;
w25683 <= not w25681 and not w25682;
w25684 <= not a(44) and not w25683;
w25685 <= a(44) and w25683;
w25686 <= not w25684 and not w25685;
w25687 <= not w25374 and w25686;
w25688 <= not w25374 and not w25687;
w25689 <= w25686 and not w25687;
w25690 <= not w25688 and not w25689;
w25691 <= not w25680 and not w25690;
w25692 <= not w25680 and not w25691;
w25693 <= not w25690 and not w25691;
w25694 <= not w25692 and not w25693;
w25695 <= b(48) and w12411;
w25696 <= b(46) and w12790;
w25697 <= b(47) and w12406;
w25698 <= not w25696 and not w25697;
w25699 <= not w25695 and w25698;
w25700 <= w7752 and w12414;
w25701 <= w25699 and not w25700;
w25702 <= a(62) and not w25701;
w25703 <= a(62) and not w25702;
w25704 <= not w25701 and not w25702;
w25705 <= not w25703 and not w25704;
w25706 <= not w25694 and not w25705;
w25707 <= not w25694 and not w25706;
w25708 <= not w25705 and not w25706;
w25709 <= not w25707 and not w25708;
w25710 <= b(51) and w11274;
w25711 <= b(49) and w11639;
w25712 <= b(50) and w11269;
w25713 <= not w25711 and not w25712;
w25714 <= not w25710 and w25713;
w25715 <= w8719 and w11277;
w25716 <= w25714 and not w25715;
w25717 <= a(59) and not w25716;
w25718 <= a(59) and not w25717;
w25719 <= not w25716 and not w25717;
w25720 <= not w25718 and not w25719;
w25721 <= w25709 and w25720;
w25722 <= not w25709 and not w25720;
w25723 <= not w25721 and not w25722;
w25724 <= not w25679 and w25723;
w25725 <= w25679 and not w25723;
w25726 <= not w25724 and not w25725;
w25727 <= w25678 and not w25726;
w25728 <= not w25678 and w25726;
w25729 <= not w25727 and not w25728;
w25730 <= not w25667 and w25729;
w25731 <= w25667 and not w25729;
w25732 <= not w25730 and not w25731;
w25733 <= w25666 and not w25732;
w25734 <= not w25666 and w25732;
w25735 <= not w25733 and not w25734;
w25736 <= not w25655 and w25735;
w25737 <= w25655 and not w25735;
w25738 <= not w25736 and not w25737;
w25739 <= w25654 and not w25738;
w25740 <= not w25654 and w25738;
w25741 <= not w25739 and not w25740;
w25742 <= not w25643 and w25741;
w25743 <= w25643 and not w25741;
w25744 <= not w25742 and not w25743;
w25745 <= not w25642 and w25744;
w25746 <= w25744 and not w25745;
w25747 <= not w25642 and not w25745;
w25748 <= not w25746 and not w25747;
w25749 <= not w25603 and not w25618;
w25750 <= w25748 and w25749;
w25751 <= not w25748 and not w25749;
w25752 <= not w25750 and not w25751;
w25753 <= not w25501 and not w25621;
w25754 <= not w25498 and not w25753;
w25755 <= w25752 and not w25754;
w25756 <= not w25752 and w25754;
w25757 <= not w25755 and not w25756;
w25758 <= not w25631 and w25757;
w25759 <= w25631 and not w25757;
w25760 <= not w25758 and not w25759;
w25761 <= not w25740 and not w25742;
w25762 <= b(62) and w7530;
w25763 <= b(63) and w7184;
w25764 <= not w25762 and not w25763;
w25765 <= not w7192 and w25764;
w25766 <= w13543 and w25764;
w25767 <= not w25765 and not w25766;
w25768 <= a(47) and not w25767;
w25769 <= not a(47) and w25767;
w25770 <= not w25768 and not w25769;
w25771 <= not w25761 and not w25770;
w25772 <= w25761 and w25770;
w25773 <= not w25771 and not w25772;
w25774 <= b(61) and w8105;
w25775 <= b(59) and w8458;
w25776 <= b(60) and w8100;
w25777 <= not w25775 and not w25776;
w25778 <= not w25774 and w25777;
w25779 <= w8108 and w12712;
w25780 <= w25778 and not w25779;
w25781 <= a(50) and not w25780;
w25782 <= a(50) and not w25781;
w25783 <= not w25780 and not w25781;
w25784 <= not w25782 and not w25783;
w25785 <= not w25734 and not w25736;
w25786 <= not w25728 and not w25730;
w25787 <= b(55) and w10169;
w25788 <= b(53) and w10539;
w25789 <= b(54) and w10164;
w25790 <= not w25788 and not w25789;
w25791 <= not w25787 and w25790;
w25792 <= w10172 and w10427;
w25793 <= w25791 and not w25792;
w25794 <= a(56) and not w25793;
w25795 <= a(56) and not w25794;
w25796 <= not w25793 and not w25794;
w25797 <= not w25795 and not w25796;
w25798 <= not w25722 and not w25724;
w25799 <= b(52) and w11274;
w25800 <= b(50) and w11639;
w25801 <= b(51) and w11269;
w25802 <= not w25800 and not w25801;
w25803 <= not w25799 and w25802;
w25804 <= w9371 and w11277;
w25805 <= w25803 and not w25804;
w25806 <= a(59) and not w25805;
w25807 <= a(59) and not w25806;
w25808 <= not w25805 and not w25806;
w25809 <= not w25807 and not w25808;
w25810 <= not w25691 and not w25706;
w25811 <= b(45) and w13646;
w25812 <= b(46) and not w13231;
w25813 <= not w25811 and not w25812;
w25814 <= not w25684 and not w25687;
w25815 <= not w25813 and w25814;
w25816 <= w25813 and not w25814;
w25817 <= not w25815 and not w25816;
w25818 <= b(49) and w12411;
w25819 <= b(47) and w12790;
w25820 <= b(48) and w12406;
w25821 <= not w25819 and not w25820;
w25822 <= not w25818 and w25821;
w25823 <= w8368 and w12414;
w25824 <= w25822 and not w25823;
w25825 <= a(62) and not w25824;
w25826 <= a(62) and not w25825;
w25827 <= not w25824 and not w25825;
w25828 <= not w25826 and not w25827;
w25829 <= not w25817 and w25828;
w25830 <= w25817 and not w25828;
w25831 <= not w25829 and not w25830;
w25832 <= not w25810 and w25831;
w25833 <= not w25810 and not w25832;
w25834 <= w25831 and not w25832;
w25835 <= not w25833 and not w25834;
w25836 <= not w25809 and not w25835;
w25837 <= w25809 and not w25834;
w25838 <= not w25833 and w25837;
w25839 <= not w25836 and not w25838;
w25840 <= not w25798 and w25839;
w25841 <= w25798 and not w25839;
w25842 <= not w25840 and not w25841;
w25843 <= not w25797 and w25842;
w25844 <= w25842 and not w25843;
w25845 <= not w25797 and not w25843;
w25846 <= not w25844 and not w25845;
w25847 <= not w25786 and w25846;
w25848 <= w25786 and not w25846;
w25849 <= not w25847 and not w25848;
w25850 <= b(58) and w9082;
w25851 <= b(56) and w9475;
w25852 <= b(57) and w9077;
w25853 <= not w25851 and not w25852;
w25854 <= not w25850 and w25853;
w25855 <= w9085 and w11179;
w25856 <= w25854 and not w25855;
w25857 <= a(53) and not w25856;
w25858 <= a(53) and not w25857;
w25859 <= not w25856 and not w25857;
w25860 <= not w25858 and not w25859;
w25861 <= w25849 and w25860;
w25862 <= not w25849 and not w25860;
w25863 <= not w25861 and not w25862;
w25864 <= not w25785 and w25863;
w25865 <= not w25785 and not w25864;
w25866 <= w25863 and not w25864;
w25867 <= not w25865 and not w25866;
w25868 <= not w25784 and not w25867;
w25869 <= not w25784 and not w25868;
w25870 <= not w25867 and not w25868;
w25871 <= not w25869 and not w25870;
w25872 <= w25773 and not w25871;
w25873 <= w25773 and not w25872;
w25874 <= not w25871 and not w25872;
w25875 <= not w25873 and not w25874;
w25876 <= not w25745 and not w25751;
w25877 <= w25875 and w25876;
w25878 <= not w25875 and not w25876;
w25879 <= not w25877 and not w25878;
w25880 <= not w25755 and not w25758;
w25881 <= w25879 and not w25880;
w25882 <= not w25879 and w25880;
w25883 <= not w25881 and not w25882;
w25884 <= b(59) and w9082;
w25885 <= b(57) and w9475;
w25886 <= b(58) and w9077;
w25887 <= not w25885 and not w25886;
w25888 <= not w25884 and w25887;
w25889 <= w9085 and w11922;
w25890 <= w25888 and not w25889;
w25891 <= a(53) and not w25890;
w25892 <= a(53) and not w25891;
w25893 <= not w25890 and not w25891;
w25894 <= not w25892 and not w25893;
w25895 <= not w25840 and not w25843;
w25896 <= b(56) and w10169;
w25897 <= b(54) and w10539;
w25898 <= b(55) and w10164;
w25899 <= not w25897 and not w25898;
w25900 <= not w25896 and w25899;
w25901 <= w10172 and w10451;
w25902 <= w25900 and not w25901;
w25903 <= a(56) and not w25902;
w25904 <= a(56) and not w25903;
w25905 <= not w25902 and not w25903;
w25906 <= not w25904 and not w25905;
w25907 <= not w25832 and not w25836;
w25908 <= b(53) and w11274;
w25909 <= b(51) and w11639;
w25910 <= b(52) and w11269;
w25911 <= not w25909 and not w25910;
w25912 <= not w25908 and w25911;
w25913 <= w9715 and w11277;
w25914 <= w25912 and not w25913;
w25915 <= a(59) and not w25914;
w25916 <= a(59) and not w25915;
w25917 <= not w25914 and not w25915;
w25918 <= not w25916 and not w25917;
w25919 <= not w25816 and not w25830;
w25920 <= b(46) and w13646;
w25921 <= b(47) and not w13231;
w25922 <= not w25920 and not w25921;
w25923 <= w25813 and not w25922;
w25924 <= not w25813 and w25922;
w25925 <= not w25919 and not w25924;
w25926 <= not w25923 and w25925;
w25927 <= not w25919 and not w25926;
w25928 <= not w25924 and not w25926;
w25929 <= not w25923 and w25928;
w25930 <= not w25927 and not w25929;
w25931 <= b(50) and w12411;
w25932 <= b(48) and w12790;
w25933 <= b(49) and w12406;
w25934 <= not w25932 and not w25933;
w25935 <= not w25931 and w25934;
w25936 <= w8692 and w12414;
w25937 <= w25935 and not w25936;
w25938 <= a(62) and not w25937;
w25939 <= a(62) and not w25938;
w25940 <= not w25937 and not w25938;
w25941 <= not w25939 and not w25940;
w25942 <= not w25930 and w25941;
w25943 <= w25930 and not w25941;
w25944 <= not w25942 and not w25943;
w25945 <= not w25918 and not w25944;
w25946 <= w25918 and w25944;
w25947 <= not w25945 and not w25946;
w25948 <= not w25907 and w25947;
w25949 <= not w25907 and not w25948;
w25950 <= w25947 and not w25948;
w25951 <= not w25949 and not w25950;
w25952 <= not w25906 and not w25951;
w25953 <= w25906 and not w25950;
w25954 <= not w25949 and w25953;
w25955 <= not w25952 and not w25954;
w25956 <= not w25895 and w25955;
w25957 <= w25895 and not w25955;
w25958 <= not w25956 and not w25957;
w25959 <= not w25894 and w25958;
w25960 <= w25958 and not w25959;
w25961 <= not w25894 and not w25959;
w25962 <= not w25960 and not w25961;
w25963 <= not w25786 and not w25846;
w25964 <= not w25862 and not w25963;
w25965 <= not w25962 and not w25964;
w25966 <= not w25962 and not w25965;
w25967 <= not w25964 and not w25965;
w25968 <= not w25966 and not w25967;
w25969 <= b(62) and w8105;
w25970 <= b(60) and w8458;
w25971 <= b(61) and w8100;
w25972 <= not w25970 and not w25971;
w25973 <= not w25969 and w25972;
w25974 <= w8108 and w13113;
w25975 <= w25973 and not w25974;
w25976 <= a(50) and not w25975;
w25977 <= a(50) and not w25976;
w25978 <= not w25975 and not w25976;
w25979 <= not w25977 and not w25978;
w25980 <= not w25968 and not w25979;
w25981 <= not w25968 and not w25980;
w25982 <= not w25979 and not w25980;
w25983 <= not w25981 and not w25982;
w25984 <= not w25864 and not w25868;
w25985 <= b(63) and w7530;
w25986 <= not w7192 and not w25985;
w25987 <= not w13540 and not w25985;
w25988 <= not w25986 and not w25987;
w25989 <= a(47) and not w25988;
w25990 <= not a(47) and w25988;
w25991 <= not w25989 and not w25990;
w25992 <= not w25984 and not w25991;
w25993 <= w25984 and w25991;
w25994 <= not w25992 and not w25993;
w25995 <= not w25983 and w25994;
w25996 <= not w25983 and not w25995;
w25997 <= w25994 and not w25995;
w25998 <= not w25996 and not w25997;
w25999 <= not w25771 and not w25872;
w26000 <= w25998 and w25999;
w26001 <= not w25998 and not w25999;
w26002 <= not w26000 and not w26001;
w26003 <= not w25878 and not w25881;
w26004 <= w26002 and not w26003;
w26005 <= not w26002 and w26003;
w26006 <= not w26004 and not w26005;
w26007 <= b(63) and w8105;
w26008 <= b(61) and w8458;
w26009 <= b(62) and w8100;
w26010 <= not w26008 and not w26009;
w26011 <= not w26007 and w26010;
w26012 <= w8108 and w13514;
w26013 <= w26011 and not w26012;
w26014 <= a(50) and not w26013;
w26015 <= a(50) and not w26014;
w26016 <= not w26013 and not w26014;
w26017 <= not w26015 and not w26016;
w26018 <= not w25956 and not w25959;
w26019 <= b(60) and w9082;
w26020 <= b(58) and w9475;
w26021 <= b(59) and w9077;
w26022 <= not w26020 and not w26021;
w26023 <= not w26019 and w26022;
w26024 <= w9085 and w11954;
w26025 <= w26023 and not w26024;
w26026 <= a(53) and not w26025;
w26027 <= a(53) and not w26026;
w26028 <= not w26025 and not w26026;
w26029 <= not w26027 and not w26028;
w26030 <= not w25948 and not w25952;
w26031 <= b(57) and w10169;
w26032 <= b(55) and w10539;
w26033 <= b(56) and w10164;
w26034 <= not w26032 and not w26033;
w26035 <= not w26031 and w26034;
w26036 <= w10172 and w11153;
w26037 <= w26035 and not w26036;
w26038 <= a(56) and not w26037;
w26039 <= a(56) and not w26038;
w26040 <= not w26037 and not w26038;
w26041 <= not w26039 and not w26040;
w26042 <= not w25930 and not w25941;
w26043 <= not w25945 and not w26042;
w26044 <= b(51) and w12411;
w26045 <= b(49) and w12790;
w26046 <= b(50) and w12406;
w26047 <= not w26045 and not w26046;
w26048 <= not w26044 and w26047;
w26049 <= w8719 and w12414;
w26050 <= w26048 and not w26049;
w26051 <= a(62) and not w26050;
w26052 <= a(62) and not w26051;
w26053 <= not w26050 and not w26051;
w26054 <= not w26052 and not w26053;
w26055 <= b(47) and w13646;
w26056 <= b(48) and not w13231;
w26057 <= not w26055 and not w26056;
w26058 <= a(47) and not w25922;
w26059 <= not a(47) and w25922;
w26060 <= not w26058 and not w26059;
w26061 <= not w26057 and not w26060;
w26062 <= w26057 and w26060;
w26063 <= not w26061 and not w26062;
w26064 <= not w26054 and w26063;
w26065 <= not w26054 and not w26064;
w26066 <= w26063 and not w26064;
w26067 <= not w26065 and not w26066;
w26068 <= not w25928 and not w26067;
w26069 <= not w25928 and not w26068;
w26070 <= not w26067 and not w26068;
w26071 <= not w26069 and not w26070;
w26072 <= b(54) and w11274;
w26073 <= b(52) and w11639;
w26074 <= b(53) and w11269;
w26075 <= not w26073 and not w26074;
w26076 <= not w26072 and w26075;
w26077 <= w9741 and w11277;
w26078 <= w26076 and not w26077;
w26079 <= a(59) and not w26078;
w26080 <= a(59) and not w26079;
w26081 <= not w26078 and not w26079;
w26082 <= not w26080 and not w26081;
w26083 <= w26071 and w26082;
w26084 <= not w26071 and not w26082;
w26085 <= not w26083 and not w26084;
w26086 <= not w26043 and w26085;
w26087 <= w26043 and not w26085;
w26088 <= not w26086 and not w26087;
w26089 <= w26041 and not w26088;
w26090 <= not w26041 and w26088;
w26091 <= not w26089 and not w26090;
w26092 <= not w26030 and w26091;
w26093 <= w26030 and not w26091;
w26094 <= not w26092 and not w26093;
w26095 <= w26029 and not w26094;
w26096 <= not w26029 and w26094;
w26097 <= not w26095 and not w26096;
w26098 <= not w26018 and w26097;
w26099 <= w26018 and not w26097;
w26100 <= not w26098 and not w26099;
w26101 <= not w26017 and w26100;
w26102 <= w26100 and not w26101;
w26103 <= not w26017 and not w26101;
w26104 <= not w26102 and not w26103;
w26105 <= not w25965 and not w25980;
w26106 <= w26104 and w26105;
w26107 <= not w26104 and not w26105;
w26108 <= not w26106 and not w26107;
w26109 <= not w25992 and not w25995;
w26110 <= not w26108 and w26109;
w26111 <= w26108 and not w26109;
w26112 <= not w26110 and not w26111;
w26113 <= not w26001 and not w26004;
w26114 <= w26112 and not w26113;
w26115 <= not w26112 and w26113;
w26116 <= not w26114 and not w26115;
w26117 <= b(62) and w8458;
w26118 <= b(63) and w8100;
w26119 <= not w26117 and not w26118;
w26120 <= w8108 and not w13543;
w26121 <= w26119 and not w26120;
w26122 <= a(50) and not w26121;
w26123 <= a(50) and not w26122;
w26124 <= not w26121 and not w26122;
w26125 <= not w26123 and not w26124;
w26126 <= not w26096 and not w26098;
w26127 <= b(61) and w9082;
w26128 <= b(59) and w9475;
w26129 <= b(60) and w9077;
w26130 <= not w26128 and not w26129;
w26131 <= not w26127 and w26130;
w26132 <= w9085 and w12712;
w26133 <= w26131 and not w26132;
w26134 <= a(53) and not w26133;
w26135 <= a(53) and not w26134;
w26136 <= not w26133 and not w26134;
w26137 <= not w26135 and not w26136;
w26138 <= not w26090 and not w26092;
w26139 <= b(58) and w10169;
w26140 <= b(56) and w10539;
w26141 <= b(57) and w10164;
w26142 <= not w26140 and not w26141;
w26143 <= not w26139 and w26142;
w26144 <= w10172 and w11179;
w26145 <= w26143 and not w26144;
w26146 <= a(56) and not w26145;
w26147 <= a(56) and not w26146;
w26148 <= not w26145 and not w26146;
w26149 <= not w26147 and not w26148;
w26150 <= not w26084 and not w26086;
w26151 <= b(55) and w11274;
w26152 <= b(53) and w11639;
w26153 <= b(54) and w11269;
w26154 <= not w26152 and not w26153;
w26155 <= not w26151 and w26154;
w26156 <= w10427 and w11277;
w26157 <= w26155 and not w26156;
w26158 <= a(59) and not w26157;
w26159 <= a(59) and not w26158;
w26160 <= not w26157 and not w26158;
w26161 <= not w26159 and not w26160;
w26162 <= not w26064 and not w26068;
w26163 <= b(48) and w13646;
w26164 <= b(49) and not w13231;
w26165 <= not w26163 and not w26164;
w26166 <= not a(47) and not w25922;
w26167 <= not w26061 and not w26166;
w26168 <= w26165 and not w26167;
w26169 <= not w26165 and w26167;
w26170 <= not w26168 and not w26169;
w26171 <= b(52) and w12411;
w26172 <= b(50) and w12790;
w26173 <= b(51) and w12406;
w26174 <= not w26172 and not w26173;
w26175 <= not w26171 and w26174;
w26176 <= not w12414 and w26175;
w26177 <= not w9371 and w26175;
w26178 <= not w26176 and not w26177;
w26179 <= a(62) and not w26178;
w26180 <= not a(62) and w26178;
w26181 <= not w26179 and not w26180;
w26182 <= w26170 and not w26181;
w26183 <= not w26170 and w26181;
w26184 <= not w26182 and not w26183;
w26185 <= not w26162 and w26184;
w26186 <= not w26162 and not w26185;
w26187 <= w26184 and not w26185;
w26188 <= not w26186 and not w26187;
w26189 <= not w26161 and not w26188;
w26190 <= w26161 and not w26187;
w26191 <= not w26186 and w26190;
w26192 <= not w26189 and not w26191;
w26193 <= not w26150 and w26192;
w26194 <= w26150 and not w26192;
w26195 <= not w26193 and not w26194;
w26196 <= not w26149 and w26195;
w26197 <= w26149 and not w26195;
w26198 <= not w26196 and not w26197;
w26199 <= not w26138 and w26198;
w26200 <= not w26138 and not w26199;
w26201 <= w26198 and not w26199;
w26202 <= not w26200 and not w26201;
w26203 <= not w26137 and not w26202;
w26204 <= w26137 and not w26201;
w26205 <= not w26200 and w26204;
w26206 <= not w26203 and not w26205;
w26207 <= not w26126 and w26206;
w26208 <= w26126 and not w26206;
w26209 <= not w26207 and not w26208;
w26210 <= not w26125 and w26209;
w26211 <= w26209 and not w26210;
w26212 <= not w26125 and not w26210;
w26213 <= not w26211 and not w26212;
w26214 <= not w26101 and not w26107;
w26215 <= w26213 and w26214;
w26216 <= not w26213 and not w26214;
w26217 <= not w26215 and not w26216;
w26218 <= not w26111 and not w26114;
w26219 <= w26217 and not w26218;
w26220 <= not w26217 and w26218;
w26221 <= not w26219 and not w26220;
w26222 <= b(59) and w10169;
w26223 <= b(57) and w10539;
w26224 <= b(58) and w10164;
w26225 <= not w26223 and not w26224;
w26226 <= not w26222 and w26225;
w26227 <= w10172 and w11922;
w26228 <= w26226 and not w26227;
w26229 <= a(56) and not w26228;
w26230 <= a(56) and not w26229;
w26231 <= not w26228 and not w26229;
w26232 <= not w26230 and not w26231;
w26233 <= not w26185 and not w26189;
w26234 <= b(53) and w12411;
w26235 <= b(51) and w12790;
w26236 <= b(52) and w12406;
w26237 <= not w26235 and not w26236;
w26238 <= not w26234 and w26237;
w26239 <= w9715 and w12414;
w26240 <= w26238 and not w26239;
w26241 <= a(62) and not w26240;
w26242 <= a(62) and not w26241;
w26243 <= not w26240 and not w26241;
w26244 <= not w26242 and not w26243;
w26245 <= b(49) and w13646;
w26246 <= b(50) and not w13231;
w26247 <= not w26245 and not w26246;
w26248 <= w26165 and not w26247;
w26249 <= w26165 and not w26248;
w26250 <= not w26247 and not w26248;
w26251 <= not w26249 and not w26250;
w26252 <= not w26244 and not w26251;
w26253 <= not w26244 and not w26252;
w26254 <= not w26251 and not w26252;
w26255 <= not w26253 and not w26254;
w26256 <= not w26168 and not w26182;
w26257 <= w26255 and w26256;
w26258 <= not w26255 and not w26256;
w26259 <= not w26257 and not w26258;
w26260 <= b(56) and w11274;
w26261 <= b(54) and w11639;
w26262 <= b(55) and w11269;
w26263 <= not w26261 and not w26262;
w26264 <= not w26260 and w26263;
w26265 <= w10451 and w11277;
w26266 <= w26264 and not w26265;
w26267 <= a(59) and not w26266;
w26268 <= a(59) and not w26267;
w26269 <= not w26266 and not w26267;
w26270 <= not w26268 and not w26269;
w26271 <= not w26259 and w26270;
w26272 <= w26259 and not w26270;
w26273 <= not w26271 and not w26272;
w26274 <= not w26233 and w26273;
w26275 <= w26233 and not w26273;
w26276 <= not w26274 and not w26275;
w26277 <= not w26232 and w26276;
w26278 <= w26276 and not w26277;
w26279 <= not w26232 and not w26277;
w26280 <= not w26278 and not w26279;
w26281 <= not w26193 and not w26196;
w26282 <= w26280 and w26281;
w26283 <= not w26280 and not w26281;
w26284 <= not w26282 and not w26283;
w26285 <= b(62) and w9082;
w26286 <= b(60) and w9475;
w26287 <= b(61) and w9077;
w26288 <= not w26286 and not w26287;
w26289 <= not w26285 and w26288;
w26290 <= w9085 and w13113;
w26291 <= w26289 and not w26290;
w26292 <= a(53) and not w26291;
w26293 <= a(53) and not w26292;
w26294 <= not w26291 and not w26292;
w26295 <= not w26293 and not w26294;
w26296 <= w26284 and not w26295;
w26297 <= w26284 and not w26296;
w26298 <= not w26295 and not w26296;
w26299 <= not w26297 and not w26298;
w26300 <= not w26199 and not w26203;
w26301 <= b(63) and w8458;
w26302 <= not w8108 and not w26301;
w26303 <= not w13540 and not w26301;
w26304 <= not w26302 and not w26303;
w26305 <= a(50) and not w26304;
w26306 <= not a(50) and w26304;
w26307 <= not w26305 and not w26306;
w26308 <= not w26300 and not w26307;
w26309 <= w26300 and w26307;
w26310 <= not w26308 and not w26309;
w26311 <= not w26299 and w26310;
w26312 <= not w26299 and not w26311;
w26313 <= w26310 and not w26311;
w26314 <= not w26312 and not w26313;
w26315 <= not w26207 and not w26210;
w26316 <= w26314 and w26315;
w26317 <= not w26314 and not w26315;
w26318 <= not w26316 and not w26317;
w26319 <= not w26216 and not w26219;
w26320 <= w26318 and not w26319;
w26321 <= not w26318 and w26319;
w26322 <= not w26320 and not w26321;
w26323 <= not w26274 and not w26277;
w26324 <= b(60) and w10169;
w26325 <= b(58) and w10539;
w26326 <= b(59) and w10164;
w26327 <= not w26325 and not w26326;
w26328 <= not w26324 and w26327;
w26329 <= w10172 and w11954;
w26330 <= w26328 and not w26329;
w26331 <= a(56) and not w26330;
w26332 <= a(56) and not w26331;
w26333 <= not w26330 and not w26331;
w26334 <= not w26332 and not w26333;
w26335 <= not w26258 and not w26272;
w26336 <= b(57) and w11274;
w26337 <= b(55) and w11639;
w26338 <= b(56) and w11269;
w26339 <= not w26337 and not w26338;
w26340 <= not w26336 and w26339;
w26341 <= w11153 and w11277;
w26342 <= w26340 and not w26341;
w26343 <= a(59) and not w26342;
w26344 <= a(59) and not w26343;
w26345 <= not w26342 and not w26343;
w26346 <= not w26344 and not w26345;
w26347 <= b(54) and w12411;
w26348 <= b(52) and w12790;
w26349 <= b(53) and w12406;
w26350 <= not w26348 and not w26349;
w26351 <= not w26347 and w26350;
w26352 <= w9741 and w12414;
w26353 <= w26351 and not w26352;
w26354 <= a(62) and not w26353;
w26355 <= a(62) and not w26354;
w26356 <= not w26353 and not w26354;
w26357 <= not w26355 and not w26356;
w26358 <= not w26248 and not w26252;
w26359 <= b(50) and w13646;
w26360 <= b(51) and not w13231;
w26361 <= not w26359 and not w26360;
w26362 <= not a(50) and not w26361;
w26363 <= a(50) and w26361;
w26364 <= not w26362 and not w26363;
w26365 <= not w26165 and w26364;
w26366 <= w26165 and not w26364;
w26367 <= not w26365 and not w26366;
w26368 <= not w26358 and w26367;
w26369 <= not w26358 and not w26368;
w26370 <= w26367 and not w26368;
w26371 <= not w26369 and not w26370;
w26372 <= not w26357 and not w26371;
w26373 <= w26357 and not w26370;
w26374 <= not w26369 and w26373;
w26375 <= not w26372 and not w26374;
w26376 <= not w26346 and w26375;
w26377 <= not w26346 and not w26376;
w26378 <= w26375 and not w26376;
w26379 <= not w26377 and not w26378;
w26380 <= not w26335 and not w26379;
w26381 <= w26335 and not w26378;
w26382 <= not w26377 and w26381;
w26383 <= not w26380 and not w26382;
w26384 <= not w26334 and w26383;
w26385 <= w26334 and not w26383;
w26386 <= not w26384 and not w26385;
w26387 <= not w26323 and w26386;
w26388 <= w26323 and not w26386;
w26389 <= not w26387 and not w26388;
w26390 <= b(63) and w9082;
w26391 <= b(61) and w9475;
w26392 <= b(62) and w9077;
w26393 <= not w26391 and not w26392;
w26394 <= not w26390 and w26393;
w26395 <= w9085 and w13514;
w26396 <= w26394 and not w26395;
w26397 <= a(53) and not w26396;
w26398 <= a(53) and not w26397;
w26399 <= not w26396 and not w26397;
w26400 <= not w26398 and not w26399;
w26401 <= w26389 and not w26400;
w26402 <= w26389 and not w26401;
w26403 <= not w26400 and not w26401;
w26404 <= not w26402 and not w26403;
w26405 <= not w26283 and not w26296;
w26406 <= w26404 and w26405;
w26407 <= not w26404 and not w26405;
w26408 <= not w26406 and not w26407;
w26409 <= not w26308 and not w26311;
w26410 <= not w26408 and w26409;
w26411 <= w26408 and not w26409;
w26412 <= not w26410 and not w26411;
w26413 <= not w26317 and not w26320;
w26414 <= w26412 and not w26413;
w26415 <= not w26412 and w26413;
w26416 <= not w26414 and not w26415;
w26417 <= b(62) and w9475;
w26418 <= b(63) and w9077;
w26419 <= not w26417 and not w26418;
w26420 <= w9085 and not w13543;
w26421 <= w26419 and not w26420;
w26422 <= a(53) and not w26421;
w26423 <= a(53) and not w26422;
w26424 <= not w26421 and not w26422;
w26425 <= not w26423 and not w26424;
w26426 <= not w26384 and not w26387;
w26427 <= b(61) and w10169;
w26428 <= b(59) and w10539;
w26429 <= b(60) and w10164;
w26430 <= not w26428 and not w26429;
w26431 <= not w26427 and w26430;
w26432 <= w10172 and w12712;
w26433 <= w26431 and not w26432;
w26434 <= a(56) and not w26433;
w26435 <= a(56) and not w26434;
w26436 <= not w26433 and not w26434;
w26437 <= not w26435 and not w26436;
w26438 <= not w26376 and not w26380;
w26439 <= b(58) and w11274;
w26440 <= b(56) and w11639;
w26441 <= b(57) and w11269;
w26442 <= not w26440 and not w26441;
w26443 <= not w26439 and w26442;
w26444 <= w11179 and w11277;
w26445 <= w26443 and not w26444;
w26446 <= a(59) and not w26445;
w26447 <= a(59) and not w26446;
w26448 <= not w26445 and not w26446;
w26449 <= not w26447 and not w26448;
w26450 <= not w26368 and not w26372;
w26451 <= b(51) and w13646;
w26452 <= b(52) and not w13231;
w26453 <= not w26451 and not w26452;
w26454 <= not w26362 and not w26365;
w26455 <= not w26453 and w26454;
w26456 <= w26453 and not w26454;
w26457 <= not w26455 and not w26456;
w26458 <= b(55) and w12411;
w26459 <= b(53) and w12790;
w26460 <= b(54) and w12406;
w26461 <= not w26459 and not w26460;
w26462 <= not w26458 and w26461;
w26463 <= w10427 and w12414;
w26464 <= w26462 and not w26463;
w26465 <= a(62) and not w26464;
w26466 <= a(62) and not w26465;
w26467 <= not w26464 and not w26465;
w26468 <= not w26466 and not w26467;
w26469 <= not w26457 and w26468;
w26470 <= w26457 and not w26468;
w26471 <= not w26469 and not w26470;
w26472 <= not w26450 and w26471;
w26473 <= w26450 and not w26471;
w26474 <= not w26472 and not w26473;
w26475 <= not w26449 and w26474;
w26476 <= w26449 and not w26474;
w26477 <= not w26475 and not w26476;
w26478 <= not w26438 and w26477;
w26479 <= not w26438 and not w26478;
w26480 <= w26477 and not w26478;
w26481 <= not w26479 and not w26480;
w26482 <= not w26437 and not w26481;
w26483 <= w26437 and not w26480;
w26484 <= not w26479 and w26483;
w26485 <= not w26482 and not w26484;
w26486 <= not w26426 and w26485;
w26487 <= w26426 and not w26485;
w26488 <= not w26486 and not w26487;
w26489 <= not w26425 and w26488;
w26490 <= w26488 and not w26489;
w26491 <= not w26425 and not w26489;
w26492 <= not w26490 and not w26491;
w26493 <= not w26401 and not w26407;
w26494 <= w26492 and w26493;
w26495 <= not w26492 and not w26493;
w26496 <= not w26494 and not w26495;
w26497 <= not w26411 and not w26414;
w26498 <= w26496 and not w26497;
w26499 <= not w26496 and w26497;
w26500 <= not w26498 and not w26499;
w26501 <= not w26472 and not w26475;
w26502 <= not w26456 and not w26470;
w26503 <= b(52) and w13646;
w26504 <= b(53) and not w13231;
w26505 <= not w26503 and not w26504;
w26506 <= w26453 and not w26505;
w26507 <= not w26453 and w26505;
w26508 <= not w26502 and not w26507;
w26509 <= not w26506 and w26508;
w26510 <= not w26502 and not w26509;
w26511 <= not w26507 and not w26509;
w26512 <= not w26506 and w26511;
w26513 <= not w26510 and not w26512;
w26514 <= b(56) and w12411;
w26515 <= b(54) and w12790;
w26516 <= b(55) and w12406;
w26517 <= not w26515 and not w26516;
w26518 <= not w26514 and w26517;
w26519 <= w10451 and w12414;
w26520 <= w26518 and not w26519;
w26521 <= a(62) and not w26520;
w26522 <= a(62) and not w26521;
w26523 <= not w26520 and not w26521;
w26524 <= not w26522 and not w26523;
w26525 <= not w26513 and w26524;
w26526 <= w26513 and not w26524;
w26527 <= not w26525 and not w26526;
w26528 <= b(59) and w11274;
w26529 <= b(57) and w11639;
w26530 <= b(58) and w11269;
w26531 <= not w26529 and not w26530;
w26532 <= not w26528 and w26531;
w26533 <= w11277 and w11922;
w26534 <= w26532 and not w26533;
w26535 <= a(59) and not w26534;
w26536 <= a(59) and not w26535;
w26537 <= not w26534 and not w26535;
w26538 <= not w26536 and not w26537;
w26539 <= not w26527 and not w26538;
w26540 <= w26527 and w26538;
w26541 <= not w26539 and not w26540;
w26542 <= w26501 and not w26541;
w26543 <= not w26501 and w26541;
w26544 <= not w26542 and not w26543;
w26545 <= b(62) and w10169;
w26546 <= b(60) and w10539;
w26547 <= b(61) and w10164;
w26548 <= not w26546 and not w26547;
w26549 <= not w26545 and w26548;
w26550 <= w10172 and w13113;
w26551 <= w26549 and not w26550;
w26552 <= a(56) and not w26551;
w26553 <= a(56) and not w26552;
w26554 <= not w26551 and not w26552;
w26555 <= not w26553 and not w26554;
w26556 <= w26544 and not w26555;
w26557 <= w26544 and not w26556;
w26558 <= not w26555 and not w26556;
w26559 <= not w26557 and not w26558;
w26560 <= not w26478 and not w26482;
w26561 <= b(63) and w9475;
w26562 <= not w9085 and not w26561;
w26563 <= not w13540 and not w26561;
w26564 <= not w26562 and not w26563;
w26565 <= a(53) and not w26564;
w26566 <= not a(53) and w26564;
w26567 <= not w26565 and not w26566;
w26568 <= not w26560 and not w26567;
w26569 <= w26560 and w26567;
w26570 <= not w26568 and not w26569;
w26571 <= not w26559 and w26570;
w26572 <= not w26559 and not w26571;
w26573 <= w26570 and not w26571;
w26574 <= not w26572 and not w26573;
w26575 <= not w26486 and not w26489;
w26576 <= w26574 and w26575;
w26577 <= not w26574 and not w26575;
w26578 <= not w26576 and not w26577;
w26579 <= not w26495 and not w26498;
w26580 <= w26578 and not w26579;
w26581 <= not w26578 and w26579;
w26582 <= not w26580 and not w26581;
w26583 <= not w26577 and not w26580;
w26584 <= not w26568 and not w26571;
w26585 <= not w26543 and not w26556;
w26586 <= b(63) and w10169;
w26587 <= b(61) and w10539;
w26588 <= b(62) and w10164;
w26589 <= not w26587 and not w26588;
w26590 <= not w26586 and w26589;
w26591 <= w10172 and w13514;
w26592 <= w26590 and not w26591;
w26593 <= a(56) and not w26592;
w26594 <= a(56) and not w26593;
w26595 <= not w26592 and not w26593;
w26596 <= not w26594 and not w26595;
w26597 <= not w26585 and not w26596;
w26598 <= not w26585 and not w26597;
w26599 <= not w26596 and not w26597;
w26600 <= not w26598 and not w26599;
w26601 <= not w26513 and not w26524;
w26602 <= not w26539 and not w26601;
w26603 <= b(60) and w11274;
w26604 <= b(58) and w11639;
w26605 <= b(59) and w11269;
w26606 <= not w26604 and not w26605;
w26607 <= not w26603 and w26606;
w26608 <= w11277 and w11954;
w26609 <= w26607 and not w26608;
w26610 <= a(59) and not w26609;
w26611 <= a(59) and not w26610;
w26612 <= not w26609 and not w26610;
w26613 <= not w26611 and not w26612;
w26614 <= a(53) and not w26505;
w26615 <= not a(53) and w26505;
w26616 <= not w26614 and not w26615;
w26617 <= b(53) and w13646;
w26618 <= b(54) and not w13231;
w26619 <= not w26617 and not w26618;
w26620 <= w26616 and w26619;
w26621 <= not w26616 and not w26619;
w26622 <= not w26620 and not w26621;
w26623 <= b(57) and w12411;
w26624 <= b(55) and w12790;
w26625 <= b(56) and w12406;
w26626 <= not w26624 and not w26625;
w26627 <= not w26623 and w26626;
w26628 <= w11153 and w12414;
w26629 <= w26627 and not w26628;
w26630 <= a(62) and not w26629;
w26631 <= a(62) and not w26630;
w26632 <= not w26629 and not w26630;
w26633 <= not w26631 and not w26632;
w26634 <= w26622 and not w26633;
w26635 <= w26622 and not w26634;
w26636 <= not w26633 and not w26634;
w26637 <= not w26635 and not w26636;
w26638 <= not w26511 and not w26637;
w26639 <= w26511 and w26637;
w26640 <= not w26638 and not w26639;
w26641 <= not w26613 and w26640;
w26642 <= not w26613 and not w26641;
w26643 <= w26640 and not w26641;
w26644 <= not w26642 and not w26643;
w26645 <= not w26602 and not w26644;
w26646 <= not w26602 and not w26645;
w26647 <= not w26644 and not w26645;
w26648 <= not w26646 and not w26647;
w26649 <= not w26600 and w26648;
w26650 <= w26600 and not w26648;
w26651 <= not w26649 and not w26650;
w26652 <= not w26584 and not w26651;
w26653 <= w26584 and w26651;
w26654 <= not w26652 and not w26653;
w26655 <= not w26583 and w26654;
w26656 <= w26583 and not w26654;
w26657 <= not w26655 and not w26656;
w26658 <= b(62) and w10539;
w26659 <= b(63) and w10164;
w26660 <= not w26658 and not w26659;
w26661 <= w10172 and not w13543;
w26662 <= w26660 and not w26661;
w26663 <= a(56) and not w26662;
w26664 <= a(56) and not w26663;
w26665 <= not w26662 and not w26663;
w26666 <= not w26664 and not w26665;
w26667 <= not w26641 and not w26645;
w26668 <= b(61) and w11274;
w26669 <= b(59) and w11639;
w26670 <= b(60) and w11269;
w26671 <= not w26669 and not w26670;
w26672 <= not w26668 and w26671;
w26673 <= w11277 and w12712;
w26674 <= w26672 and not w26673;
w26675 <= a(59) and not w26674;
w26676 <= a(59) and not w26675;
w26677 <= not w26674 and not w26675;
w26678 <= not w26676 and not w26677;
w26679 <= not w26634 and not w26638;
w26680 <= b(54) and w13646;
w26681 <= b(55) and not w13231;
w26682 <= not w26680 and not w26681;
w26683 <= not a(53) and not w26505;
w26684 <= not w26621 and not w26683;
w26685 <= w26682 and not w26684;
w26686 <= not w26682 and w26684;
w26687 <= not w26685 and not w26686;
w26688 <= b(58) and w12411;
w26689 <= b(56) and w12790;
w26690 <= b(57) and w12406;
w26691 <= not w26689 and not w26690;
w26692 <= not w26688 and w26691;
w26693 <= not w12414 and w26692;
w26694 <= not w11179 and w26692;
w26695 <= not w26693 and not w26694;
w26696 <= a(62) and not w26695;
w26697 <= not a(62) and w26695;
w26698 <= not w26696 and not w26697;
w26699 <= w26687 and not w26698;
w26700 <= not w26687 and w26698;
w26701 <= not w26699 and not w26700;
w26702 <= not w26679 and w26701;
w26703 <= not w26679 and not w26702;
w26704 <= w26701 and not w26702;
w26705 <= not w26703 and not w26704;
w26706 <= not w26678 and not w26705;
w26707 <= w26678 and not w26704;
w26708 <= not w26703 and w26707;
w26709 <= not w26706 and not w26708;
w26710 <= not w26667 and w26709;
w26711 <= w26667 and not w26709;
w26712 <= not w26710 and not w26711;
w26713 <= not w26666 and w26712;
w26714 <= w26712 and not w26713;
w26715 <= not w26666 and not w26713;
w26716 <= not w26714 and not w26715;
w26717 <= not w26600 and not w26648;
w26718 <= not w26597 and not w26717;
w26719 <= not w26716 and not w26718;
w26720 <= not w26716 and not w26719;
w26721 <= not w26718 and not w26719;
w26722 <= not w26720 and not w26721;
w26723 <= not w26652 and not w26655;
w26724 <= not w26722 and not w26723;
w26725 <= w26722 and w26723;
w26726 <= not w26724 and not w26725;
w26727 <= b(59) and w12411;
w26728 <= b(57) and w12790;
w26729 <= b(58) and w12406;
w26730 <= not w26728 and not w26729;
w26731 <= not w26727 and w26730;
w26732 <= w11922 and w12414;
w26733 <= w26731 and not w26732;
w26734 <= a(62) and not w26733;
w26735 <= a(62) and not w26734;
w26736 <= not w26733 and not w26734;
w26737 <= not w26735 and not w26736;
w26738 <= b(55) and w13646;
w26739 <= b(56) and not w13231;
w26740 <= not w26738 and not w26739;
w26741 <= w26682 and not w26740;
w26742 <= w26682 and not w26741;
w26743 <= not w26740 and not w26741;
w26744 <= not w26742 and not w26743;
w26745 <= not w26737 and not w26744;
w26746 <= not w26737 and not w26745;
w26747 <= not w26744 and not w26745;
w26748 <= not w26746 and not w26747;
w26749 <= not w26685 and not w26699;
w26750 <= w26748 and w26749;
w26751 <= not w26748 and not w26749;
w26752 <= not w26750 and not w26751;
w26753 <= b(62) and w11274;
w26754 <= b(60) and w11639;
w26755 <= b(61) and w11269;
w26756 <= not w26754 and not w26755;
w26757 <= not w26753 and w26756;
w26758 <= w11277 and w13113;
w26759 <= w26757 and not w26758;
w26760 <= a(59) and not w26759;
w26761 <= a(59) and not w26760;
w26762 <= not w26759 and not w26760;
w26763 <= not w26761 and not w26762;
w26764 <= w26752 and not w26763;
w26765 <= w26752 and not w26764;
w26766 <= not w26763 and not w26764;
w26767 <= not w26765 and not w26766;
w26768 <= not w26702 and not w26706;
w26769 <= b(63) and w10539;
w26770 <= not w10172 and not w26769;
w26771 <= not w13540 and not w26769;
w26772 <= not w26770 and not w26771;
w26773 <= a(56) and not w26772;
w26774 <= not a(56) and w26772;
w26775 <= not w26773 and not w26774;
w26776 <= not w26768 and not w26775;
w26777 <= w26768 and w26775;
w26778 <= not w26776 and not w26777;
w26779 <= not w26767 and w26778;
w26780 <= not w26767 and not w26779;
w26781 <= w26778 and not w26779;
w26782 <= not w26780 and not w26781;
w26783 <= not w26710 and not w26713;
w26784 <= w26782 and w26783;
w26785 <= not w26782 and not w26783;
w26786 <= not w26784 and not w26785;
w26787 <= not w26719 and not w26724;
w26788 <= w26786 and not w26787;
w26789 <= not w26786 and w26787;
w26790 <= not w26788 and not w26789;
w26791 <= not w26751 and not w26764;
w26792 <= b(63) and w11274;
w26793 <= b(61) and w11639;
w26794 <= b(62) and w11269;
w26795 <= not w26793 and not w26794;
w26796 <= not w26792 and w26795;
w26797 <= w11277 and w13514;
w26798 <= w26796 and not w26797;
w26799 <= a(59) and not w26798;
w26800 <= a(59) and not w26799;
w26801 <= not w26798 and not w26799;
w26802 <= not w26800 and not w26801;
w26803 <= not w26791 and not w26802;
w26804 <= not w26791 and not w26803;
w26805 <= not w26802 and not w26803;
w26806 <= not w26804 and not w26805;
w26807 <= b(56) and w13646;
w26808 <= b(57) and not w13231;
w26809 <= not w26807 and not w26808;
w26810 <= not a(56) and not w26809;
w26811 <= not a(56) and not w26810;
w26812 <= not w26809 and not w26810;
w26813 <= not w26811 and not w26812;
w26814 <= not w26682 and not w26813;
w26815 <= not w26682 and not w26814;
w26816 <= not w26813 and not w26814;
w26817 <= not w26815 and not w26816;
w26818 <= not w26741 and not w26745;
w26819 <= w26817 and w26818;
w26820 <= not w26817 and not w26818;
w26821 <= not w26819 and not w26820;
w26822 <= b(60) and w12411;
w26823 <= b(58) and w12790;
w26824 <= b(59) and w12406;
w26825 <= not w26823 and not w26824;
w26826 <= not w26822 and w26825;
w26827 <= w11954 and w12414;
w26828 <= w26826 and not w26827;
w26829 <= a(62) and not w26828;
w26830 <= a(62) and not w26829;
w26831 <= not w26828 and not w26829;
w26832 <= not w26830 and not w26831;
w26833 <= w26821 and not w26832;
w26834 <= not w26821 and w26832;
w26835 <= not w26806 and not w26834;
w26836 <= not w26833 and w26835;
w26837 <= not w26806 and not w26836;
w26838 <= not w26834 and not w26836;
w26839 <= not w26833 and w26838;
w26840 <= not w26837 and not w26839;
w26841 <= not w26776 and not w26779;
w26842 <= w26840 and w26841;
w26843 <= not w26840 and not w26841;
w26844 <= not w26842 and not w26843;
w26845 <= not w26785 and not w26788;
w26846 <= w26844 and not w26845;
w26847 <= not w26844 and w26845;
w26848 <= not w26846 and not w26847;
w26849 <= not w26820 and not w26833;
w26850 <= b(57) and w13646;
w26851 <= b(58) and not w13231;
w26852 <= not w26850 and not w26851;
w26853 <= not w26810 and not w26814;
w26854 <= not w26852 and w26853;
w26855 <= w26852 and not w26853;
w26856 <= not w26854 and not w26855;
w26857 <= b(61) and w12411;
w26858 <= b(59) and w12790;
w26859 <= b(60) and w12406;
w26860 <= not w26858 and not w26859;
w26861 <= not w26857 and w26860;
w26862 <= not w12414 and w26861;
w26863 <= not w12712 and w26861;
w26864 <= not w26862 and not w26863;
w26865 <= a(62) and not w26864;
w26866 <= not a(62) and w26864;
w26867 <= not w26865 and not w26866;
w26868 <= w26856 and not w26867;
w26869 <= not w26856 and w26867;
w26870 <= not w26868 and not w26869;
w26871 <= not w26849 and w26870;
w26872 <= w26849 and not w26870;
w26873 <= not w26871 and not w26872;
w26874 <= b(62) and w11639;
w26875 <= b(63) and w11269;
w26876 <= not w26874 and not w26875;
w26877 <= w11277 and not w13543;
w26878 <= w26876 and not w26877;
w26879 <= a(59) and not w26878;
w26880 <= a(59) and not w26879;
w26881 <= not w26878 and not w26879;
w26882 <= not w26880 and not w26881;
w26883 <= w26873 and not w26882;
w26884 <= w26873 and not w26883;
w26885 <= not w26882 and not w26883;
w26886 <= not w26884 and not w26885;
w26887 <= not w26803 and not w26836;
w26888 <= w26886 and w26887;
w26889 <= not w26886 and not w26887;
w26890 <= not w26888 and not w26889;
w26891 <= not w26843 and not w26846;
w26892 <= w26890 and not w26891;
w26893 <= not w26890 and w26891;
w26894 <= not w26892 and not w26893;
w26895 <= not w26889 and not w26892;
w26896 <= not w26871 and not w26883;
w26897 <= not w26855 and not w26868;
w26898 <= b(58) and w13646;
w26899 <= b(59) and not w13231;
w26900 <= not w26898 and not w26899;
w26901 <= w26852 and not w26900;
w26902 <= not w26852 and w26900;
w26903 <= not w26897 and not w26902;
w26904 <= not w26901 and w26903;
w26905 <= not w26897 and not w26904;
w26906 <= not w26902 and not w26904;
w26907 <= not w26901 and w26906;
w26908 <= not w26905 and not w26907;
w26909 <= b(62) and w12411;
w26910 <= b(60) and w12790;
w26911 <= b(61) and w12406;
w26912 <= not w26910 and not w26911;
w26913 <= not w26909 and w26912;
w26914 <= w12414 and w13113;
w26915 <= w26913 and not w26914;
w26916 <= a(62) and not w26915;
w26917 <= a(62) and not w26916;
w26918 <= not w26915 and not w26916;
w26919 <= not w26917 and not w26918;
w26920 <= b(63) and w11639;
w26921 <= w11277 and w13540;
w26922 <= not w26920 and not w26921;
w26923 <= a(59) and not w26922;
w26924 <= a(59) and not w26923;
w26925 <= not w26922 and not w26923;
w26926 <= not w26924 and not w26925;
w26927 <= not w26919 and not w26926;
w26928 <= not w26919 and not w26927;
w26929 <= not w26926 and not w26927;
w26930 <= not w26928 and not w26929;
w26931 <= not w26908 and w26930;
w26932 <= w26908 and not w26930;
w26933 <= not w26931 and not w26932;
w26934 <= not w26896 and not w26933;
w26935 <= not w26896 and not w26934;
w26936 <= not w26933 and not w26934;
w26937 <= not w26935 and not w26936;
w26938 <= not w26895 and not w26937;
w26939 <= w26895 and not w26936;
w26940 <= not w26935 and w26939;
w26941 <= not w26938 and not w26940;
w26942 <= not w26934 and not w26938;
w26943 <= not w26908 and not w26930;
w26944 <= not w26927 and not w26943;
w26945 <= a(59) and not w26900;
w26946 <= not a(59) and w26900;
w26947 <= not w26945 and not w26946;
w26948 <= b(59) and w13646;
w26949 <= b(60) and not w13231;
w26950 <= not w26948 and not w26949;
w26951 <= w26947 and w26950;
w26952 <= not w26947 and not w26950;
w26953 <= not w26951 and not w26952;
w26954 <= b(63) and w12411;
w26955 <= b(61) and w12790;
w26956 <= b(62) and w12406;
w26957 <= not w26955 and not w26956;
w26958 <= not w26954 and w26957;
w26959 <= w12414 and w13514;
w26960 <= w26958 and not w26959;
w26961 <= a(62) and not w26960;
w26962 <= a(62) and not w26961;
w26963 <= not w26960 and not w26961;
w26964 <= not w26962 and not w26963;
w26965 <= w26953 and not w26964;
w26966 <= w26953 and not w26965;
w26967 <= not w26964 and not w26965;
w26968 <= not w26966 and not w26967;
w26969 <= not w26906 and not w26968;
w26970 <= w26906 and w26968;
w26971 <= not w26969 and not w26970;
w26972 <= not w26944 and w26971;
w26973 <= not w26944 and not w26972;
w26974 <= w26971 and not w26972;
w26975 <= not w26973 and not w26974;
w26976 <= not w26942 and not w26975;
w26977 <= w26942 and not w26974;
w26978 <= not w26973 and w26977;
w26979 <= not w26976 and not w26978;
w26980 <= not w26972 and not w26976;
w26981 <= not w26965 and not w26969;
w26982 <= b(60) and w13646;
w26983 <= b(61) and not w13231;
w26984 <= not w26982 and not w26983;
w26985 <= not a(59) and not w26900;
w26986 <= not w26952 and not w26985;
w26987 <= w26984 and not w26986;
w26988 <= not w26984 and w26986;
w26989 <= not w26987 and not w26988;
w26990 <= b(62) and w12790;
w26991 <= b(63) and w12406;
w26992 <= not w26990 and not w26991;
w26993 <= not w12414 and w26992;
w26994 <= w13543 and w26992;
w26995 <= not w26993 and not w26994;
w26996 <= a(62) and not w26995;
w26997 <= not a(62) and w26995;
w26998 <= not w26996 and not w26997;
w26999 <= w26989 and not w26998;
w27000 <= not w26989 and w26998;
w27001 <= not w26999 and not w27000;
w27002 <= not w26981 and w27001;
w27003 <= not w26981 and not w27002;
w27004 <= w27001 and not w27002;
w27005 <= not w27003 and not w27004;
w27006 <= not w26980 and not w27005;
w27007 <= w26980 and not w27004;
w27008 <= not w27003 and w27007;
w27009 <= not w27006 and not w27008;
w27010 <= not w27002 and not w27006;
w27011 <= not w26987 and not w26999;
w27012 <= b(61) and w13646;
w27013 <= b(62) and not w13231;
w27014 <= not w27012 and not w27013;
w27015 <= w26984 and not w27014;
w27016 <= not w26984 and w27014;
w27017 <= not w27015 and not w27016;
w27018 <= b(63) and w12790;
w27019 <= not w12414 and not w27018;
w27020 <= not w13540 and not w27018;
w27021 <= not w27019 and not w27020;
w27022 <= a(62) and not w27021;
w27023 <= not a(62) and w27021;
w27024 <= not w27022 and not w27023;
w27025 <= w27017 and not w27024;
w27026 <= not w27017 and w27024;
w27027 <= not w27025 and not w27026;
w27028 <= not w27011 and w27027;
w27029 <= not w27011 and not w27028;
w27030 <= w27027 and not w27028;
w27031 <= not w27029 and not w27030;
w27032 <= not w27010 and not w27031;
w27033 <= w27010 and not w27030;
w27034 <= not w27029 and w27033;
w27035 <= not w27032 and not w27034;
w27036 <= not w27028 and not w27032;
w27037 <= not w27015 and not w27025;
w27038 <= b(62) and w13646;
w27039 <= b(63) and not w13231;
w27040 <= not w27038 and not w27039;
w27041 <= not a(62) and not w27040;
w27042 <= a(62) and w27040;
w27043 <= not w27041 and not w27042;
w27044 <= not w26984 and w27043;
w27045 <= w26984 and not w27043;
w27046 <= not w27044 and not w27045;
w27047 <= not w27037 and w27046;
w27048 <= w27037 and not w27046;
w27049 <= not w27047 and not w27048;
w27050 <= not w27036 and w27049;
w27051 <= w27036 and not w27049;
w27052 <= not w27050 and not w27051;
w27053 <= not w27041 and not w27044;
w27054 <= b(63) and w13646;
w27055 <= not w27053 and w27054;
w27056 <= w27053 and not w27054;
w27057 <= not w27055 and not w27056;
w27058 <= not w27047 and not w27050;
w27059 <= w27057 and w27058;
w27060 <= not w27057 and not w27058;
w27061 <= not w27059 and not w27060;
one <= '1';
f(0) <= w3;-- level 3
f(1) <= w24;-- level 11
f(2) <= w48;-- level 13
f(3) <= w77;-- level 15
f(4) <= w125;-- level 17
f(5) <= w167;-- level 19
f(6) <= w214;-- level 21
f(7) <= w281;-- level 23
f(8) <= w342;-- level 26
f(9) <= w408;-- level 28
f(10) <= w493;-- level 30
f(11) <= w573;-- level 32
f(12) <= w658;-- level 34
f(13) <= w763;-- level 38
f(14) <= w860;-- level 40
f(15) <= w967;-- level 43
f(16) <= w1087;-- level 44
f(17) <= w1204;-- level 46
f(18) <= w1323;-- level 48
f(19) <= w1465;-- level 50
f(20) <= w1603;-- level 52
f(21) <= w1741;-- level 54
f(22) <= w1900;-- level 56
f(23) <= w2057;-- level 58
f(24) <= w2215;-- level 60
f(25) <= w2394;-- level 62
f(26) <= w2568;-- level 64
f(27) <= w2745;-- level 66
f(28) <= w2944;-- level 68
f(29) <= w3140;-- level 70
f(30) <= w3334;-- level 72
f(31) <= w3553;-- level 74
f(32) <= w3768;-- level 77
f(33) <= w3978;-- level 79
f(34) <= w4221;-- level 82
f(35) <= w4451;-- level 85
f(36) <= w4680;-- level 87
f(37) <= w4936;-- level 89
f(38) <= w5182;-- level 91
f(39) <= w5433;-- level 93
f(40) <= w5710;-- level 95
f(41) <= w5974;-- level 97
f(42) <= w6246;-- level 99
f(43) <= w6544;-- level 101
f(44) <= w6827;-- level 103
f(45) <= w7116;-- level 105
f(46) <= w7434;-- level 108
f(47) <= w7739;-- level 110
f(48) <= w8044;-- level 112
f(49) <= w8380;-- level 114
f(50) <= w8706;-- level 118
f(51) <= w9028;-- level 120
f(52) <= w9383;-- level 122
f(53) <= w9727;-- level 126
f(54) <= w10071;-- level 128
f(55) <= w10439;-- level 130
f(56) <= w10802;-- level 132
f(57) <= w11167;-- level 134
f(58) <= w11556;-- level 136
f(59) <= w11939;-- level 139
f(60) <= w12322;-- level 140
f(61) <= w12730;-- level 142
f(62) <= w13128;-- level 144
f(63) <= w13533;-- level 146
f(64) <= w13936;-- level 148
f(65) <= w14334;-- level 150
f(66) <= w14723;-- level 152
f(67) <= w15119;-- level 155
f(68) <= w15510;-- level 157
f(69) <= w15888;-- level 158
f(70) <= w16260;-- level 160
f(71) <= w16633;-- level 163
f(72) <= w16997;-- level 165
f(73) <= w17362;-- level 167
f(74) <= w17713;-- level 169
f(75) <= w18059;-- level 171
f(76) <= w18405;-- level 173
f(77) <= w18731;-- level 174
f(78) <= w19056;-- level 176
f(79) <= w19371;-- level 178
f(80) <= w19682;-- level 181
f(81) <= w19984;-- level 183
f(82) <= w20282;-- level 185
f(83) <= w20568;-- level 186
f(84) <= w20855;-- level 188
f(85) <= w21129;-- level 190
f(86) <= w21400;-- level 193
f(87) <= w21666;-- level 195
f(88) <= w21926;-- level 197
f(89) <= w22175;-- level 198
f(90) <= w22418;-- level 200
f(91) <= w22655;-- level 202
f(92) <= w22890;-- level 205
f(93) <= w23116;-- level 206
f(94) <= w23336;-- level 208
f(95) <= w23552;-- level 211
f(96) <= w23760;-- level 212
f(97) <= w23959;-- level 214
f(98) <= w24155;-- level 216
f(99) <= w24342;-- level 218
f(100) <= w24525;-- level 220
f(101) <= w24702;-- level 222
f(102) <= w24872;-- level 224
f(103) <= w25034;-- level 226
f(104) <= w25193;-- level 228
f(105) <= w25344;-- level 230
f(106) <= w25487;-- level 232
f(107) <= w25630;-- level 234
f(108) <= w25760;-- level 236
f(109) <= w25883;-- level 238
f(110) <= w26006;-- level 240
f(111) <= w26116;-- level 242
f(112) <= w26221;-- level 244
f(113) <= w26322;-- level 246
f(114) <= w26416;-- level 248
f(115) <= w26500;-- level 250
f(116) <= w26582;-- level 252
f(117) <= w26657;-- level 254
f(118) <= w26726;-- level 256
f(119) <= w26790;-- level 258
f(120) <= w26848;-- level 260
f(121) <= w26894;-- level 262
f(122) <= w26941;-- level 265
f(123) <= w26979;-- level 267
f(124) <= w27009;-- level 269
f(125) <= w27035;-- level 271
f(126) <= w27052;-- level 272
f(127) <= w27061;-- level 274
end Behavioral;