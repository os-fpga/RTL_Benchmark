// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_bpu_bht (
    core_clk,
    core_reset_n,
    bht_update_p0,
    bht_update_p0_dir_addr,
    bht_update_p0_sel_addr,
    bht_update_p0_sel_data,
    bht_update_p0_dir_data,
    bht_update_p1,
    bht_update_p1_dir_addr,
    bht_update_p1_sel_addr,
    bht_update_p1_sel_data,
    bht_update_p1_dir_data,
    bht_dir_rd_addr,
    bht_sel_rd_addr,
    bht_taken_rdata,
    bht_ntaken_rdata,
    bht_sel_rdata
);
parameter BTB_SIZE = 256;
input core_clk;
input core_reset_n;
input bht_update_p0;
input [7:0] bht_update_p0_dir_addr;
input [7:0] bht_update_p0_sel_addr;
input [1:0] bht_update_p0_sel_data;
input [1:0] bht_update_p0_dir_data;
input bht_update_p1;
input [7:0] bht_update_p1_dir_addr;
input [7:0] bht_update_p1_sel_addr;
input [1:0] bht_update_p1_sel_data;
input [1:0] bht_update_p1_dir_data;
input [7:0] bht_dir_rd_addr;
input [7:0] bht_sel_rd_addr;
output [1:0] bht_taken_rdata;
output [1:0] bht_ntaken_rdata;
output [1:0] bht_sel_rdata;


generate
    if (BTB_SIZE != 0) begin:gen_bht_yes
        reg [1:0] s0[0:255];
        reg [1:0] s1[0:255];
        reg [1:0] s2[0:255];
        wire [7:0] s3;
        wire [7:0] s4;
        wire [7:0] s5;
        wire [7:0] s6;
        wire [255:0] s7;
        wire [255:0] s8;
        wire [255:0] s9;
        wire [255:0] s10;
        wire [255:0] s11;
        wire [255:0] s12;
        assign s3[7:0] = bht_update_p0_dir_addr[7:0];
        assign s4[7:0] = bht_update_p1_dir_addr[7:0];
        assign s5[7:0] = bht_update_p0_sel_addr[7:0];
        assign s6[7:0] = bht_update_p1_sel_addr[7:0];
        assign s7[0] = ((s3 == 8'd0) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[0] = ((s4 == 8'd0) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[0] = ((s3 == 8'd0) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[0] = ((s4 == 8'd0) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[0] = ((s5 == 8'd0) & bht_update_p0);
        assign s12[0] = ((s6 == 8'd0) & bht_update_p1);
        assign s7[1] = ((s3 == 8'd1) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[1] = ((s4 == 8'd1) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[1] = ((s3 == 8'd1) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[1] = ((s4 == 8'd1) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[1] = ((s5 == 8'd1) & bht_update_p0);
        assign s12[1] = ((s6 == 8'd1) & bht_update_p1);
        assign s7[2] = ((s3 == 8'd2) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[2] = ((s4 == 8'd2) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[2] = ((s3 == 8'd2) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[2] = ((s4 == 8'd2) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[2] = ((s5 == 8'd2) & bht_update_p0);
        assign s12[2] = ((s6 == 8'd2) & bht_update_p1);
        assign s7[3] = ((s3 == 8'd3) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[3] = ((s4 == 8'd3) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[3] = ((s3 == 8'd3) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[3] = ((s4 == 8'd3) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[3] = ((s5 == 8'd3) & bht_update_p0);
        assign s12[3] = ((s6 == 8'd3) & bht_update_p1);
        assign s7[4] = ((s3 == 8'd4) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[4] = ((s4 == 8'd4) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[4] = ((s3 == 8'd4) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[4] = ((s4 == 8'd4) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[4] = ((s5 == 8'd4) & bht_update_p0);
        assign s12[4] = ((s6 == 8'd4) & bht_update_p1);
        assign s7[5] = ((s3 == 8'd5) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[5] = ((s4 == 8'd5) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[5] = ((s3 == 8'd5) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[5] = ((s4 == 8'd5) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[5] = ((s5 == 8'd5) & bht_update_p0);
        assign s12[5] = ((s6 == 8'd5) & bht_update_p1);
        assign s7[6] = ((s3 == 8'd6) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[6] = ((s4 == 8'd6) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[6] = ((s3 == 8'd6) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[6] = ((s4 == 8'd6) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[6] = ((s5 == 8'd6) & bht_update_p0);
        assign s12[6] = ((s6 == 8'd6) & bht_update_p1);
        assign s7[7] = ((s3 == 8'd7) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[7] = ((s4 == 8'd7) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[7] = ((s3 == 8'd7) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[7] = ((s4 == 8'd7) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[7] = ((s5 == 8'd7) & bht_update_p0);
        assign s12[7] = ((s6 == 8'd7) & bht_update_p1);
        assign s7[8] = ((s3 == 8'd8) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[8] = ((s4 == 8'd8) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[8] = ((s3 == 8'd8) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[8] = ((s4 == 8'd8) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[8] = ((s5 == 8'd8) & bht_update_p0);
        assign s12[8] = ((s6 == 8'd8) & bht_update_p1);
        assign s7[9] = ((s3 == 8'd9) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[9] = ((s4 == 8'd9) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[9] = ((s3 == 8'd9) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[9] = ((s4 == 8'd9) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[9] = ((s5 == 8'd9) & bht_update_p0);
        assign s12[9] = ((s6 == 8'd9) & bht_update_p1);
        assign s7[10] = ((s3 == 8'd10) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[10] = ((s4 == 8'd10) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[10] = ((s3 == 8'd10) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[10] = ((s4 == 8'd10) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[10] = ((s5 == 8'd10) & bht_update_p0);
        assign s12[10] = ((s6 == 8'd10) & bht_update_p1);
        assign s7[11] = ((s3 == 8'd11) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[11] = ((s4 == 8'd11) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[11] = ((s3 == 8'd11) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[11] = ((s4 == 8'd11) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[11] = ((s5 == 8'd11) & bht_update_p0);
        assign s12[11] = ((s6 == 8'd11) & bht_update_p1);
        assign s7[12] = ((s3 == 8'd12) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[12] = ((s4 == 8'd12) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[12] = ((s3 == 8'd12) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[12] = ((s4 == 8'd12) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[12] = ((s5 == 8'd12) & bht_update_p0);
        assign s12[12] = ((s6 == 8'd12) & bht_update_p1);
        assign s7[13] = ((s3 == 8'd13) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[13] = ((s4 == 8'd13) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[13] = ((s3 == 8'd13) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[13] = ((s4 == 8'd13) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[13] = ((s5 == 8'd13) & bht_update_p0);
        assign s12[13] = ((s6 == 8'd13) & bht_update_p1);
        assign s7[14] = ((s3 == 8'd14) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[14] = ((s4 == 8'd14) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[14] = ((s3 == 8'd14) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[14] = ((s4 == 8'd14) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[14] = ((s5 == 8'd14) & bht_update_p0);
        assign s12[14] = ((s6 == 8'd14) & bht_update_p1);
        assign s7[15] = ((s3 == 8'd15) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[15] = ((s4 == 8'd15) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[15] = ((s3 == 8'd15) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[15] = ((s4 == 8'd15) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[15] = ((s5 == 8'd15) & bht_update_p0);
        assign s12[15] = ((s6 == 8'd15) & bht_update_p1);
        assign s7[16] = ((s3 == 8'd16) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[16] = ((s4 == 8'd16) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[16] = ((s3 == 8'd16) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[16] = ((s4 == 8'd16) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[16] = ((s5 == 8'd16) & bht_update_p0);
        assign s12[16] = ((s6 == 8'd16) & bht_update_p1);
        assign s7[17] = ((s3 == 8'd17) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[17] = ((s4 == 8'd17) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[17] = ((s3 == 8'd17) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[17] = ((s4 == 8'd17) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[17] = ((s5 == 8'd17) & bht_update_p0);
        assign s12[17] = ((s6 == 8'd17) & bht_update_p1);
        assign s7[18] = ((s3 == 8'd18) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[18] = ((s4 == 8'd18) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[18] = ((s3 == 8'd18) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[18] = ((s4 == 8'd18) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[18] = ((s5 == 8'd18) & bht_update_p0);
        assign s12[18] = ((s6 == 8'd18) & bht_update_p1);
        assign s7[19] = ((s3 == 8'd19) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[19] = ((s4 == 8'd19) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[19] = ((s3 == 8'd19) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[19] = ((s4 == 8'd19) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[19] = ((s5 == 8'd19) & bht_update_p0);
        assign s12[19] = ((s6 == 8'd19) & bht_update_p1);
        assign s7[20] = ((s3 == 8'd20) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[20] = ((s4 == 8'd20) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[20] = ((s3 == 8'd20) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[20] = ((s4 == 8'd20) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[20] = ((s5 == 8'd20) & bht_update_p0);
        assign s12[20] = ((s6 == 8'd20) & bht_update_p1);
        assign s7[21] = ((s3 == 8'd21) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[21] = ((s4 == 8'd21) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[21] = ((s3 == 8'd21) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[21] = ((s4 == 8'd21) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[21] = ((s5 == 8'd21) & bht_update_p0);
        assign s12[21] = ((s6 == 8'd21) & bht_update_p1);
        assign s7[22] = ((s3 == 8'd22) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[22] = ((s4 == 8'd22) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[22] = ((s3 == 8'd22) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[22] = ((s4 == 8'd22) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[22] = ((s5 == 8'd22) & bht_update_p0);
        assign s12[22] = ((s6 == 8'd22) & bht_update_p1);
        assign s7[23] = ((s3 == 8'd23) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[23] = ((s4 == 8'd23) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[23] = ((s3 == 8'd23) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[23] = ((s4 == 8'd23) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[23] = ((s5 == 8'd23) & bht_update_p0);
        assign s12[23] = ((s6 == 8'd23) & bht_update_p1);
        assign s7[24] = ((s3 == 8'd24) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[24] = ((s4 == 8'd24) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[24] = ((s3 == 8'd24) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[24] = ((s4 == 8'd24) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[24] = ((s5 == 8'd24) & bht_update_p0);
        assign s12[24] = ((s6 == 8'd24) & bht_update_p1);
        assign s7[25] = ((s3 == 8'd25) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[25] = ((s4 == 8'd25) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[25] = ((s3 == 8'd25) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[25] = ((s4 == 8'd25) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[25] = ((s5 == 8'd25) & bht_update_p0);
        assign s12[25] = ((s6 == 8'd25) & bht_update_p1);
        assign s7[26] = ((s3 == 8'd26) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[26] = ((s4 == 8'd26) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[26] = ((s3 == 8'd26) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[26] = ((s4 == 8'd26) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[26] = ((s5 == 8'd26) & bht_update_p0);
        assign s12[26] = ((s6 == 8'd26) & bht_update_p1);
        assign s7[27] = ((s3 == 8'd27) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[27] = ((s4 == 8'd27) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[27] = ((s3 == 8'd27) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[27] = ((s4 == 8'd27) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[27] = ((s5 == 8'd27) & bht_update_p0);
        assign s12[27] = ((s6 == 8'd27) & bht_update_p1);
        assign s7[28] = ((s3 == 8'd28) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[28] = ((s4 == 8'd28) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[28] = ((s3 == 8'd28) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[28] = ((s4 == 8'd28) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[28] = ((s5 == 8'd28) & bht_update_p0);
        assign s12[28] = ((s6 == 8'd28) & bht_update_p1);
        assign s7[29] = ((s3 == 8'd29) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[29] = ((s4 == 8'd29) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[29] = ((s3 == 8'd29) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[29] = ((s4 == 8'd29) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[29] = ((s5 == 8'd29) & bht_update_p0);
        assign s12[29] = ((s6 == 8'd29) & bht_update_p1);
        assign s7[30] = ((s3 == 8'd30) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[30] = ((s4 == 8'd30) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[30] = ((s3 == 8'd30) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[30] = ((s4 == 8'd30) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[30] = ((s5 == 8'd30) & bht_update_p0);
        assign s12[30] = ((s6 == 8'd30) & bht_update_p1);
        assign s7[31] = ((s3 == 8'd31) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[31] = ((s4 == 8'd31) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[31] = ((s3 == 8'd31) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[31] = ((s4 == 8'd31) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[31] = ((s5 == 8'd31) & bht_update_p0);
        assign s12[31] = ((s6 == 8'd31) & bht_update_p1);
        assign s7[32] = ((s3 == 8'd32) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[32] = ((s4 == 8'd32) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[32] = ((s3 == 8'd32) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[32] = ((s4 == 8'd32) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[32] = ((s5 == 8'd32) & bht_update_p0);
        assign s12[32] = ((s6 == 8'd32) & bht_update_p1);
        assign s7[33] = ((s3 == 8'd33) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[33] = ((s4 == 8'd33) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[33] = ((s3 == 8'd33) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[33] = ((s4 == 8'd33) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[33] = ((s5 == 8'd33) & bht_update_p0);
        assign s12[33] = ((s6 == 8'd33) & bht_update_p1);
        assign s7[34] = ((s3 == 8'd34) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[34] = ((s4 == 8'd34) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[34] = ((s3 == 8'd34) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[34] = ((s4 == 8'd34) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[34] = ((s5 == 8'd34) & bht_update_p0);
        assign s12[34] = ((s6 == 8'd34) & bht_update_p1);
        assign s7[35] = ((s3 == 8'd35) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[35] = ((s4 == 8'd35) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[35] = ((s3 == 8'd35) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[35] = ((s4 == 8'd35) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[35] = ((s5 == 8'd35) & bht_update_p0);
        assign s12[35] = ((s6 == 8'd35) & bht_update_p1);
        assign s7[36] = ((s3 == 8'd36) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[36] = ((s4 == 8'd36) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[36] = ((s3 == 8'd36) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[36] = ((s4 == 8'd36) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[36] = ((s5 == 8'd36) & bht_update_p0);
        assign s12[36] = ((s6 == 8'd36) & bht_update_p1);
        assign s7[37] = ((s3 == 8'd37) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[37] = ((s4 == 8'd37) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[37] = ((s3 == 8'd37) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[37] = ((s4 == 8'd37) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[37] = ((s5 == 8'd37) & bht_update_p0);
        assign s12[37] = ((s6 == 8'd37) & bht_update_p1);
        assign s7[38] = ((s3 == 8'd38) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[38] = ((s4 == 8'd38) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[38] = ((s3 == 8'd38) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[38] = ((s4 == 8'd38) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[38] = ((s5 == 8'd38) & bht_update_p0);
        assign s12[38] = ((s6 == 8'd38) & bht_update_p1);
        assign s7[39] = ((s3 == 8'd39) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[39] = ((s4 == 8'd39) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[39] = ((s3 == 8'd39) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[39] = ((s4 == 8'd39) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[39] = ((s5 == 8'd39) & bht_update_p0);
        assign s12[39] = ((s6 == 8'd39) & bht_update_p1);
        assign s7[40] = ((s3 == 8'd40) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[40] = ((s4 == 8'd40) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[40] = ((s3 == 8'd40) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[40] = ((s4 == 8'd40) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[40] = ((s5 == 8'd40) & bht_update_p0);
        assign s12[40] = ((s6 == 8'd40) & bht_update_p1);
        assign s7[41] = ((s3 == 8'd41) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[41] = ((s4 == 8'd41) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[41] = ((s3 == 8'd41) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[41] = ((s4 == 8'd41) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[41] = ((s5 == 8'd41) & bht_update_p0);
        assign s12[41] = ((s6 == 8'd41) & bht_update_p1);
        assign s7[42] = ((s3 == 8'd42) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[42] = ((s4 == 8'd42) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[42] = ((s3 == 8'd42) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[42] = ((s4 == 8'd42) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[42] = ((s5 == 8'd42) & bht_update_p0);
        assign s12[42] = ((s6 == 8'd42) & bht_update_p1);
        assign s7[43] = ((s3 == 8'd43) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[43] = ((s4 == 8'd43) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[43] = ((s3 == 8'd43) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[43] = ((s4 == 8'd43) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[43] = ((s5 == 8'd43) & bht_update_p0);
        assign s12[43] = ((s6 == 8'd43) & bht_update_p1);
        assign s7[44] = ((s3 == 8'd44) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[44] = ((s4 == 8'd44) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[44] = ((s3 == 8'd44) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[44] = ((s4 == 8'd44) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[44] = ((s5 == 8'd44) & bht_update_p0);
        assign s12[44] = ((s6 == 8'd44) & bht_update_p1);
        assign s7[45] = ((s3 == 8'd45) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[45] = ((s4 == 8'd45) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[45] = ((s3 == 8'd45) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[45] = ((s4 == 8'd45) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[45] = ((s5 == 8'd45) & bht_update_p0);
        assign s12[45] = ((s6 == 8'd45) & bht_update_p1);
        assign s7[46] = ((s3 == 8'd46) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[46] = ((s4 == 8'd46) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[46] = ((s3 == 8'd46) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[46] = ((s4 == 8'd46) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[46] = ((s5 == 8'd46) & bht_update_p0);
        assign s12[46] = ((s6 == 8'd46) & bht_update_p1);
        assign s7[47] = ((s3 == 8'd47) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[47] = ((s4 == 8'd47) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[47] = ((s3 == 8'd47) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[47] = ((s4 == 8'd47) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[47] = ((s5 == 8'd47) & bht_update_p0);
        assign s12[47] = ((s6 == 8'd47) & bht_update_p1);
        assign s7[48] = ((s3 == 8'd48) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[48] = ((s4 == 8'd48) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[48] = ((s3 == 8'd48) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[48] = ((s4 == 8'd48) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[48] = ((s5 == 8'd48) & bht_update_p0);
        assign s12[48] = ((s6 == 8'd48) & bht_update_p1);
        assign s7[49] = ((s3 == 8'd49) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[49] = ((s4 == 8'd49) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[49] = ((s3 == 8'd49) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[49] = ((s4 == 8'd49) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[49] = ((s5 == 8'd49) & bht_update_p0);
        assign s12[49] = ((s6 == 8'd49) & bht_update_p1);
        assign s7[50] = ((s3 == 8'd50) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[50] = ((s4 == 8'd50) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[50] = ((s3 == 8'd50) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[50] = ((s4 == 8'd50) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[50] = ((s5 == 8'd50) & bht_update_p0);
        assign s12[50] = ((s6 == 8'd50) & bht_update_p1);
        assign s7[51] = ((s3 == 8'd51) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[51] = ((s4 == 8'd51) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[51] = ((s3 == 8'd51) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[51] = ((s4 == 8'd51) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[51] = ((s5 == 8'd51) & bht_update_p0);
        assign s12[51] = ((s6 == 8'd51) & bht_update_p1);
        assign s7[52] = ((s3 == 8'd52) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[52] = ((s4 == 8'd52) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[52] = ((s3 == 8'd52) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[52] = ((s4 == 8'd52) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[52] = ((s5 == 8'd52) & bht_update_p0);
        assign s12[52] = ((s6 == 8'd52) & bht_update_p1);
        assign s7[53] = ((s3 == 8'd53) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[53] = ((s4 == 8'd53) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[53] = ((s3 == 8'd53) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[53] = ((s4 == 8'd53) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[53] = ((s5 == 8'd53) & bht_update_p0);
        assign s12[53] = ((s6 == 8'd53) & bht_update_p1);
        assign s7[54] = ((s3 == 8'd54) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[54] = ((s4 == 8'd54) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[54] = ((s3 == 8'd54) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[54] = ((s4 == 8'd54) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[54] = ((s5 == 8'd54) & bht_update_p0);
        assign s12[54] = ((s6 == 8'd54) & bht_update_p1);
        assign s7[55] = ((s3 == 8'd55) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[55] = ((s4 == 8'd55) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[55] = ((s3 == 8'd55) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[55] = ((s4 == 8'd55) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[55] = ((s5 == 8'd55) & bht_update_p0);
        assign s12[55] = ((s6 == 8'd55) & bht_update_p1);
        assign s7[56] = ((s3 == 8'd56) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[56] = ((s4 == 8'd56) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[56] = ((s3 == 8'd56) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[56] = ((s4 == 8'd56) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[56] = ((s5 == 8'd56) & bht_update_p0);
        assign s12[56] = ((s6 == 8'd56) & bht_update_p1);
        assign s7[57] = ((s3 == 8'd57) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[57] = ((s4 == 8'd57) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[57] = ((s3 == 8'd57) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[57] = ((s4 == 8'd57) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[57] = ((s5 == 8'd57) & bht_update_p0);
        assign s12[57] = ((s6 == 8'd57) & bht_update_p1);
        assign s7[58] = ((s3 == 8'd58) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[58] = ((s4 == 8'd58) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[58] = ((s3 == 8'd58) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[58] = ((s4 == 8'd58) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[58] = ((s5 == 8'd58) & bht_update_p0);
        assign s12[58] = ((s6 == 8'd58) & bht_update_p1);
        assign s7[59] = ((s3 == 8'd59) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[59] = ((s4 == 8'd59) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[59] = ((s3 == 8'd59) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[59] = ((s4 == 8'd59) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[59] = ((s5 == 8'd59) & bht_update_p0);
        assign s12[59] = ((s6 == 8'd59) & bht_update_p1);
        assign s7[60] = ((s3 == 8'd60) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[60] = ((s4 == 8'd60) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[60] = ((s3 == 8'd60) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[60] = ((s4 == 8'd60) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[60] = ((s5 == 8'd60) & bht_update_p0);
        assign s12[60] = ((s6 == 8'd60) & bht_update_p1);
        assign s7[61] = ((s3 == 8'd61) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[61] = ((s4 == 8'd61) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[61] = ((s3 == 8'd61) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[61] = ((s4 == 8'd61) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[61] = ((s5 == 8'd61) & bht_update_p0);
        assign s12[61] = ((s6 == 8'd61) & bht_update_p1);
        assign s7[62] = ((s3 == 8'd62) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[62] = ((s4 == 8'd62) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[62] = ((s3 == 8'd62) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[62] = ((s4 == 8'd62) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[62] = ((s5 == 8'd62) & bht_update_p0);
        assign s12[62] = ((s6 == 8'd62) & bht_update_p1);
        assign s7[63] = ((s3 == 8'd63) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[63] = ((s4 == 8'd63) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[63] = ((s3 == 8'd63) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[63] = ((s4 == 8'd63) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[63] = ((s5 == 8'd63) & bht_update_p0);
        assign s12[63] = ((s6 == 8'd63) & bht_update_p1);
        assign s7[64] = ((s3 == 8'd64) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[64] = ((s4 == 8'd64) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[64] = ((s3 == 8'd64) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[64] = ((s4 == 8'd64) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[64] = ((s5 == 8'd64) & bht_update_p0);
        assign s12[64] = ((s6 == 8'd64) & bht_update_p1);
        assign s7[65] = ((s3 == 8'd65) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[65] = ((s4 == 8'd65) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[65] = ((s3 == 8'd65) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[65] = ((s4 == 8'd65) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[65] = ((s5 == 8'd65) & bht_update_p0);
        assign s12[65] = ((s6 == 8'd65) & bht_update_p1);
        assign s7[66] = ((s3 == 8'd66) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[66] = ((s4 == 8'd66) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[66] = ((s3 == 8'd66) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[66] = ((s4 == 8'd66) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[66] = ((s5 == 8'd66) & bht_update_p0);
        assign s12[66] = ((s6 == 8'd66) & bht_update_p1);
        assign s7[67] = ((s3 == 8'd67) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[67] = ((s4 == 8'd67) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[67] = ((s3 == 8'd67) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[67] = ((s4 == 8'd67) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[67] = ((s5 == 8'd67) & bht_update_p0);
        assign s12[67] = ((s6 == 8'd67) & bht_update_p1);
        assign s7[68] = ((s3 == 8'd68) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[68] = ((s4 == 8'd68) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[68] = ((s3 == 8'd68) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[68] = ((s4 == 8'd68) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[68] = ((s5 == 8'd68) & bht_update_p0);
        assign s12[68] = ((s6 == 8'd68) & bht_update_p1);
        assign s7[69] = ((s3 == 8'd69) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[69] = ((s4 == 8'd69) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[69] = ((s3 == 8'd69) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[69] = ((s4 == 8'd69) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[69] = ((s5 == 8'd69) & bht_update_p0);
        assign s12[69] = ((s6 == 8'd69) & bht_update_p1);
        assign s7[70] = ((s3 == 8'd70) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[70] = ((s4 == 8'd70) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[70] = ((s3 == 8'd70) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[70] = ((s4 == 8'd70) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[70] = ((s5 == 8'd70) & bht_update_p0);
        assign s12[70] = ((s6 == 8'd70) & bht_update_p1);
        assign s7[71] = ((s3 == 8'd71) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[71] = ((s4 == 8'd71) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[71] = ((s3 == 8'd71) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[71] = ((s4 == 8'd71) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[71] = ((s5 == 8'd71) & bht_update_p0);
        assign s12[71] = ((s6 == 8'd71) & bht_update_p1);
        assign s7[72] = ((s3 == 8'd72) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[72] = ((s4 == 8'd72) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[72] = ((s3 == 8'd72) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[72] = ((s4 == 8'd72) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[72] = ((s5 == 8'd72) & bht_update_p0);
        assign s12[72] = ((s6 == 8'd72) & bht_update_p1);
        assign s7[73] = ((s3 == 8'd73) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[73] = ((s4 == 8'd73) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[73] = ((s3 == 8'd73) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[73] = ((s4 == 8'd73) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[73] = ((s5 == 8'd73) & bht_update_p0);
        assign s12[73] = ((s6 == 8'd73) & bht_update_p1);
        assign s7[74] = ((s3 == 8'd74) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[74] = ((s4 == 8'd74) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[74] = ((s3 == 8'd74) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[74] = ((s4 == 8'd74) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[74] = ((s5 == 8'd74) & bht_update_p0);
        assign s12[74] = ((s6 == 8'd74) & bht_update_p1);
        assign s7[75] = ((s3 == 8'd75) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[75] = ((s4 == 8'd75) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[75] = ((s3 == 8'd75) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[75] = ((s4 == 8'd75) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[75] = ((s5 == 8'd75) & bht_update_p0);
        assign s12[75] = ((s6 == 8'd75) & bht_update_p1);
        assign s7[76] = ((s3 == 8'd76) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[76] = ((s4 == 8'd76) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[76] = ((s3 == 8'd76) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[76] = ((s4 == 8'd76) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[76] = ((s5 == 8'd76) & bht_update_p0);
        assign s12[76] = ((s6 == 8'd76) & bht_update_p1);
        assign s7[77] = ((s3 == 8'd77) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[77] = ((s4 == 8'd77) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[77] = ((s3 == 8'd77) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[77] = ((s4 == 8'd77) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[77] = ((s5 == 8'd77) & bht_update_p0);
        assign s12[77] = ((s6 == 8'd77) & bht_update_p1);
        assign s7[78] = ((s3 == 8'd78) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[78] = ((s4 == 8'd78) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[78] = ((s3 == 8'd78) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[78] = ((s4 == 8'd78) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[78] = ((s5 == 8'd78) & bht_update_p0);
        assign s12[78] = ((s6 == 8'd78) & bht_update_p1);
        assign s7[79] = ((s3 == 8'd79) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[79] = ((s4 == 8'd79) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[79] = ((s3 == 8'd79) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[79] = ((s4 == 8'd79) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[79] = ((s5 == 8'd79) & bht_update_p0);
        assign s12[79] = ((s6 == 8'd79) & bht_update_p1);
        assign s7[80] = ((s3 == 8'd80) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[80] = ((s4 == 8'd80) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[80] = ((s3 == 8'd80) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[80] = ((s4 == 8'd80) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[80] = ((s5 == 8'd80) & bht_update_p0);
        assign s12[80] = ((s6 == 8'd80) & bht_update_p1);
        assign s7[81] = ((s3 == 8'd81) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[81] = ((s4 == 8'd81) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[81] = ((s3 == 8'd81) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[81] = ((s4 == 8'd81) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[81] = ((s5 == 8'd81) & bht_update_p0);
        assign s12[81] = ((s6 == 8'd81) & bht_update_p1);
        assign s7[82] = ((s3 == 8'd82) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[82] = ((s4 == 8'd82) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[82] = ((s3 == 8'd82) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[82] = ((s4 == 8'd82) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[82] = ((s5 == 8'd82) & bht_update_p0);
        assign s12[82] = ((s6 == 8'd82) & bht_update_p1);
        assign s7[83] = ((s3 == 8'd83) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[83] = ((s4 == 8'd83) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[83] = ((s3 == 8'd83) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[83] = ((s4 == 8'd83) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[83] = ((s5 == 8'd83) & bht_update_p0);
        assign s12[83] = ((s6 == 8'd83) & bht_update_p1);
        assign s7[84] = ((s3 == 8'd84) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[84] = ((s4 == 8'd84) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[84] = ((s3 == 8'd84) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[84] = ((s4 == 8'd84) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[84] = ((s5 == 8'd84) & bht_update_p0);
        assign s12[84] = ((s6 == 8'd84) & bht_update_p1);
        assign s7[85] = ((s3 == 8'd85) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[85] = ((s4 == 8'd85) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[85] = ((s3 == 8'd85) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[85] = ((s4 == 8'd85) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[85] = ((s5 == 8'd85) & bht_update_p0);
        assign s12[85] = ((s6 == 8'd85) & bht_update_p1);
        assign s7[86] = ((s3 == 8'd86) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[86] = ((s4 == 8'd86) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[86] = ((s3 == 8'd86) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[86] = ((s4 == 8'd86) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[86] = ((s5 == 8'd86) & bht_update_p0);
        assign s12[86] = ((s6 == 8'd86) & bht_update_p1);
        assign s7[87] = ((s3 == 8'd87) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[87] = ((s4 == 8'd87) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[87] = ((s3 == 8'd87) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[87] = ((s4 == 8'd87) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[87] = ((s5 == 8'd87) & bht_update_p0);
        assign s12[87] = ((s6 == 8'd87) & bht_update_p1);
        assign s7[88] = ((s3 == 8'd88) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[88] = ((s4 == 8'd88) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[88] = ((s3 == 8'd88) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[88] = ((s4 == 8'd88) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[88] = ((s5 == 8'd88) & bht_update_p0);
        assign s12[88] = ((s6 == 8'd88) & bht_update_p1);
        assign s7[89] = ((s3 == 8'd89) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[89] = ((s4 == 8'd89) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[89] = ((s3 == 8'd89) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[89] = ((s4 == 8'd89) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[89] = ((s5 == 8'd89) & bht_update_p0);
        assign s12[89] = ((s6 == 8'd89) & bht_update_p1);
        assign s7[90] = ((s3 == 8'd90) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[90] = ((s4 == 8'd90) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[90] = ((s3 == 8'd90) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[90] = ((s4 == 8'd90) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[90] = ((s5 == 8'd90) & bht_update_p0);
        assign s12[90] = ((s6 == 8'd90) & bht_update_p1);
        assign s7[91] = ((s3 == 8'd91) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[91] = ((s4 == 8'd91) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[91] = ((s3 == 8'd91) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[91] = ((s4 == 8'd91) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[91] = ((s5 == 8'd91) & bht_update_p0);
        assign s12[91] = ((s6 == 8'd91) & bht_update_p1);
        assign s7[92] = ((s3 == 8'd92) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[92] = ((s4 == 8'd92) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[92] = ((s3 == 8'd92) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[92] = ((s4 == 8'd92) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[92] = ((s5 == 8'd92) & bht_update_p0);
        assign s12[92] = ((s6 == 8'd92) & bht_update_p1);
        assign s7[93] = ((s3 == 8'd93) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[93] = ((s4 == 8'd93) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[93] = ((s3 == 8'd93) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[93] = ((s4 == 8'd93) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[93] = ((s5 == 8'd93) & bht_update_p0);
        assign s12[93] = ((s6 == 8'd93) & bht_update_p1);
        assign s7[94] = ((s3 == 8'd94) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[94] = ((s4 == 8'd94) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[94] = ((s3 == 8'd94) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[94] = ((s4 == 8'd94) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[94] = ((s5 == 8'd94) & bht_update_p0);
        assign s12[94] = ((s6 == 8'd94) & bht_update_p1);
        assign s7[95] = ((s3 == 8'd95) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[95] = ((s4 == 8'd95) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[95] = ((s3 == 8'd95) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[95] = ((s4 == 8'd95) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[95] = ((s5 == 8'd95) & bht_update_p0);
        assign s12[95] = ((s6 == 8'd95) & bht_update_p1);
        assign s7[96] = ((s3 == 8'd96) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[96] = ((s4 == 8'd96) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[96] = ((s3 == 8'd96) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[96] = ((s4 == 8'd96) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[96] = ((s5 == 8'd96) & bht_update_p0);
        assign s12[96] = ((s6 == 8'd96) & bht_update_p1);
        assign s7[97] = ((s3 == 8'd97) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[97] = ((s4 == 8'd97) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[97] = ((s3 == 8'd97) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[97] = ((s4 == 8'd97) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[97] = ((s5 == 8'd97) & bht_update_p0);
        assign s12[97] = ((s6 == 8'd97) & bht_update_p1);
        assign s7[98] = ((s3 == 8'd98) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[98] = ((s4 == 8'd98) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[98] = ((s3 == 8'd98) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[98] = ((s4 == 8'd98) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[98] = ((s5 == 8'd98) & bht_update_p0);
        assign s12[98] = ((s6 == 8'd98) & bht_update_p1);
        assign s7[99] = ((s3 == 8'd99) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[99] = ((s4 == 8'd99) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[99] = ((s3 == 8'd99) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[99] = ((s4 == 8'd99) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[99] = ((s5 == 8'd99) & bht_update_p0);
        assign s12[99] = ((s6 == 8'd99) & bht_update_p1);
        assign s7[100] = ((s3 == 8'd100) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[100] = ((s4 == 8'd100) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[100] = ((s3 == 8'd100) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[100] = ((s4 == 8'd100) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[100] = ((s5 == 8'd100) & bht_update_p0);
        assign s12[100] = ((s6 == 8'd100) & bht_update_p1);
        assign s7[101] = ((s3 == 8'd101) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[101] = ((s4 == 8'd101) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[101] = ((s3 == 8'd101) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[101] = ((s4 == 8'd101) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[101] = ((s5 == 8'd101) & bht_update_p0);
        assign s12[101] = ((s6 == 8'd101) & bht_update_p1);
        assign s7[102] = ((s3 == 8'd102) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[102] = ((s4 == 8'd102) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[102] = ((s3 == 8'd102) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[102] = ((s4 == 8'd102) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[102] = ((s5 == 8'd102) & bht_update_p0);
        assign s12[102] = ((s6 == 8'd102) & bht_update_p1);
        assign s7[103] = ((s3 == 8'd103) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[103] = ((s4 == 8'd103) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[103] = ((s3 == 8'd103) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[103] = ((s4 == 8'd103) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[103] = ((s5 == 8'd103) & bht_update_p0);
        assign s12[103] = ((s6 == 8'd103) & bht_update_p1);
        assign s7[104] = ((s3 == 8'd104) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[104] = ((s4 == 8'd104) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[104] = ((s3 == 8'd104) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[104] = ((s4 == 8'd104) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[104] = ((s5 == 8'd104) & bht_update_p0);
        assign s12[104] = ((s6 == 8'd104) & bht_update_p1);
        assign s7[105] = ((s3 == 8'd105) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[105] = ((s4 == 8'd105) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[105] = ((s3 == 8'd105) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[105] = ((s4 == 8'd105) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[105] = ((s5 == 8'd105) & bht_update_p0);
        assign s12[105] = ((s6 == 8'd105) & bht_update_p1);
        assign s7[106] = ((s3 == 8'd106) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[106] = ((s4 == 8'd106) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[106] = ((s3 == 8'd106) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[106] = ((s4 == 8'd106) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[106] = ((s5 == 8'd106) & bht_update_p0);
        assign s12[106] = ((s6 == 8'd106) & bht_update_p1);
        assign s7[107] = ((s3 == 8'd107) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[107] = ((s4 == 8'd107) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[107] = ((s3 == 8'd107) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[107] = ((s4 == 8'd107) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[107] = ((s5 == 8'd107) & bht_update_p0);
        assign s12[107] = ((s6 == 8'd107) & bht_update_p1);
        assign s7[108] = ((s3 == 8'd108) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[108] = ((s4 == 8'd108) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[108] = ((s3 == 8'd108) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[108] = ((s4 == 8'd108) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[108] = ((s5 == 8'd108) & bht_update_p0);
        assign s12[108] = ((s6 == 8'd108) & bht_update_p1);
        assign s7[109] = ((s3 == 8'd109) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[109] = ((s4 == 8'd109) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[109] = ((s3 == 8'd109) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[109] = ((s4 == 8'd109) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[109] = ((s5 == 8'd109) & bht_update_p0);
        assign s12[109] = ((s6 == 8'd109) & bht_update_p1);
        assign s7[110] = ((s3 == 8'd110) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[110] = ((s4 == 8'd110) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[110] = ((s3 == 8'd110) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[110] = ((s4 == 8'd110) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[110] = ((s5 == 8'd110) & bht_update_p0);
        assign s12[110] = ((s6 == 8'd110) & bht_update_p1);
        assign s7[111] = ((s3 == 8'd111) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[111] = ((s4 == 8'd111) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[111] = ((s3 == 8'd111) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[111] = ((s4 == 8'd111) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[111] = ((s5 == 8'd111) & bht_update_p0);
        assign s12[111] = ((s6 == 8'd111) & bht_update_p1);
        assign s7[112] = ((s3 == 8'd112) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[112] = ((s4 == 8'd112) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[112] = ((s3 == 8'd112) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[112] = ((s4 == 8'd112) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[112] = ((s5 == 8'd112) & bht_update_p0);
        assign s12[112] = ((s6 == 8'd112) & bht_update_p1);
        assign s7[113] = ((s3 == 8'd113) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[113] = ((s4 == 8'd113) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[113] = ((s3 == 8'd113) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[113] = ((s4 == 8'd113) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[113] = ((s5 == 8'd113) & bht_update_p0);
        assign s12[113] = ((s6 == 8'd113) & bht_update_p1);
        assign s7[114] = ((s3 == 8'd114) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[114] = ((s4 == 8'd114) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[114] = ((s3 == 8'd114) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[114] = ((s4 == 8'd114) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[114] = ((s5 == 8'd114) & bht_update_p0);
        assign s12[114] = ((s6 == 8'd114) & bht_update_p1);
        assign s7[115] = ((s3 == 8'd115) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[115] = ((s4 == 8'd115) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[115] = ((s3 == 8'd115) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[115] = ((s4 == 8'd115) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[115] = ((s5 == 8'd115) & bht_update_p0);
        assign s12[115] = ((s6 == 8'd115) & bht_update_p1);
        assign s7[116] = ((s3 == 8'd116) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[116] = ((s4 == 8'd116) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[116] = ((s3 == 8'd116) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[116] = ((s4 == 8'd116) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[116] = ((s5 == 8'd116) & bht_update_p0);
        assign s12[116] = ((s6 == 8'd116) & bht_update_p1);
        assign s7[117] = ((s3 == 8'd117) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[117] = ((s4 == 8'd117) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[117] = ((s3 == 8'd117) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[117] = ((s4 == 8'd117) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[117] = ((s5 == 8'd117) & bht_update_p0);
        assign s12[117] = ((s6 == 8'd117) & bht_update_p1);
        assign s7[118] = ((s3 == 8'd118) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[118] = ((s4 == 8'd118) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[118] = ((s3 == 8'd118) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[118] = ((s4 == 8'd118) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[118] = ((s5 == 8'd118) & bht_update_p0);
        assign s12[118] = ((s6 == 8'd118) & bht_update_p1);
        assign s7[119] = ((s3 == 8'd119) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[119] = ((s4 == 8'd119) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[119] = ((s3 == 8'd119) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[119] = ((s4 == 8'd119) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[119] = ((s5 == 8'd119) & bht_update_p0);
        assign s12[119] = ((s6 == 8'd119) & bht_update_p1);
        assign s7[120] = ((s3 == 8'd120) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[120] = ((s4 == 8'd120) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[120] = ((s3 == 8'd120) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[120] = ((s4 == 8'd120) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[120] = ((s5 == 8'd120) & bht_update_p0);
        assign s12[120] = ((s6 == 8'd120) & bht_update_p1);
        assign s7[121] = ((s3 == 8'd121) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[121] = ((s4 == 8'd121) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[121] = ((s3 == 8'd121) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[121] = ((s4 == 8'd121) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[121] = ((s5 == 8'd121) & bht_update_p0);
        assign s12[121] = ((s6 == 8'd121) & bht_update_p1);
        assign s7[122] = ((s3 == 8'd122) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[122] = ((s4 == 8'd122) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[122] = ((s3 == 8'd122) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[122] = ((s4 == 8'd122) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[122] = ((s5 == 8'd122) & bht_update_p0);
        assign s12[122] = ((s6 == 8'd122) & bht_update_p1);
        assign s7[123] = ((s3 == 8'd123) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[123] = ((s4 == 8'd123) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[123] = ((s3 == 8'd123) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[123] = ((s4 == 8'd123) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[123] = ((s5 == 8'd123) & bht_update_p0);
        assign s12[123] = ((s6 == 8'd123) & bht_update_p1);
        assign s7[124] = ((s3 == 8'd124) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[124] = ((s4 == 8'd124) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[124] = ((s3 == 8'd124) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[124] = ((s4 == 8'd124) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[124] = ((s5 == 8'd124) & bht_update_p0);
        assign s12[124] = ((s6 == 8'd124) & bht_update_p1);
        assign s7[125] = ((s3 == 8'd125) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[125] = ((s4 == 8'd125) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[125] = ((s3 == 8'd125) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[125] = ((s4 == 8'd125) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[125] = ((s5 == 8'd125) & bht_update_p0);
        assign s12[125] = ((s6 == 8'd125) & bht_update_p1);
        assign s7[126] = ((s3 == 8'd126) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[126] = ((s4 == 8'd126) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[126] = ((s3 == 8'd126) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[126] = ((s4 == 8'd126) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[126] = ((s5 == 8'd126) & bht_update_p0);
        assign s12[126] = ((s6 == 8'd126) & bht_update_p1);
        assign s7[127] = ((s3 == 8'd127) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[127] = ((s4 == 8'd127) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[127] = ((s3 == 8'd127) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[127] = ((s4 == 8'd127) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[127] = ((s5 == 8'd127) & bht_update_p0);
        assign s12[127] = ((s6 == 8'd127) & bht_update_p1);
        assign s7[128] = ((s3 == 8'd128) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[128] = ((s4 == 8'd128) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[128] = ((s3 == 8'd128) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[128] = ((s4 == 8'd128) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[128] = ((s5 == 8'd128) & bht_update_p0);
        assign s12[128] = ((s6 == 8'd128) & bht_update_p1);
        assign s7[129] = ((s3 == 8'd129) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[129] = ((s4 == 8'd129) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[129] = ((s3 == 8'd129) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[129] = ((s4 == 8'd129) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[129] = ((s5 == 8'd129) & bht_update_p0);
        assign s12[129] = ((s6 == 8'd129) & bht_update_p1);
        assign s7[130] = ((s3 == 8'd130) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[130] = ((s4 == 8'd130) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[130] = ((s3 == 8'd130) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[130] = ((s4 == 8'd130) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[130] = ((s5 == 8'd130) & bht_update_p0);
        assign s12[130] = ((s6 == 8'd130) & bht_update_p1);
        assign s7[131] = ((s3 == 8'd131) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[131] = ((s4 == 8'd131) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[131] = ((s3 == 8'd131) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[131] = ((s4 == 8'd131) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[131] = ((s5 == 8'd131) & bht_update_p0);
        assign s12[131] = ((s6 == 8'd131) & bht_update_p1);
        assign s7[132] = ((s3 == 8'd132) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[132] = ((s4 == 8'd132) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[132] = ((s3 == 8'd132) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[132] = ((s4 == 8'd132) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[132] = ((s5 == 8'd132) & bht_update_p0);
        assign s12[132] = ((s6 == 8'd132) & bht_update_p1);
        assign s7[133] = ((s3 == 8'd133) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[133] = ((s4 == 8'd133) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[133] = ((s3 == 8'd133) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[133] = ((s4 == 8'd133) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[133] = ((s5 == 8'd133) & bht_update_p0);
        assign s12[133] = ((s6 == 8'd133) & bht_update_p1);
        assign s7[134] = ((s3 == 8'd134) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[134] = ((s4 == 8'd134) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[134] = ((s3 == 8'd134) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[134] = ((s4 == 8'd134) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[134] = ((s5 == 8'd134) & bht_update_p0);
        assign s12[134] = ((s6 == 8'd134) & bht_update_p1);
        assign s7[135] = ((s3 == 8'd135) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[135] = ((s4 == 8'd135) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[135] = ((s3 == 8'd135) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[135] = ((s4 == 8'd135) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[135] = ((s5 == 8'd135) & bht_update_p0);
        assign s12[135] = ((s6 == 8'd135) & bht_update_p1);
        assign s7[136] = ((s3 == 8'd136) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[136] = ((s4 == 8'd136) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[136] = ((s3 == 8'd136) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[136] = ((s4 == 8'd136) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[136] = ((s5 == 8'd136) & bht_update_p0);
        assign s12[136] = ((s6 == 8'd136) & bht_update_p1);
        assign s7[137] = ((s3 == 8'd137) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[137] = ((s4 == 8'd137) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[137] = ((s3 == 8'd137) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[137] = ((s4 == 8'd137) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[137] = ((s5 == 8'd137) & bht_update_p0);
        assign s12[137] = ((s6 == 8'd137) & bht_update_p1);
        assign s7[138] = ((s3 == 8'd138) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[138] = ((s4 == 8'd138) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[138] = ((s3 == 8'd138) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[138] = ((s4 == 8'd138) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[138] = ((s5 == 8'd138) & bht_update_p0);
        assign s12[138] = ((s6 == 8'd138) & bht_update_p1);
        assign s7[139] = ((s3 == 8'd139) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[139] = ((s4 == 8'd139) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[139] = ((s3 == 8'd139) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[139] = ((s4 == 8'd139) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[139] = ((s5 == 8'd139) & bht_update_p0);
        assign s12[139] = ((s6 == 8'd139) & bht_update_p1);
        assign s7[140] = ((s3 == 8'd140) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[140] = ((s4 == 8'd140) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[140] = ((s3 == 8'd140) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[140] = ((s4 == 8'd140) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[140] = ((s5 == 8'd140) & bht_update_p0);
        assign s12[140] = ((s6 == 8'd140) & bht_update_p1);
        assign s7[141] = ((s3 == 8'd141) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[141] = ((s4 == 8'd141) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[141] = ((s3 == 8'd141) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[141] = ((s4 == 8'd141) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[141] = ((s5 == 8'd141) & bht_update_p0);
        assign s12[141] = ((s6 == 8'd141) & bht_update_p1);
        assign s7[142] = ((s3 == 8'd142) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[142] = ((s4 == 8'd142) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[142] = ((s3 == 8'd142) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[142] = ((s4 == 8'd142) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[142] = ((s5 == 8'd142) & bht_update_p0);
        assign s12[142] = ((s6 == 8'd142) & bht_update_p1);
        assign s7[143] = ((s3 == 8'd143) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[143] = ((s4 == 8'd143) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[143] = ((s3 == 8'd143) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[143] = ((s4 == 8'd143) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[143] = ((s5 == 8'd143) & bht_update_p0);
        assign s12[143] = ((s6 == 8'd143) & bht_update_p1);
        assign s7[144] = ((s3 == 8'd144) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[144] = ((s4 == 8'd144) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[144] = ((s3 == 8'd144) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[144] = ((s4 == 8'd144) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[144] = ((s5 == 8'd144) & bht_update_p0);
        assign s12[144] = ((s6 == 8'd144) & bht_update_p1);
        assign s7[145] = ((s3 == 8'd145) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[145] = ((s4 == 8'd145) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[145] = ((s3 == 8'd145) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[145] = ((s4 == 8'd145) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[145] = ((s5 == 8'd145) & bht_update_p0);
        assign s12[145] = ((s6 == 8'd145) & bht_update_p1);
        assign s7[146] = ((s3 == 8'd146) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[146] = ((s4 == 8'd146) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[146] = ((s3 == 8'd146) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[146] = ((s4 == 8'd146) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[146] = ((s5 == 8'd146) & bht_update_p0);
        assign s12[146] = ((s6 == 8'd146) & bht_update_p1);
        assign s7[147] = ((s3 == 8'd147) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[147] = ((s4 == 8'd147) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[147] = ((s3 == 8'd147) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[147] = ((s4 == 8'd147) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[147] = ((s5 == 8'd147) & bht_update_p0);
        assign s12[147] = ((s6 == 8'd147) & bht_update_p1);
        assign s7[148] = ((s3 == 8'd148) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[148] = ((s4 == 8'd148) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[148] = ((s3 == 8'd148) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[148] = ((s4 == 8'd148) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[148] = ((s5 == 8'd148) & bht_update_p0);
        assign s12[148] = ((s6 == 8'd148) & bht_update_p1);
        assign s7[149] = ((s3 == 8'd149) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[149] = ((s4 == 8'd149) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[149] = ((s3 == 8'd149) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[149] = ((s4 == 8'd149) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[149] = ((s5 == 8'd149) & bht_update_p0);
        assign s12[149] = ((s6 == 8'd149) & bht_update_p1);
        assign s7[150] = ((s3 == 8'd150) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[150] = ((s4 == 8'd150) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[150] = ((s3 == 8'd150) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[150] = ((s4 == 8'd150) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[150] = ((s5 == 8'd150) & bht_update_p0);
        assign s12[150] = ((s6 == 8'd150) & bht_update_p1);
        assign s7[151] = ((s3 == 8'd151) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[151] = ((s4 == 8'd151) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[151] = ((s3 == 8'd151) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[151] = ((s4 == 8'd151) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[151] = ((s5 == 8'd151) & bht_update_p0);
        assign s12[151] = ((s6 == 8'd151) & bht_update_p1);
        assign s7[152] = ((s3 == 8'd152) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[152] = ((s4 == 8'd152) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[152] = ((s3 == 8'd152) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[152] = ((s4 == 8'd152) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[152] = ((s5 == 8'd152) & bht_update_p0);
        assign s12[152] = ((s6 == 8'd152) & bht_update_p1);
        assign s7[153] = ((s3 == 8'd153) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[153] = ((s4 == 8'd153) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[153] = ((s3 == 8'd153) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[153] = ((s4 == 8'd153) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[153] = ((s5 == 8'd153) & bht_update_p0);
        assign s12[153] = ((s6 == 8'd153) & bht_update_p1);
        assign s7[154] = ((s3 == 8'd154) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[154] = ((s4 == 8'd154) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[154] = ((s3 == 8'd154) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[154] = ((s4 == 8'd154) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[154] = ((s5 == 8'd154) & bht_update_p0);
        assign s12[154] = ((s6 == 8'd154) & bht_update_p1);
        assign s7[155] = ((s3 == 8'd155) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[155] = ((s4 == 8'd155) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[155] = ((s3 == 8'd155) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[155] = ((s4 == 8'd155) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[155] = ((s5 == 8'd155) & bht_update_p0);
        assign s12[155] = ((s6 == 8'd155) & bht_update_p1);
        assign s7[156] = ((s3 == 8'd156) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[156] = ((s4 == 8'd156) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[156] = ((s3 == 8'd156) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[156] = ((s4 == 8'd156) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[156] = ((s5 == 8'd156) & bht_update_p0);
        assign s12[156] = ((s6 == 8'd156) & bht_update_p1);
        assign s7[157] = ((s3 == 8'd157) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[157] = ((s4 == 8'd157) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[157] = ((s3 == 8'd157) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[157] = ((s4 == 8'd157) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[157] = ((s5 == 8'd157) & bht_update_p0);
        assign s12[157] = ((s6 == 8'd157) & bht_update_p1);
        assign s7[158] = ((s3 == 8'd158) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[158] = ((s4 == 8'd158) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[158] = ((s3 == 8'd158) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[158] = ((s4 == 8'd158) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[158] = ((s5 == 8'd158) & bht_update_p0);
        assign s12[158] = ((s6 == 8'd158) & bht_update_p1);
        assign s7[159] = ((s3 == 8'd159) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[159] = ((s4 == 8'd159) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[159] = ((s3 == 8'd159) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[159] = ((s4 == 8'd159) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[159] = ((s5 == 8'd159) & bht_update_p0);
        assign s12[159] = ((s6 == 8'd159) & bht_update_p1);
        assign s7[160] = ((s3 == 8'd160) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[160] = ((s4 == 8'd160) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[160] = ((s3 == 8'd160) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[160] = ((s4 == 8'd160) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[160] = ((s5 == 8'd160) & bht_update_p0);
        assign s12[160] = ((s6 == 8'd160) & bht_update_p1);
        assign s7[161] = ((s3 == 8'd161) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[161] = ((s4 == 8'd161) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[161] = ((s3 == 8'd161) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[161] = ((s4 == 8'd161) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[161] = ((s5 == 8'd161) & bht_update_p0);
        assign s12[161] = ((s6 == 8'd161) & bht_update_p1);
        assign s7[162] = ((s3 == 8'd162) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[162] = ((s4 == 8'd162) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[162] = ((s3 == 8'd162) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[162] = ((s4 == 8'd162) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[162] = ((s5 == 8'd162) & bht_update_p0);
        assign s12[162] = ((s6 == 8'd162) & bht_update_p1);
        assign s7[163] = ((s3 == 8'd163) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[163] = ((s4 == 8'd163) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[163] = ((s3 == 8'd163) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[163] = ((s4 == 8'd163) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[163] = ((s5 == 8'd163) & bht_update_p0);
        assign s12[163] = ((s6 == 8'd163) & bht_update_p1);
        assign s7[164] = ((s3 == 8'd164) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[164] = ((s4 == 8'd164) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[164] = ((s3 == 8'd164) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[164] = ((s4 == 8'd164) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[164] = ((s5 == 8'd164) & bht_update_p0);
        assign s12[164] = ((s6 == 8'd164) & bht_update_p1);
        assign s7[165] = ((s3 == 8'd165) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[165] = ((s4 == 8'd165) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[165] = ((s3 == 8'd165) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[165] = ((s4 == 8'd165) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[165] = ((s5 == 8'd165) & bht_update_p0);
        assign s12[165] = ((s6 == 8'd165) & bht_update_p1);
        assign s7[166] = ((s3 == 8'd166) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[166] = ((s4 == 8'd166) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[166] = ((s3 == 8'd166) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[166] = ((s4 == 8'd166) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[166] = ((s5 == 8'd166) & bht_update_p0);
        assign s12[166] = ((s6 == 8'd166) & bht_update_p1);
        assign s7[167] = ((s3 == 8'd167) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[167] = ((s4 == 8'd167) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[167] = ((s3 == 8'd167) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[167] = ((s4 == 8'd167) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[167] = ((s5 == 8'd167) & bht_update_p0);
        assign s12[167] = ((s6 == 8'd167) & bht_update_p1);
        assign s7[168] = ((s3 == 8'd168) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[168] = ((s4 == 8'd168) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[168] = ((s3 == 8'd168) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[168] = ((s4 == 8'd168) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[168] = ((s5 == 8'd168) & bht_update_p0);
        assign s12[168] = ((s6 == 8'd168) & bht_update_p1);
        assign s7[169] = ((s3 == 8'd169) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[169] = ((s4 == 8'd169) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[169] = ((s3 == 8'd169) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[169] = ((s4 == 8'd169) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[169] = ((s5 == 8'd169) & bht_update_p0);
        assign s12[169] = ((s6 == 8'd169) & bht_update_p1);
        assign s7[170] = ((s3 == 8'd170) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[170] = ((s4 == 8'd170) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[170] = ((s3 == 8'd170) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[170] = ((s4 == 8'd170) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[170] = ((s5 == 8'd170) & bht_update_p0);
        assign s12[170] = ((s6 == 8'd170) & bht_update_p1);
        assign s7[171] = ((s3 == 8'd171) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[171] = ((s4 == 8'd171) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[171] = ((s3 == 8'd171) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[171] = ((s4 == 8'd171) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[171] = ((s5 == 8'd171) & bht_update_p0);
        assign s12[171] = ((s6 == 8'd171) & bht_update_p1);
        assign s7[172] = ((s3 == 8'd172) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[172] = ((s4 == 8'd172) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[172] = ((s3 == 8'd172) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[172] = ((s4 == 8'd172) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[172] = ((s5 == 8'd172) & bht_update_p0);
        assign s12[172] = ((s6 == 8'd172) & bht_update_p1);
        assign s7[173] = ((s3 == 8'd173) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[173] = ((s4 == 8'd173) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[173] = ((s3 == 8'd173) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[173] = ((s4 == 8'd173) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[173] = ((s5 == 8'd173) & bht_update_p0);
        assign s12[173] = ((s6 == 8'd173) & bht_update_p1);
        assign s7[174] = ((s3 == 8'd174) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[174] = ((s4 == 8'd174) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[174] = ((s3 == 8'd174) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[174] = ((s4 == 8'd174) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[174] = ((s5 == 8'd174) & bht_update_p0);
        assign s12[174] = ((s6 == 8'd174) & bht_update_p1);
        assign s7[175] = ((s3 == 8'd175) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[175] = ((s4 == 8'd175) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[175] = ((s3 == 8'd175) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[175] = ((s4 == 8'd175) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[175] = ((s5 == 8'd175) & bht_update_p0);
        assign s12[175] = ((s6 == 8'd175) & bht_update_p1);
        assign s7[176] = ((s3 == 8'd176) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[176] = ((s4 == 8'd176) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[176] = ((s3 == 8'd176) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[176] = ((s4 == 8'd176) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[176] = ((s5 == 8'd176) & bht_update_p0);
        assign s12[176] = ((s6 == 8'd176) & bht_update_p1);
        assign s7[177] = ((s3 == 8'd177) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[177] = ((s4 == 8'd177) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[177] = ((s3 == 8'd177) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[177] = ((s4 == 8'd177) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[177] = ((s5 == 8'd177) & bht_update_p0);
        assign s12[177] = ((s6 == 8'd177) & bht_update_p1);
        assign s7[178] = ((s3 == 8'd178) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[178] = ((s4 == 8'd178) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[178] = ((s3 == 8'd178) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[178] = ((s4 == 8'd178) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[178] = ((s5 == 8'd178) & bht_update_p0);
        assign s12[178] = ((s6 == 8'd178) & bht_update_p1);
        assign s7[179] = ((s3 == 8'd179) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[179] = ((s4 == 8'd179) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[179] = ((s3 == 8'd179) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[179] = ((s4 == 8'd179) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[179] = ((s5 == 8'd179) & bht_update_p0);
        assign s12[179] = ((s6 == 8'd179) & bht_update_p1);
        assign s7[180] = ((s3 == 8'd180) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[180] = ((s4 == 8'd180) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[180] = ((s3 == 8'd180) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[180] = ((s4 == 8'd180) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[180] = ((s5 == 8'd180) & bht_update_p0);
        assign s12[180] = ((s6 == 8'd180) & bht_update_p1);
        assign s7[181] = ((s3 == 8'd181) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[181] = ((s4 == 8'd181) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[181] = ((s3 == 8'd181) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[181] = ((s4 == 8'd181) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[181] = ((s5 == 8'd181) & bht_update_p0);
        assign s12[181] = ((s6 == 8'd181) & bht_update_p1);
        assign s7[182] = ((s3 == 8'd182) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[182] = ((s4 == 8'd182) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[182] = ((s3 == 8'd182) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[182] = ((s4 == 8'd182) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[182] = ((s5 == 8'd182) & bht_update_p0);
        assign s12[182] = ((s6 == 8'd182) & bht_update_p1);
        assign s7[183] = ((s3 == 8'd183) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[183] = ((s4 == 8'd183) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[183] = ((s3 == 8'd183) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[183] = ((s4 == 8'd183) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[183] = ((s5 == 8'd183) & bht_update_p0);
        assign s12[183] = ((s6 == 8'd183) & bht_update_p1);
        assign s7[184] = ((s3 == 8'd184) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[184] = ((s4 == 8'd184) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[184] = ((s3 == 8'd184) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[184] = ((s4 == 8'd184) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[184] = ((s5 == 8'd184) & bht_update_p0);
        assign s12[184] = ((s6 == 8'd184) & bht_update_p1);
        assign s7[185] = ((s3 == 8'd185) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[185] = ((s4 == 8'd185) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[185] = ((s3 == 8'd185) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[185] = ((s4 == 8'd185) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[185] = ((s5 == 8'd185) & bht_update_p0);
        assign s12[185] = ((s6 == 8'd185) & bht_update_p1);
        assign s7[186] = ((s3 == 8'd186) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[186] = ((s4 == 8'd186) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[186] = ((s3 == 8'd186) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[186] = ((s4 == 8'd186) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[186] = ((s5 == 8'd186) & bht_update_p0);
        assign s12[186] = ((s6 == 8'd186) & bht_update_p1);
        assign s7[187] = ((s3 == 8'd187) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[187] = ((s4 == 8'd187) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[187] = ((s3 == 8'd187) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[187] = ((s4 == 8'd187) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[187] = ((s5 == 8'd187) & bht_update_p0);
        assign s12[187] = ((s6 == 8'd187) & bht_update_p1);
        assign s7[188] = ((s3 == 8'd188) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[188] = ((s4 == 8'd188) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[188] = ((s3 == 8'd188) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[188] = ((s4 == 8'd188) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[188] = ((s5 == 8'd188) & bht_update_p0);
        assign s12[188] = ((s6 == 8'd188) & bht_update_p1);
        assign s7[189] = ((s3 == 8'd189) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[189] = ((s4 == 8'd189) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[189] = ((s3 == 8'd189) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[189] = ((s4 == 8'd189) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[189] = ((s5 == 8'd189) & bht_update_p0);
        assign s12[189] = ((s6 == 8'd189) & bht_update_p1);
        assign s7[190] = ((s3 == 8'd190) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[190] = ((s4 == 8'd190) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[190] = ((s3 == 8'd190) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[190] = ((s4 == 8'd190) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[190] = ((s5 == 8'd190) & bht_update_p0);
        assign s12[190] = ((s6 == 8'd190) & bht_update_p1);
        assign s7[191] = ((s3 == 8'd191) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[191] = ((s4 == 8'd191) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[191] = ((s3 == 8'd191) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[191] = ((s4 == 8'd191) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[191] = ((s5 == 8'd191) & bht_update_p0);
        assign s12[191] = ((s6 == 8'd191) & bht_update_p1);
        assign s7[192] = ((s3 == 8'd192) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[192] = ((s4 == 8'd192) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[192] = ((s3 == 8'd192) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[192] = ((s4 == 8'd192) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[192] = ((s5 == 8'd192) & bht_update_p0);
        assign s12[192] = ((s6 == 8'd192) & bht_update_p1);
        assign s7[193] = ((s3 == 8'd193) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[193] = ((s4 == 8'd193) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[193] = ((s3 == 8'd193) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[193] = ((s4 == 8'd193) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[193] = ((s5 == 8'd193) & bht_update_p0);
        assign s12[193] = ((s6 == 8'd193) & bht_update_p1);
        assign s7[194] = ((s3 == 8'd194) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[194] = ((s4 == 8'd194) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[194] = ((s3 == 8'd194) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[194] = ((s4 == 8'd194) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[194] = ((s5 == 8'd194) & bht_update_p0);
        assign s12[194] = ((s6 == 8'd194) & bht_update_p1);
        assign s7[195] = ((s3 == 8'd195) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[195] = ((s4 == 8'd195) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[195] = ((s3 == 8'd195) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[195] = ((s4 == 8'd195) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[195] = ((s5 == 8'd195) & bht_update_p0);
        assign s12[195] = ((s6 == 8'd195) & bht_update_p1);
        assign s7[196] = ((s3 == 8'd196) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[196] = ((s4 == 8'd196) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[196] = ((s3 == 8'd196) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[196] = ((s4 == 8'd196) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[196] = ((s5 == 8'd196) & bht_update_p0);
        assign s12[196] = ((s6 == 8'd196) & bht_update_p1);
        assign s7[197] = ((s3 == 8'd197) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[197] = ((s4 == 8'd197) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[197] = ((s3 == 8'd197) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[197] = ((s4 == 8'd197) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[197] = ((s5 == 8'd197) & bht_update_p0);
        assign s12[197] = ((s6 == 8'd197) & bht_update_p1);
        assign s7[198] = ((s3 == 8'd198) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[198] = ((s4 == 8'd198) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[198] = ((s3 == 8'd198) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[198] = ((s4 == 8'd198) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[198] = ((s5 == 8'd198) & bht_update_p0);
        assign s12[198] = ((s6 == 8'd198) & bht_update_p1);
        assign s7[199] = ((s3 == 8'd199) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[199] = ((s4 == 8'd199) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[199] = ((s3 == 8'd199) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[199] = ((s4 == 8'd199) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[199] = ((s5 == 8'd199) & bht_update_p0);
        assign s12[199] = ((s6 == 8'd199) & bht_update_p1);
        assign s7[200] = ((s3 == 8'd200) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[200] = ((s4 == 8'd200) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[200] = ((s3 == 8'd200) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[200] = ((s4 == 8'd200) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[200] = ((s5 == 8'd200) & bht_update_p0);
        assign s12[200] = ((s6 == 8'd200) & bht_update_p1);
        assign s7[201] = ((s3 == 8'd201) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[201] = ((s4 == 8'd201) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[201] = ((s3 == 8'd201) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[201] = ((s4 == 8'd201) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[201] = ((s5 == 8'd201) & bht_update_p0);
        assign s12[201] = ((s6 == 8'd201) & bht_update_p1);
        assign s7[202] = ((s3 == 8'd202) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[202] = ((s4 == 8'd202) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[202] = ((s3 == 8'd202) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[202] = ((s4 == 8'd202) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[202] = ((s5 == 8'd202) & bht_update_p0);
        assign s12[202] = ((s6 == 8'd202) & bht_update_p1);
        assign s7[203] = ((s3 == 8'd203) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[203] = ((s4 == 8'd203) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[203] = ((s3 == 8'd203) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[203] = ((s4 == 8'd203) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[203] = ((s5 == 8'd203) & bht_update_p0);
        assign s12[203] = ((s6 == 8'd203) & bht_update_p1);
        assign s7[204] = ((s3 == 8'd204) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[204] = ((s4 == 8'd204) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[204] = ((s3 == 8'd204) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[204] = ((s4 == 8'd204) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[204] = ((s5 == 8'd204) & bht_update_p0);
        assign s12[204] = ((s6 == 8'd204) & bht_update_p1);
        assign s7[205] = ((s3 == 8'd205) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[205] = ((s4 == 8'd205) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[205] = ((s3 == 8'd205) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[205] = ((s4 == 8'd205) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[205] = ((s5 == 8'd205) & bht_update_p0);
        assign s12[205] = ((s6 == 8'd205) & bht_update_p1);
        assign s7[206] = ((s3 == 8'd206) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[206] = ((s4 == 8'd206) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[206] = ((s3 == 8'd206) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[206] = ((s4 == 8'd206) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[206] = ((s5 == 8'd206) & bht_update_p0);
        assign s12[206] = ((s6 == 8'd206) & bht_update_p1);
        assign s7[207] = ((s3 == 8'd207) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[207] = ((s4 == 8'd207) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[207] = ((s3 == 8'd207) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[207] = ((s4 == 8'd207) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[207] = ((s5 == 8'd207) & bht_update_p0);
        assign s12[207] = ((s6 == 8'd207) & bht_update_p1);
        assign s7[208] = ((s3 == 8'd208) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[208] = ((s4 == 8'd208) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[208] = ((s3 == 8'd208) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[208] = ((s4 == 8'd208) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[208] = ((s5 == 8'd208) & bht_update_p0);
        assign s12[208] = ((s6 == 8'd208) & bht_update_p1);
        assign s7[209] = ((s3 == 8'd209) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[209] = ((s4 == 8'd209) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[209] = ((s3 == 8'd209) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[209] = ((s4 == 8'd209) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[209] = ((s5 == 8'd209) & bht_update_p0);
        assign s12[209] = ((s6 == 8'd209) & bht_update_p1);
        assign s7[210] = ((s3 == 8'd210) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[210] = ((s4 == 8'd210) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[210] = ((s3 == 8'd210) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[210] = ((s4 == 8'd210) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[210] = ((s5 == 8'd210) & bht_update_p0);
        assign s12[210] = ((s6 == 8'd210) & bht_update_p1);
        assign s7[211] = ((s3 == 8'd211) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[211] = ((s4 == 8'd211) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[211] = ((s3 == 8'd211) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[211] = ((s4 == 8'd211) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[211] = ((s5 == 8'd211) & bht_update_p0);
        assign s12[211] = ((s6 == 8'd211) & bht_update_p1);
        assign s7[212] = ((s3 == 8'd212) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[212] = ((s4 == 8'd212) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[212] = ((s3 == 8'd212) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[212] = ((s4 == 8'd212) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[212] = ((s5 == 8'd212) & bht_update_p0);
        assign s12[212] = ((s6 == 8'd212) & bht_update_p1);
        assign s7[213] = ((s3 == 8'd213) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[213] = ((s4 == 8'd213) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[213] = ((s3 == 8'd213) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[213] = ((s4 == 8'd213) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[213] = ((s5 == 8'd213) & bht_update_p0);
        assign s12[213] = ((s6 == 8'd213) & bht_update_p1);
        assign s7[214] = ((s3 == 8'd214) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[214] = ((s4 == 8'd214) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[214] = ((s3 == 8'd214) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[214] = ((s4 == 8'd214) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[214] = ((s5 == 8'd214) & bht_update_p0);
        assign s12[214] = ((s6 == 8'd214) & bht_update_p1);
        assign s7[215] = ((s3 == 8'd215) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[215] = ((s4 == 8'd215) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[215] = ((s3 == 8'd215) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[215] = ((s4 == 8'd215) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[215] = ((s5 == 8'd215) & bht_update_p0);
        assign s12[215] = ((s6 == 8'd215) & bht_update_p1);
        assign s7[216] = ((s3 == 8'd216) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[216] = ((s4 == 8'd216) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[216] = ((s3 == 8'd216) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[216] = ((s4 == 8'd216) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[216] = ((s5 == 8'd216) & bht_update_p0);
        assign s12[216] = ((s6 == 8'd216) & bht_update_p1);
        assign s7[217] = ((s3 == 8'd217) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[217] = ((s4 == 8'd217) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[217] = ((s3 == 8'd217) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[217] = ((s4 == 8'd217) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[217] = ((s5 == 8'd217) & bht_update_p0);
        assign s12[217] = ((s6 == 8'd217) & bht_update_p1);
        assign s7[218] = ((s3 == 8'd218) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[218] = ((s4 == 8'd218) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[218] = ((s3 == 8'd218) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[218] = ((s4 == 8'd218) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[218] = ((s5 == 8'd218) & bht_update_p0);
        assign s12[218] = ((s6 == 8'd218) & bht_update_p1);
        assign s7[219] = ((s3 == 8'd219) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[219] = ((s4 == 8'd219) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[219] = ((s3 == 8'd219) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[219] = ((s4 == 8'd219) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[219] = ((s5 == 8'd219) & bht_update_p0);
        assign s12[219] = ((s6 == 8'd219) & bht_update_p1);
        assign s7[220] = ((s3 == 8'd220) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[220] = ((s4 == 8'd220) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[220] = ((s3 == 8'd220) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[220] = ((s4 == 8'd220) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[220] = ((s5 == 8'd220) & bht_update_p0);
        assign s12[220] = ((s6 == 8'd220) & bht_update_p1);
        assign s7[221] = ((s3 == 8'd221) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[221] = ((s4 == 8'd221) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[221] = ((s3 == 8'd221) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[221] = ((s4 == 8'd221) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[221] = ((s5 == 8'd221) & bht_update_p0);
        assign s12[221] = ((s6 == 8'd221) & bht_update_p1);
        assign s7[222] = ((s3 == 8'd222) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[222] = ((s4 == 8'd222) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[222] = ((s3 == 8'd222) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[222] = ((s4 == 8'd222) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[222] = ((s5 == 8'd222) & bht_update_p0);
        assign s12[222] = ((s6 == 8'd222) & bht_update_p1);
        assign s7[223] = ((s3 == 8'd223) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[223] = ((s4 == 8'd223) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[223] = ((s3 == 8'd223) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[223] = ((s4 == 8'd223) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[223] = ((s5 == 8'd223) & bht_update_p0);
        assign s12[223] = ((s6 == 8'd223) & bht_update_p1);
        assign s7[224] = ((s3 == 8'd224) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[224] = ((s4 == 8'd224) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[224] = ((s3 == 8'd224) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[224] = ((s4 == 8'd224) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[224] = ((s5 == 8'd224) & bht_update_p0);
        assign s12[224] = ((s6 == 8'd224) & bht_update_p1);
        assign s7[225] = ((s3 == 8'd225) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[225] = ((s4 == 8'd225) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[225] = ((s3 == 8'd225) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[225] = ((s4 == 8'd225) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[225] = ((s5 == 8'd225) & bht_update_p0);
        assign s12[225] = ((s6 == 8'd225) & bht_update_p1);
        assign s7[226] = ((s3 == 8'd226) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[226] = ((s4 == 8'd226) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[226] = ((s3 == 8'd226) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[226] = ((s4 == 8'd226) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[226] = ((s5 == 8'd226) & bht_update_p0);
        assign s12[226] = ((s6 == 8'd226) & bht_update_p1);
        assign s7[227] = ((s3 == 8'd227) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[227] = ((s4 == 8'd227) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[227] = ((s3 == 8'd227) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[227] = ((s4 == 8'd227) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[227] = ((s5 == 8'd227) & bht_update_p0);
        assign s12[227] = ((s6 == 8'd227) & bht_update_p1);
        assign s7[228] = ((s3 == 8'd228) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[228] = ((s4 == 8'd228) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[228] = ((s3 == 8'd228) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[228] = ((s4 == 8'd228) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[228] = ((s5 == 8'd228) & bht_update_p0);
        assign s12[228] = ((s6 == 8'd228) & bht_update_p1);
        assign s7[229] = ((s3 == 8'd229) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[229] = ((s4 == 8'd229) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[229] = ((s3 == 8'd229) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[229] = ((s4 == 8'd229) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[229] = ((s5 == 8'd229) & bht_update_p0);
        assign s12[229] = ((s6 == 8'd229) & bht_update_p1);
        assign s7[230] = ((s3 == 8'd230) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[230] = ((s4 == 8'd230) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[230] = ((s3 == 8'd230) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[230] = ((s4 == 8'd230) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[230] = ((s5 == 8'd230) & bht_update_p0);
        assign s12[230] = ((s6 == 8'd230) & bht_update_p1);
        assign s7[231] = ((s3 == 8'd231) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[231] = ((s4 == 8'd231) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[231] = ((s3 == 8'd231) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[231] = ((s4 == 8'd231) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[231] = ((s5 == 8'd231) & bht_update_p0);
        assign s12[231] = ((s6 == 8'd231) & bht_update_p1);
        assign s7[232] = ((s3 == 8'd232) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[232] = ((s4 == 8'd232) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[232] = ((s3 == 8'd232) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[232] = ((s4 == 8'd232) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[232] = ((s5 == 8'd232) & bht_update_p0);
        assign s12[232] = ((s6 == 8'd232) & bht_update_p1);
        assign s7[233] = ((s3 == 8'd233) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[233] = ((s4 == 8'd233) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[233] = ((s3 == 8'd233) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[233] = ((s4 == 8'd233) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[233] = ((s5 == 8'd233) & bht_update_p0);
        assign s12[233] = ((s6 == 8'd233) & bht_update_p1);
        assign s7[234] = ((s3 == 8'd234) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[234] = ((s4 == 8'd234) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[234] = ((s3 == 8'd234) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[234] = ((s4 == 8'd234) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[234] = ((s5 == 8'd234) & bht_update_p0);
        assign s12[234] = ((s6 == 8'd234) & bht_update_p1);
        assign s7[235] = ((s3 == 8'd235) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[235] = ((s4 == 8'd235) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[235] = ((s3 == 8'd235) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[235] = ((s4 == 8'd235) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[235] = ((s5 == 8'd235) & bht_update_p0);
        assign s12[235] = ((s6 == 8'd235) & bht_update_p1);
        assign s7[236] = ((s3 == 8'd236) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[236] = ((s4 == 8'd236) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[236] = ((s3 == 8'd236) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[236] = ((s4 == 8'd236) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[236] = ((s5 == 8'd236) & bht_update_p0);
        assign s12[236] = ((s6 == 8'd236) & bht_update_p1);
        assign s7[237] = ((s3 == 8'd237) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[237] = ((s4 == 8'd237) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[237] = ((s3 == 8'd237) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[237] = ((s4 == 8'd237) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[237] = ((s5 == 8'd237) & bht_update_p0);
        assign s12[237] = ((s6 == 8'd237) & bht_update_p1);
        assign s7[238] = ((s3 == 8'd238) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[238] = ((s4 == 8'd238) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[238] = ((s3 == 8'd238) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[238] = ((s4 == 8'd238) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[238] = ((s5 == 8'd238) & bht_update_p0);
        assign s12[238] = ((s6 == 8'd238) & bht_update_p1);
        assign s7[239] = ((s3 == 8'd239) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[239] = ((s4 == 8'd239) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[239] = ((s3 == 8'd239) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[239] = ((s4 == 8'd239) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[239] = ((s5 == 8'd239) & bht_update_p0);
        assign s12[239] = ((s6 == 8'd239) & bht_update_p1);
        assign s7[240] = ((s3 == 8'd240) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[240] = ((s4 == 8'd240) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[240] = ((s3 == 8'd240) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[240] = ((s4 == 8'd240) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[240] = ((s5 == 8'd240) & bht_update_p0);
        assign s12[240] = ((s6 == 8'd240) & bht_update_p1);
        assign s7[241] = ((s3 == 8'd241) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[241] = ((s4 == 8'd241) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[241] = ((s3 == 8'd241) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[241] = ((s4 == 8'd241) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[241] = ((s5 == 8'd241) & bht_update_p0);
        assign s12[241] = ((s6 == 8'd241) & bht_update_p1);
        assign s7[242] = ((s3 == 8'd242) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[242] = ((s4 == 8'd242) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[242] = ((s3 == 8'd242) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[242] = ((s4 == 8'd242) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[242] = ((s5 == 8'd242) & bht_update_p0);
        assign s12[242] = ((s6 == 8'd242) & bht_update_p1);
        assign s7[243] = ((s3 == 8'd243) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[243] = ((s4 == 8'd243) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[243] = ((s3 == 8'd243) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[243] = ((s4 == 8'd243) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[243] = ((s5 == 8'd243) & bht_update_p0);
        assign s12[243] = ((s6 == 8'd243) & bht_update_p1);
        assign s7[244] = ((s3 == 8'd244) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[244] = ((s4 == 8'd244) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[244] = ((s3 == 8'd244) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[244] = ((s4 == 8'd244) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[244] = ((s5 == 8'd244) & bht_update_p0);
        assign s12[244] = ((s6 == 8'd244) & bht_update_p1);
        assign s7[245] = ((s3 == 8'd245) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[245] = ((s4 == 8'd245) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[245] = ((s3 == 8'd245) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[245] = ((s4 == 8'd245) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[245] = ((s5 == 8'd245) & bht_update_p0);
        assign s12[245] = ((s6 == 8'd245) & bht_update_p1);
        assign s7[246] = ((s3 == 8'd246) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[246] = ((s4 == 8'd246) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[246] = ((s3 == 8'd246) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[246] = ((s4 == 8'd246) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[246] = ((s5 == 8'd246) & bht_update_p0);
        assign s12[246] = ((s6 == 8'd246) & bht_update_p1);
        assign s7[247] = ((s3 == 8'd247) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[247] = ((s4 == 8'd247) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[247] = ((s3 == 8'd247) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[247] = ((s4 == 8'd247) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[247] = ((s5 == 8'd247) & bht_update_p0);
        assign s12[247] = ((s6 == 8'd247) & bht_update_p1);
        assign s7[248] = ((s3 == 8'd248) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[248] = ((s4 == 8'd248) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[248] = ((s3 == 8'd248) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[248] = ((s4 == 8'd248) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[248] = ((s5 == 8'd248) & bht_update_p0);
        assign s12[248] = ((s6 == 8'd248) & bht_update_p1);
        assign s7[249] = ((s3 == 8'd249) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[249] = ((s4 == 8'd249) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[249] = ((s3 == 8'd249) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[249] = ((s4 == 8'd249) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[249] = ((s5 == 8'd249) & bht_update_p0);
        assign s12[249] = ((s6 == 8'd249) & bht_update_p1);
        assign s7[250] = ((s3 == 8'd250) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[250] = ((s4 == 8'd250) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[250] = ((s3 == 8'd250) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[250] = ((s4 == 8'd250) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[250] = ((s5 == 8'd250) & bht_update_p0);
        assign s12[250] = ((s6 == 8'd250) & bht_update_p1);
        assign s7[251] = ((s3 == 8'd251) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[251] = ((s4 == 8'd251) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[251] = ((s3 == 8'd251) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[251] = ((s4 == 8'd251) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[251] = ((s5 == 8'd251) & bht_update_p0);
        assign s12[251] = ((s6 == 8'd251) & bht_update_p1);
        assign s7[252] = ((s3 == 8'd252) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[252] = ((s4 == 8'd252) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[252] = ((s3 == 8'd252) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[252] = ((s4 == 8'd252) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[252] = ((s5 == 8'd252) & bht_update_p0);
        assign s12[252] = ((s6 == 8'd252) & bht_update_p1);
        assign s7[253] = ((s3 == 8'd253) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[253] = ((s4 == 8'd253) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[253] = ((s3 == 8'd253) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[253] = ((s4 == 8'd253) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[253] = ((s5 == 8'd253) & bht_update_p0);
        assign s12[253] = ((s6 == 8'd253) & bht_update_p1);
        assign s7[254] = ((s3 == 8'd254) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[254] = ((s4 == 8'd254) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[254] = ((s3 == 8'd254) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[254] = ((s4 == 8'd254) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[254] = ((s5 == 8'd254) & bht_update_p0);
        assign s12[254] = ((s6 == 8'd254) & bht_update_p1);
        assign s7[255] = ((s3 == 8'd255) & bht_update_p0 & bht_update_p0_sel_data[1]);
        assign s8[255] = ((s4 == 8'd255) & bht_update_p1 & bht_update_p1_sel_data[1]);
        assign s9[255] = ((s3 == 8'd255) & bht_update_p0 & ~bht_update_p0_sel_data[1]);
        assign s10[255] = ((s4 == 8'd255) & bht_update_p1 & ~bht_update_p1_sel_data[1]);
        assign s11[255] = ((s5 == 8'd255) & bht_update_p0);
        assign s12[255] = ((s6 == 8'd255) & bht_update_p1);
        integer s13;
        wire s14;
        wire s15;
        wire s16;
        assign s14 = bht_update_p0 & (bht_update_p0_sel_data[1]) & bht_update_p1 & (bht_update_p1_sel_data[1]) & (s3 == s4);
        assign s15 = bht_update_p0 & ~(bht_update_p0_sel_data[1]) & bht_update_p1 & ~(bht_update_p1_sel_data[1]) & (s3 == s4);
        assign s16 = bht_update_p0 & bht_update_p1 & (s6 == s5);
        wire s17 = (bht_update_p0 & (bht_update_p0_sel_data[1])) | (bht_update_p1 & (bht_update_p1_sel_data[1]));
        always @(posedge core_clk or negedge core_reset_n) begin
            if (!core_reset_n) begin
                for (s13 = 0; s13 < 256; s13 = s13 + 1) begin
                    s0[s13] <= 2'b01;
                end
            end
            else if (s17) begin
                for (s13 = 0; s13 < 256; s13 = s13 + 1) begin
                    if (s7[s13] | s8[s13]) begin
                        s0[s13] <= s14 ? bht_update_p1_dir_data : (({2{s7[s13]}} & bht_update_p0_dir_data) | ({2{s8[s13]}} & bht_update_p1_dir_data));
                    end
                end
            end
        end

        integer s18;
        wire s19 = (bht_update_p0 & ~(bht_update_p0_sel_data[1])) | (bht_update_p1 & ~(bht_update_p1_sel_data[1]));
        always @(posedge core_clk or negedge core_reset_n) begin
            if (!core_reset_n) begin
                for (s18 = 0; s18 < 256; s18 = s18 + 1) begin
                    s1[s18] <= 2'b01;
                end
            end
            else if (s19) begin
                for (s18 = 0; s18 < 256; s18 = s18 + 1) begin
                    if (s9[s18] | s10[s18]) begin
                        s1[s18] <= s15 ? bht_update_p1_dir_data : (({2{s9[s18]}} & bht_update_p0_dir_data) | ({2{s10[s18]}} & bht_update_p1_dir_data));
                    end
                end
            end
        end

        integer s20;
        always @(posedge core_clk or negedge core_reset_n) begin
            if (!core_reset_n) begin
                for (s20 = 0; s20 < 256; s20 = s20 + 1) begin
                    s2[s20] <= 2'b01;
                end
            end
            else if (bht_update_p0 | bht_update_p1) begin
                for (s20 = 0; s20 < 256; s20 = s20 + 1) begin
                    if (s11[s20] | s12[s20]) begin
                        s2[s20] <= s16 ? bht_update_p1_sel_data : (({2{s11[s20]}} & bht_update_p0_sel_data) | ({2{s12[s20]}} & bht_update_p1_sel_data));
                    end
                end
            end
        end

        assign bht_taken_rdata = s0[bht_dir_rd_addr];
        assign bht_ntaken_rdata = s1[bht_dir_rd_addr];
        assign bht_sel_rdata = s2[bht_sel_rd_addr];
    end
    else begin:gen_bht_no
        assign bht_taken_rdata = 2'b0;
        assign bht_ntaken_rdata = 2'b0;
        assign bht_sel_rdata = 2'b0;
    end
endgenerate
endmodule

