library ieee;
use ieee.std_logic_1164.all;

entity top is
	 port( a: in std_logic_vector(31 downto 0);
	       result: out std_logic_vector(31 downto 0));
 end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059: std_logic;

begin

w0 <= a(4) and not a(5);
w1 <= not a(4) and a(5);
w2 <= not w0 and not w1;
w3 <= a(2) and not a(3);
w4 <= not a(2) and a(3);
w5 <= not w3 and not w4;
w6 <= w2 and not w5;
w7 <= not a(29) and a(30);
w8 <= a(29) and not a(30);
w9 <= not w7 and not w8;
w10 <= a(31) and not w9;
w11 <= not a(24) and not a(25);
w12 <= not a(23) and a(26);
w13 <= w11 and w12;
w14 <= a(27) and a(28);
w15 <= w8 and w14;
w16 <= w13 and w15;
w17 <= not a(27) and not a(28);
w18 <= w8 and w17;
w19 <= a(24) and a(25);
w20 <= w12 and w19;
w21 <= w18 and w20;
w22 <= not a(23) and not a(26);
w23 <= w11 and w22;
w24 <= a(29) and a(30);
w25 <= w14 and w24;
w26 <= w23 and w25;
w27 <= a(23) and not a(26);
w28 <= not a(24) and a(25);
w29 <= w27 and w28;
w30 <= w18 and w29;
w31 <= w19 and w27;
w32 <= not a(29) and not a(30);
w33 <= w17 and w32;
w34 <= w31 and w33;
w35 <= not w30 and not w34;
w36 <= w22 and w28;
w37 <= w25 and w36;
w38 <= a(27) and not a(28);
w39 <= w24 and w38;
w40 <= a(23) and a(26);
w41 <= w28 and w40;
w42 <= w39 and w41;
w43 <= not w37 and not w42;
w44 <= not a(27) and a(28);
w45 <= w7 and w44;
w46 <= w31 and w45;
w47 <= a(24) and not a(25);
w48 <= w27 and w47;
w49 <= w7 and w38;
w50 <= w48 and w49;
w51 <= not w46 and not w50;
w52 <= w17 and w24;
w53 <= w29 and w52;
w54 <= w18 and w41;
w55 <= not w53 and not w54;
w56 <= w23 and w52;
w57 <= w22 and w47;
w58 <= w45 and w57;
w59 <= w12 and w28;
w60 <= w18 and w59;
w61 <= w40 and w47;
w62 <= w18 and w61;
w63 <= not w60 and not w62;
w64 <= w32 and w44;
w65 <= w48 and w64;
w66 <= w11 and w27;
w67 <= w64 and w66;
w68 <= not w65 and not w67;
w69 <= w7 and w17;
w70 <= w48 and w69;
w71 <= w45 and w61;
w72 <= not w70 and not w71;
w73 <= w68 and w72;
w74 <= w63 and w73;
w75 <= not w58 and w74;
w76 <= not w56 and w75;
w77 <= w33 and w61;
w78 <= w14 and w32;
w79 <= w57 and w78;
w80 <= w13 and w78;
w81 <= w39 and w61;
w82 <= w13 and w52;
w83 <= w12 and w47;
w84 <= w52 and w83;
w85 <= w49 and w59;
w86 <= w49 and w57;
w87 <= w36 and w69;
w88 <= w7 and w14;
w89 <= w61 and w88;
w90 <= w52 and w59;
w91 <= not w89 and not w90;
w92 <= w29 and w64;
w93 <= w18 and w83;
w94 <= not w92 and not w93;
w95 <= w8 and w44;
w96 <= w29 and w95;
w97 <= w19 and w40;
w98 <= w64 and w97;
w99 <= w20 and w78;
w100 <= w59 and w78;
w101 <= w32 and w38;
w102 <= w59 and w101;
w103 <= w49 and w61;
w104 <= w20 and w88;
w105 <= w64 and w83;
w106 <= w49 and w66;
w107 <= not w105 and not w106;
w108 <= w23 and w78;
w109 <= w24 and w44;
w110 <= w41 and w109;
w111 <= w19 and w22;
w112 <= w52 and w111;
w113 <= not w110 and not w112;
w114 <= not w108 and w113;
w115 <= w107 and w114;
w116 <= not w104 and w115;
w117 <= not w103 and w116;
w118 <= not w102 and w117;
w119 <= not w100 and w118;
w120 <= not w99 and w119;
w121 <= not w98 and w120;
w122 <= not w96 and w121;
w123 <= w15 and w59;
w124 <= w41 and w49;
w125 <= w57 and w88;
w126 <= w33 and w97;
w127 <= w36 and w101;
w128 <= not w126 and not w127;
w129 <= w45 and w48;
w130 <= w128 and not w129;
w131 <= not w125 and w130;
w132 <= not w124 and w131;
w133 <= not w123 and w132;
w134 <= w8 and w38;
w135 <= w111 and w134;
w136 <= w61 and w134;
w137 <= not w135 and not w136;
w138 <= w61 and w109;
w139 <= w137 and not w138;
w140 <= w29 and w78;
w141 <= w25 and w83;
w142 <= not w140 and not w141;
w143 <= w139 and w142;
w144 <= w133 and w143;
w145 <= w122 and w144;
w146 <= w94 and w145;
w147 <= w91 and w146;
w148 <= not w87 and w147;
w149 <= not w86 and w148;
w150 <= not w85 and w149;
w151 <= not w84 and w150;
w152 <= not w82 and w151;
w153 <= not w81 and w152;
w154 <= not w80 and w153;
w155 <= not w79 and w154;
w156 <= not w77 and w155;
w157 <= w15 and w20;
w158 <= w52 and w97;
w159 <= w20 and w69;
w160 <= w23 and w134;
w161 <= w29 and w39;
w162 <= not w160 and not w161;
w163 <= w25 and w57;
w164 <= w13 and w88;
w165 <= not w163 and not w164;
w166 <= w15 and w41;
w167 <= w61 and w69;
w168 <= w13 and w109;
w169 <= not w167 and not w168;
w170 <= not w166 and w169;
w171 <= w20 and w45;
w172 <= w83 and w134;
w173 <= not w171 and not w172;
w174 <= w20 and w52;
w175 <= w78 and w83;
w176 <= not w174 and not w175;
w177 <= w88 and w111;
w178 <= w78 and w111;
w179 <= not w177 and not w178;
w180 <= w33 and w59;
w181 <= w61 and w101;
w182 <= not w180 and not w181;
w183 <= w39 and w97;
w184 <= w15 and w66;
w185 <= not w183 and not w184;
w186 <= w18 and w66;
w187 <= w41 and w134;
w188 <= not w186 and not w187;
w189 <= w49 and w111;
w190 <= w41 and w69;
w191 <= not w189 and not w190;
w192 <= w188 and w191;
w193 <= w185 and w192;
w194 <= w182 and w193;
w195 <= w179 and w194;
w196 <= w176 and w195;
w197 <= w173 and w196;
w198 <= w170 and w197;
w199 <= w165 and w198;
w200 <= w162 and w199;
w201 <= not w159 and w200;
w202 <= not w158 and w201;
w203 <= not w157 and w202;
w204 <= w11 and w40;
w205 <= w15 and w204;
w206 <= w18 and w23;
w207 <= w66 and w134;
w208 <= w61 and w64;
w209 <= w66 and w78;
w210 <= w48 and w52;
w211 <= w45 and w66;
w212 <= w31 and w95;
w213 <= w69 and w97;
w214 <= not w212 and not w213;
w215 <= w36 and w49;
w216 <= w31 and w69;
w217 <= not w215 and not w216;
w218 <= w33 and w66;
w219 <= w69 and w83;
w220 <= not w218 and not w219;
w221 <= w66 and w101;
w222 <= w25 and w29;
w223 <= not w221 and not w222;
w224 <= w29 and w69;
w225 <= w31 and w39;
w226 <= not w224 and not w225;
w227 <= w39 and w66;
w228 <= w18 and w97;
w229 <= not w227 and not w228;
w230 <= w59 and w95;
w231 <= w29 and w101;
w232 <= not w230 and not w231;
w233 <= w33 and w111;
w234 <= w52 and w66;
w235 <= not w233 and not w234;
w236 <= w45 and w111;
w237 <= w25 and w59;
w238 <= not w236 and not w237;
w239 <= w23 and w95;
w240 <= w39 and w204;
w241 <= w64 and w204;
w242 <= not w240 and not w241;
w243 <= not w239 and w242;
w244 <= w238 and w243;
w245 <= w235 and w244;
w246 <= w232 and w245;
w247 <= w229 and w246;
w248 <= w226 and w247;
w249 <= w223 and w248;
w250 <= w220 and w249;
w251 <= w217 and w250;
w252 <= w214 and w251;
w253 <= not w211 and w252;
w254 <= not w210 and w253;
w255 <= not w209 and w254;
w256 <= not w208 and w255;
w257 <= not w207 and w256;
w258 <= not w206 and w257;
w259 <= not w205 and w258;
w260 <= w18 and w36;
w261 <= w25 and w97;
w262 <= w97 and w109;
w263 <= w23 and w49;
w264 <= w13 and w69;
w265 <= w29 and w88;
w266 <= w97 and w101;
w267 <= w95 and w204;
w268 <= not w266 and not w267;
w269 <= w109 and w111;
w270 <= w29 and w49;
w271 <= not w269 and not w270;
w272 <= w15 and w36;
w273 <= w20 and w134;
w274 <= w36 and w109;
w275 <= w48 and w95;
w276 <= not w274 and not w275;
w277 <= not w273 and w276;
w278 <= not w272 and w277;
w279 <= w271 and w278;
w280 <= w268 and w279;
w281 <= not w265 and w280;
w282 <= not w264 and w281;
w283 <= not w263 and w282;
w284 <= not w262 and w283;
w285 <= not w261 and w284;
w286 <= not w260 and w285;
w287 <= w57 and w109;
w288 <= w69 and w111;
w289 <= w59 and w69;
w290 <= w69 and w204;
w291 <= not w289 and not w290;
w292 <= w25 and w204;
w293 <= w18 and w204;
w294 <= not w292 and not w293;
w295 <= w291 and w294;
w296 <= not w288 and w295;
w297 <= not w287 and w296;
w298 <= w15 and w29;
w299 <= w45 and w97;
w300 <= not w298 and not w299;
w301 <= w31 and w134;
w302 <= w39 and w48;
w303 <= w33 and w48;
w304 <= not w302 and not w303;
w305 <= not w301 and w304;
w306 <= w20 and w95;
w307 <= w23 and w33;
w308 <= not w306 and not w307;
w309 <= w25 and w31;
w310 <= w13 and w64;
w311 <= not w309 and not w310;
w312 <= w308 and w311;
w313 <= w305 and w312;
w314 <= w300 and w313;
w315 <= w297 and w314;
w316 <= w286 and w315;
w317 <= w259 and w316;
w318 <= w203 and w317;
w319 <= w156 and w318;
w320 <= w76 and w319;
w321 <= w55 and w320;
w322 <= w51 and w321;
w323 <= w43 and w322;
w324 <= w35 and w323;
w325 <= not w26 and w324;
w326 <= not w21 and w325;
w327 <= not w16 and w326;
w328 <= w20 and w64;
w329 <= w59 and w64;
w330 <= w25 and w48;
w331 <= w13 and w39;
w332 <= w41 and w45;
w333 <= w66 and w88;
w334 <= not w262 and not w333;
w335 <= w23 and w39;
w336 <= not w270 and not w335;
w337 <= w36 and w39;
w338 <= w39 and w83;
w339 <= not w337 and not w338;
w340 <= not w310 and w339;
w341 <= w336 and w340;
w342 <= w334 and w341;
w343 <= not w46 and w342;
w344 <= not w332 and w343;
w345 <= not w112 and w344;
w346 <= not w234 and w345;
w347 <= not w331 and w346;
w348 <= not w330 and w347;
w349 <= not w260 and w348;
w350 <= not w228 and w349;
w351 <= w13 and w25;
w352 <= w52 and w57;
w353 <= not w299 and not w352;
w354 <= w31 and w52;
w355 <= w41 and w88;
w356 <= not w354 and not w355;
w357 <= w33 and w83;
w358 <= not w81 and not w357;
w359 <= w36 and w78;
w360 <= w101 and w204;
w361 <= w49 and w83;
w362 <= w45 and w83;
w363 <= w15 and w111;
w364 <= w15 and w83;
w365 <= w83 and w101;
w366 <= not w79 and not w365;
w367 <= not w136 and w366;
w368 <= not w364 and w367;
w369 <= not w363 and w368;
w370 <= w52 and w204;
w371 <= w95 and w111;
w372 <= not w370 and not w371;
w373 <= w23 and w101;
w374 <= not w306 and not w373;
w375 <= w372 and w374;
w376 <= w369 and w375;
w377 <= not w362 and w376;
w378 <= not w129 and w377;
w379 <= not w361 and w378;
w380 <= not w215 and w379;
w381 <= not w302 and w380;
w382 <= not w360 and w381;
w383 <= not w359 and w382;
w384 <= w15 and w57;
w385 <= not w206 and not w384;
w386 <= w134 and w204;
w387 <= w20 and w33;
w388 <= w33 and w36;
w389 <= not w387 and not w388;
w390 <= not w224 and w389;
w391 <= not w227 and w390;
w392 <= not w221 and w391;
w393 <= not w160 and w392;
w394 <= not w386 and w393;
w395 <= w39 and w111;
w396 <= w20 and w39;
w397 <= w83 and w88;
w398 <= not w396 and not w397;
w399 <= not w395 and w398;
w400 <= not w218 and w399;
w401 <= w31 and w78;
w402 <= not w168 and not w401;
w403 <= w41 and w64;
w404 <= w29 and w45;
w405 <= w29 and w134;
w406 <= not w301 and not w405;
w407 <= not w404 and w406;
w408 <= not w403 and w407;
w409 <= w36 and w95;
w410 <= not w123 and not w409;
w411 <= w408 and w410;
w412 <= w402 and w411;
w413 <= w400 and w412;
w414 <= w394 and w413;
w415 <= w385 and w414;
w416 <= w383 and w415;
w417 <= w94 and w416;
w418 <= w358 and w417;
w419 <= w356 and w418;
w420 <= w353 and w419;
w421 <= not w189 and w420;
w422 <= not w351 and w421;
w423 <= not w272 and w422;
w424 <= w18 and w111;
w425 <= w25 and w41;
w426 <= not w424 and not w425;
w427 <= w101 and w111;
w428 <= w64 and w111;
w429 <= not w102 and not w428;
w430 <= w20 and w109;
w431 <= w13 and w101;
w432 <= not w430 and not w431;
w433 <= w429 and w432;
w434 <= not w177 and w433;
w435 <= not w124 and w434;
w436 <= not w225 and w435;
w437 <= not w427 and w436;
w438 <= not w166 and w437;
w439 <= w78 and w97;
w440 <= w31 and w101;
w441 <= w31 and w109;
w442 <= not w16 and not w441;
w443 <= not w210 and not w269;
w444 <= w36 and w88;
w445 <= not w70 and not w444;
w446 <= w49 and w204;
w447 <= not w183 and not w446;
w448 <= w39 and w59;
w449 <= w109 and w204;
w450 <= not w241 and not w292;
w451 <= not w96 and w450;
w452 <= not w267 and w451;
w453 <= w31 and w88;
w454 <= w57 and w95;
w455 <= not w453 and not w454;
w456 <= w452 and w455;
w457 <= not w449 and w456;
w458 <= not w448 and w457;
w459 <= not w209 and w458;
w460 <= w95 and w97;
w461 <= not w207 and not w460;
w462 <= w39 and w57;
w463 <= not w50 and not w240;
w464 <= not w462 and w463;
w465 <= not w62 and not w158;
w466 <= w36 and w134;
w467 <= w83 and w95;
w468 <= not w275 and not w467;
w469 <= not w466 and w468;
w470 <= not w273 and w469;
w471 <= w13 and w33;
w472 <= w33 and w57;
w473 <= not w303 and not w472;
w474 <= not w471 and w473;
w475 <= not w233 and w474;
w476 <= not w293 and w475;
w477 <= w470 and w476;
w478 <= w465 and w477;
w479 <= w464 and w478;
w480 <= w461 and w479;
w481 <= w459 and w480;
w482 <= w447 and w481;
w483 <= w445 and w482;
w484 <= w443 and w483;
w485 <= w442 and w484;
w486 <= w43 and w485;
w487 <= not w104 and w486;
w488 <= not w82 and w487;
w489 <= not w440 and w488;
w490 <= not w439 and w489;
w491 <= not w180 and w490;
w492 <= w23 and w69;
w493 <= w23 and w45;
w494 <= not w492 and not w493;
w495 <= not w161 and w494;
w496 <= not w212 and w495;
w497 <= w15 and w97;
w498 <= w20 and w101;
w499 <= w13 and w95;
w500 <= not w498 and not w499;
w501 <= not w497 and w500;
w502 <= w33 and w204;
w503 <= w57 and w101;
w504 <= w18 and w57;
w505 <= not w503 and not w504;
w506 <= w23 and w109;
w507 <= w505 and not w506;
w508 <= not w502 and w507;
w509 <= w501 and w508;
w510 <= w496 and w509;
w511 <= w491 and w510;
w512 <= w438 and w511;
w513 <= w426 and w512;
w514 <= w423 and w513;
w515 <= w350 and w514;
w516 <= w128 and w515;
w517 <= not w87 and w516;
w518 <= not w237 and w517;
w519 <= not w178 and w518;
w520 <= not w329 and w519;
w521 <= not w328 and w520;
w522 <= not w184 and w521;
w523 <= not w327 and not w522;
w524 <= w31 and w64;
w525 <= not w123 and not w157;
w526 <= not w129 and not w425;
w527 <= w59 and w134;
w528 <= not w163 and not w527;
w529 <= w52 and w61;
w530 <= not w140 and not w529;
w531 <= w528 and w530;
w532 <= not w71 and w531;
w533 <= not w112 and w532;
w534 <= not w329 and w533;
w535 <= not w54 and w534;
w536 <= w41 and w78;
w537 <= w49 and w97;
w538 <= w36 and w64;
w539 <= not w428 and not w538;
w540 <= w294 and w539;
w541 <= not w537 and w540;
w542 <= not w234 and w541;
w543 <= not w42 and w542;
w544 <= not w178 and w543;
w545 <= not w536 and w544;
w546 <= not w328 and w545;
w547 <= not w405 and w546;
w548 <= not w207 and w547;
w549 <= not w275 and w548;
w550 <= not w86 and not w262;
w551 <= not w164 and w311;
w552 <= w45 and w204;
w553 <= not w106 and not w552;
w554 <= w59 and w109;
w555 <= w66 and w69;
w556 <= not w554 and not w555;
w557 <= not w110 and not w460;
w558 <= w97 and w134;
w559 <= not w70 and not w87;
w560 <= not w270 and w559;
w561 <= not w85 and w560;
w562 <= not w183 and w561;
w563 <= not w99 and w562;
w564 <= not w558 and w563;
w565 <= not w467 and w564;
w566 <= not w21 and w565;
w567 <= not w37 and not w177;
w568 <= w15 and w61;
w569 <= not w359 and not w568;
w570 <= not w89 and w569;
w571 <= not w335 and w570;
w572 <= w36 and w52;
w573 <= not w506 and not w572;
w574 <= w25 and w61;
w575 <= not w440 and not w574;
w576 <= w13 and w49;
w577 <= not w427 and not w576;
w578 <= w575 and w577;
w579 <= w573 and w578;
w580 <= w571 and w579;
w581 <= w567 and w580;
w582 <= w566 and w581;
w583 <= w557 and w582;
w584 <= w556 and w583;
w585 <= w553 and w584;
w586 <= not w333 and w585;
w587 <= not w84 and w586;
w588 <= not w158 and w587;
w589 <= not w58 and not w60;
w590 <= w15 and w48;
w591 <= w29 and w109;
w592 <= w48 and w134;
w593 <= not w387 and not w592;
w594 <= not w362 and w593;
w595 <= not w288 and w594;
w596 <= not w361 and w595;
w597 <= not w591 and w596;
w598 <= not w227 and w597;
w599 <= not w590 and w598;
w600 <= not w218 and not w502;
w601 <= w18 and w31;
w602 <= w88 and w97;
w603 <= not w216 and not w602;
w604 <= not w365 and w603;
w605 <= not w454 and w604;
w606 <= not w601 and w605;
w607 <= w41 and w95;
w608 <= w78 and w204;
w609 <= not w607 and not w608;
w610 <= not w79 and not w503;
w611 <= w609 and w610;
w612 <= w606 and w611;
w613 <= w600 and w612;
w614 <= w599 and w613;
w615 <= w589 and w614;
w616 <= w385 and w615;
w617 <= not w265 and w616;
w618 <= not w354 and w617;
w619 <= not w396 and w618;
w620 <= not w462 and w619;
w621 <= not w357 and w620;
w622 <= not w105 and w621;
w623 <= not w497 and w622;
w624 <= w48 and w78;
w625 <= not w125 and not w624;
w626 <= not w264 and not w274;
w627 <= not w355 and not w471;
w628 <= not w403 and w627;
w629 <= not w80 and not w189;
w630 <= w628 and w629;
w631 <= w626 and w630;
w632 <= w625 and w631;
w633 <= w623 and w632;
w634 <= w588 and w633;
w635 <= w551 and w634;
w636 <= w268 and w635;
w637 <= w550 and w636;
w638 <= w549 and w637;
w639 <= w535 and w638;
w640 <= w526 and w639;
w641 <= w137 and w640;
w642 <= w525 and w641;
w643 <= not w449 and w642;
w644 <= not w261 and w643;
w645 <= not w524 and w644;
w646 <= not w522 and not w645;
w647 <= w13 and w134;
w648 <= w57 and w69;
w649 <= w61 and w78;
w650 <= w25 and w66;
w651 <= w48 and w101;
w652 <= w72 and not w397;
w653 <= not w302 and w652;
w654 <= not w651 and w653;
w655 <= not w99 and not w186;
w656 <= not w90 and not w404;
w657 <= not w309 and w656;
w658 <= not w82 and not w395;
w659 <= w657 and w658;
w660 <= not w290 and w659;
w661 <= not w81 and w660;
w662 <= not w221 and w661;
w663 <= not w502 and w662;
w664 <= not w328 and w663;
w665 <= not w273 and w664;
w666 <= not w80 and not w506;
w667 <= not w306 and not w409;
w668 <= not w108 and not w454;
w669 <= not w93 and w668;
w670 <= not w471 and not w591;
w671 <= w669 and w670;
w672 <= w667 and w671;
w673 <= not w177 and w672;
w674 <= not w224 and w673;
w675 <= not w240 and w674;
w676 <= not w183 and w675;
w677 <= not w388 and w676;
w678 <= not w329 and w677;
w679 <= not w30 and w678;
w680 <= not w298 and w679;
w681 <= w36 and w45;
w682 <= not w141 and not w237;
w683 <= not w681 and w682;
w684 <= not w360 and w683;
w685 <= not w34 and w684;
w686 <= not w527 and w685;
w687 <= w59 and w88;
w688 <= not w89 and not w687;
w689 <= not w498 and w688;
w690 <= w128 and not w425;
w691 <= not w172 and w690;
w692 <= not w239 and w691;
w693 <= w689 and w692;
w694 <= w686 and w693;
w695 <= w680 and w694;
w696 <= w666 and w695;
w697 <= w665 and w696;
w698 <= w655 and w697;
w699 <= w654 and w698;
w700 <= w162 and w699;
w701 <= not w138 and w700;
w702 <= not w650 and w701;
w703 <= not w649 and w702;
w704 <= not w100 and w703;
w705 <= not w364 and w704;
w706 <= w15 and w23;
w707 <= not w386 and not w706;
w708 <= not w125 and not w175;
w709 <= not w293 and not w337;
w710 <= not w299 and not w362;
w711 <= not w213 and not w263;
w712 <= w20 and w25;
w713 <= not w272 and not w712;
w714 <= w711 and w713;
w715 <= w710 and w714;
w716 <= w709 and w715;
w717 <= w708 and w716;
w718 <= not w225 and w717;
w719 <= not w292 and w718;
w720 <= not w351 and w719;
w721 <= not w307 and w720;
w722 <= not w206 and w721;
w723 <= not w21 and not w428;
w724 <= not w405 and not w602;
w725 <= not w338 and not w448;
w726 <= w33 and w41;
w727 <= not w103 and not w726;
w728 <= not w96 and not w180;
w729 <= w727 and w728;
w730 <= w725 and w729;
w731 <= w724 and w730;
w732 <= w557 and w731;
w733 <= not w112 and w732;
w734 <= not w331 and w733;
w735 <= not w212 and w734;
w736 <= w723 and w735;
w737 <= not w384 and w736;
w738 <= w31 and w49;
w739 <= not w261 and not w446;
w740 <= not w430 and not w449;
w741 <= not w231 and not w427;
w742 <= not w357 and w741;
w743 <= not w310 and w742;
w744 <= w48 and w109;
w745 <= not w365 and not w744;
w746 <= not w85 and not w219;
w747 <= not w84 and not w352;
w748 <= not w558 and not w576;
w749 <= not w601 and w748;
w750 <= not w104 and not w555;
w751 <= not w607 and w750;
w752 <= w749 and w751;
w753 <= w747 and w752;
w754 <= w746 and w753;
w755 <= w745 and w754;
w756 <= not w163 and w755;
w757 <= not w178 and w756;
w758 <= not w301 and w757;
w759 <= not w497 and w758;
w760 <= w25 and w111;
w761 <= not w181 and not w355;
w762 <= not w230 and not w499;
w763 <= w761 and w762;
w764 <= not w56 and w763;
w765 <= not w760 and w764;
w766 <= not w439 and not w453;
w767 <= not w205 and w766;
w768 <= w402 and w767;
w769 <= w765 and w768;
w770 <= w759 and w769;
w771 <= w743 and w770;
w772 <= w740 and w771;
w773 <= w739 and w772;
w774 <= not w444 and w773;
w775 <= not w492 and w774;
w776 <= not w189 and w775;
w777 <= not w738 and w776;
w778 <= not w215 and w777;
w779 <= not w467 and w778;
w780 <= w55 and w589;
w781 <= not w124 and w780;
w782 <= w23 and w88;
w783 <= not w493 and not w782;
w784 <= not w158 and w783;
w785 <= not w552 and w784;
w786 <= not w288 and w785;
w787 <= w781 and w786;
w788 <= w779 and w787;
w789 <= w737 and w788;
w790 <= w722 and w789;
w791 <= w707 and w790;
w792 <= w705 and w791;
w793 <= not w648 and w792;
w794 <= not w86 and w793;
w795 <= not w234 and w794;
w796 <= not w574 and w795;
w797 <= not w431 and w796;
w798 <= not w77 and w797;
w799 <= not w403 and w798;
w800 <= not w647 and w799;
w801 <= not w424 and w800;
w802 <= not w123 and w801;
w803 <= not w645 and not w802;
w804 <= not w159 and not w178;
w805 <= not w90 and not w189;
w806 <= not w712 and w805;
w807 <= not w239 and w806;
w808 <= not w79 and not w648;
w809 <= not w171 and not w207;
w810 <= w15 and w31;
w811 <= not w236 and not w448;
w812 <= not w265 and not w650;
w813 <= w811 and w812;
w814 <= not w537 and w813;
w815 <= not w140 and w814;
w816 <= not w260 and w815;
w817 <= not w810 and w816;
w818 <= w13 and w18;
w819 <= w41 and w52;
w820 <= not w21 and not w231;
w821 <= w18 and w48;
w822 <= not w361 and not w497;
w823 <= not w261 and not w572;
w824 <= not w431 and w823;
w825 <= w822 and w824;
w826 <= not w529 and w825;
w827 <= not w354 and w826;
w828 <= not w352 and w827;
w829 <= not w821 and w828;
w830 <= not w364 and w829;
w831 <= not w360 and not w424;
w832 <= not w273 and not w362;
w833 <= not w289 and w654;
w834 <= not w328 and w833;
w835 <= w832 and w834;
w836 <= w786 and w835;
w837 <= w474 and w836;
w838 <= w63 and w837;
w839 <= w831 and w838;
w840 <= w334 and w839;
w841 <= w830 and w840;
w842 <= w442 and w841;
w843 <= w820 and w842;
w844 <= not w164 and w843;
w845 <= w507 and w844;
w846 <= not w554 and w845;
w847 <= not w819 and w846;
w848 <= not w760 and w847;
w849 <= not w266 and w848;
w850 <= not w818 and w849;
w851 <= not w363 and w850;
w852 <= not w177 and not w270;
w853 <= not w706 and w852;
w854 <= not w129 and not w524;
w855 <= not w65 and w854;
w856 <= not w568 and w855;
w857 <= w114 and w856;
w858 <= w853 and w857;
w859 <= not w190 and w858;
w860 <= not w124 and w859;
w861 <= not w263 and w860;
w862 <= not w744 and w861;
w863 <= not w396 and w862;
w864 <= not w330 and w863;
w865 <= not w80 and w864;
w866 <= not w186 and w865;
w867 <= w23 and w64;
w868 <= not w371 and not w867;
w869 <= w170 and w868;
w870 <= w389 and w869;
w871 <= not w77 and w870;
w872 <= not w54 and not w373;
w873 <= not w216 and w872;
w874 <= not w287 and w873;
w875 <= not w558 and w874;
w876 <= not w82 and not w230;
w877 <= w410 and w876;
w878 <= w875 and w877;
w879 <= w871 and w878;
w880 <= w866 and w879;
w881 <= w851 and w880;
w882 <= w817 and w881;
w883 <= w809 and w882;
w884 <= w808 and w883;
w885 <= w807 and w884;
w886 <= w358 and w885;
w887 <= w804 and w886;
w888 <= not w681 and w887;
w889 <= not w290 and w888;
w890 <= not w335 and w889;
w891 <= not w309 and w890;
w892 <= not w427 and w891;
w893 <= not w93 and w892;
w894 <= not w802 and not w893;
w895 <= not w46 and not w189;
w896 <= w29 and w33;
w897 <= not w332 and not w896;
w898 <= w895 and w897;
w899 <= not w287 and w898;
w900 <= not w819 and w899;
w901 <= not w37 and w900;
w902 <= not w175 and w901;
w903 <= not w16 and not w272;
w904 <= not w211 and w903;
w905 <= not w234 and w904;
w906 <= not w448 and w905;
w907 <= not w100 and w906;
w908 <= not w726 and w907;
w909 <= not w466 and w908;
w910 <= not w424 and w909;
w911 <= not w818 and w910;
w912 <= not w329 and not w364;
w913 <= not w261 and not w574;
w914 <= not w288 and not w555;
w915 <= w41 and w101;
w916 <= not w138 and not w221;
w917 <= not w301 and w916;
w918 <= w450 and w917;
w919 <= not w274 and w918;
w920 <= not w53 and w919;
w921 <= not w915 and w920;
w922 <= not w127 and w921;
w923 <= not w108 and w922;
w924 <= not w371 and not w524;
w925 <= not w401 and not w428;
w926 <= not w84 and not w552;
w927 <= not w760 and w926;
w928 <= w925 and w927;
w929 <= w924 and w928;
w930 <= w923 and w929;
w931 <= w445 and w930;
w932 <= w229 and w931;
w933 <= w173 and w932;
w934 <= w914 and w933;
w935 <= w913 and w934;
w936 <= w162 and w935;
w937 <= w353 and w936;
w938 <= not w681 and w937;
w939 <= not w112 and w938;
w940 <= not w624 and w939;
w941 <= not w99 and w940;
w942 <= not w273 and w941;
w943 <= not w60 and w942;
w944 <= not w85 and not w187;
w945 <= w66 and w95;
w946 <= w48 and w88;
w947 <= not w335 and not w607;
w948 <= not w362 and w947;
w949 <= not w946 and w948;
w950 <= not w370 and w949;
w951 <= not w867 and w950;
w952 <= not w65 and w951;
w953 <= not w558 and w952;
w954 <= not w945 and w953;
w955 <= not w499 and w954;
w956 <= not w125 and not w159;
w957 <= not w168 and w956;
w958 <= not w425 and w957;
w959 <= not w184 and w958;
w960 <= not w89 and not w208;
w961 <= w340 and w960;
w962 <= w959 and w961;
w963 <= w955 and w962;
w964 <= w366 and not w738;
w965 <= w963 and w964;
w966 <= w179 and w965;
w967 <= w944 and w966;
w968 <= w682 and w967;
w969 <= not w58 and w968;
w970 <= not w361 and w969;
w971 <= not w351 and w970;
w972 <= not w77 and w971;
w973 <= not w357 and w972;
w974 <= not w186 and w973;
w975 <= not w239 and not w492;
w976 <= w505 and w975;
w977 <= not w782 and w976;
w978 <= not w87 and w977;
w979 <= not w106 and w978;
w980 <= not w71 and w217;
w981 <= not w102 and not w181;
w982 <= not w98 and w981;
w983 <= w980 and w982;
w984 <= w979 and w983;
w985 <= w974 and w984;
w986 <= w943 and w985;
w987 <= w912 and w986;
w988 <= w557 and w987;
w989 <= w911 and w988;
w990 <= w902 and w989;
w991 <= w820 and w990;
w992 <= not w537 and w991;
w993 <= not w441 and w992;
w994 <= not w360 and w993;
w995 <= not w92 and w994;
w996 <= not w893 and not w995;
w997 <= w66 and w109;
w998 <= not w112 and not w351;
w999 <= not w354 and not w946;
w1000 <= not w272 and w999;
w1001 <= not w333 and w1000;
w1002 <= not w335 and w1001;
w1003 <= not w102 and w1002;
w1004 <= not w810 and w1003;
w1005 <= not w187 and not w444;
w1006 <= not w100 and not w172;
w1007 <= w45 and w59;
w1008 <= not w90 and not w1007;
w1009 <= w1006 and w1008;
w1010 <= w1005 and w1009;
w1011 <= not w236 and w1010;
w1012 <= not w576 and w1011;
w1013 <= not w84 and w1012;
w1014 <= not w42 and w1013;
w1015 <= not w108 and w1014;
w1016 <= not w124 and not w231;
w1017 <= not w472 and w1016;
w1018 <= not w357 and w1017;
w1019 <= not w386 and w1018;
w1020 <= not w209 and not w466;
w1021 <= w191 and w1020;
w1022 <= w1019 and w1021;
w1023 <= w1015 and w1022;
w1024 <= w1004 and w1023;
w1025 <= w998 and w1024;
w1026 <= w94 and w1025;
w1027 <= w505 and w1026;
w1028 <= not w50 and w1027;
w1029 <= not w997 and w1028;
w1030 <= not w233 and w1029;
w1031 <= not w524 and w1030;
w1032 <= not w301 and w1031;
w1033 <= not w275 and w1032;
w1034 <= not w306 and w1033;
w1035 <= not w206 and w1034;
w1036 <= w83 and w109;
w1037 <= w20 and w49;
w1038 <= not w401 and not w1037;
w1039 <= w57 and w134;
w1040 <= not w454 and not w1039;
w1041 <= not w538 and w1040;
w1042 <= not w706 and w1041;
w1043 <= not w106 and not w687;
w1044 <= not w647 and w1043;
w1045 <= w1042 and w1044;
w1046 <= w1038 and w1045;
w1047 <= not w71 and w1046;
w1048 <= not w332 and w1047;
w1049 <= not w397 and w1048;
w1050 <= not w782 and w1049;
w1051 <= not w1036 and w1050;
w1052 <= not w370 and w1051;
w1053 <= not w330 and w1052;
w1054 <= not w62 and w1053;
w1055 <= not w174 and not w181;
w1056 <= not w208 and w1055;
w1057 <= not w337 and w1056;
w1058 <= not w651 and w1057;
w1059 <= not w79 and w1058;
w1060 <= not w136 and w1059;
w1061 <= not w267 and w1060;
w1062 <= w61 and w95;
w1063 <= not w818 and not w1062;
w1064 <= not w363 and not w404;
w1065 <= not w86 and not w492;
w1066 <= not w441 and w1065;
w1067 <= not w359 and not w738;
w1068 <= not w56 and not w211;
w1069 <= not w425 and w1068;
w1070 <= not w601 and w1069;
w1071 <= not w234 and not w361;
w1072 <= not w608 and w1071;
w1073 <= not w329 and w1072;
w1074 <= not w140 and not w227;
w1075 <= not w499 and w1074;
w1076 <= not w205 and not w273;
w1077 <= not w210 and w1076;
w1078 <= not w98 and w1077;
w1079 <= w1075 and w1078;
w1080 <= w1073 and w1079;
w1081 <= w1070 and w1080;
w1082 <= w1067 and w1081;
w1083 <= w871 and w1082;
w1084 <= w1066 and w1083;
w1085 <= w1064 and w1084;
w1086 <= w589 and w1085;
w1087 <= w1063 and w1086;
w1088 <= not w572 and w1087;
w1089 <= not w302 and w1088;
w1090 <= not w239 and not w945;
w1091 <= w708 and w914;
w1092 <= not w67 and w1091;
w1093 <= not w590 and w1092;
w1094 <= not w34 and not w240;
w1095 <= not w228 and w1094;
w1096 <= not w126 and not w403;
w1097 <= not w216 and w1096;
w1098 <= not w649 and w1097;
w1099 <= w1095 and w1098;
w1100 <= w711 and w1099;
w1101 <= w1093 and w1100;
w1102 <= w1090 and w1101;
w1103 <= w1089 and w1102;
w1104 <= w1061 and w1103;
w1105 <= w1054 and w1104;
w1106 <= w600 and w1105;
w1107 <= w1035 and w1106;
w1108 <= w831 and w1107;
w1109 <= w872 and w1108;
w1110 <= not w552 and w1109;
w1111 <= not w430 and w1110;
w1112 <= not w395 and w1111;
w1113 <= not w497 and w1112;
w1114 <= not w995 and not w1113;
w1115 <= not w70 and not w592;
w1116 <= not w87 and not w440;
w1117 <= not w16 and not w264;
w1118 <= not w354 and not w370;
w1119 <= w173 and w872;
w1120 <= not w129 and w1119;
w1121 <= w610 and w1120;
w1122 <= w686 and w1121;
w1123 <= w1090 and w1122;
w1124 <= w722 and w1123;
w1125 <= w1118 and w1124;
w1126 <= w1117 and w1125;
w1127 <= not w236 and w1126;
w1128 <= not w71 and w1127;
w1129 <= not w46 and w1128;
w1130 <= not w289 and w1129;
w1131 <= not w159 and w1130;
w1132 <= not w819 and w1131;
w1133 <= not w108 and w1132;
w1134 <= not w99 and w1133;
w1135 <= not w471 and w1134;
w1136 <= not w538 and w1135;
w1137 <= not w590 and w1136;
w1138 <= w57 and w64;
w1139 <= not w504 and not w915;
w1140 <= not w275 and not w462;
w1141 <= not w810 and w1140;
w1142 <= w1139 and w1141;
w1143 <= not w262 and w1142;
w1144 <= not w163 and w1143;
w1145 <= not w1138 and w1144;
w1146 <= not w260 and w1145;
w1147 <= not w89 and not w189;
w1148 <= not w335 and w1147;
w1149 <= not w37 and w1148;
w1150 <= not w266 and w1149;
w1151 <= not w524 and w1150;
w1152 <= not w102 and not w498;
w1153 <= not w241 and w1152;
w1154 <= not w186 and w1153;
w1155 <= not w357 and not w591;
w1156 <= not w157 and w1155;
w1157 <= w917 and w1156;
w1158 <= w1154 and w1157;
w1159 <= w1151 and w1158;
w1160 <= w1089 and w1159;
w1161 <= w737 and w1160;
w1162 <= w1146 and w1161;
w1163 <= w1137 and w1162;
w1164 <= w1116 and w1163;
w1165 <= w1115 and w1164;
w1166 <= not w453 and w1165;
w1167 <= not w309 and w1166;
w1168 <= not w536 and w1167;
w1169 <= not w135 and w1168;
w1170 <= not w230 and w1169;
w1171 <= not w1113 and not w1170;
w1172 <= not w159 and not w332;
w1173 <= not w85 and not w352;
w1174 <= not w240 and w1173;
w1175 <= not w309 and w1174;
w1176 <= w525 and w1175;
w1177 <= not w337 and w1176;
w1178 <= not w431 and w1177;
w1179 <= not w359 and w1178;
w1180 <= not w212 and w1179;
w1181 <= w88 and w204;
w1182 <= not w209 and not w404;
w1183 <= not w287 and not w1036;
w1184 <= not w127 and not w186;
w1185 <= w238 and w1184;
w1186 <= not w608 and w1185;
w1187 <= not w306 and not w439;
w1188 <= not w303 and not w706;
w1189 <= not w190 and not w497;
w1190 <= not w34 and not w184;
w1191 <= w749 and w1190;
w1192 <= w669 and w1191;
w1193 <= w1189 and w1192;
w1194 <= w1188 and w1193;
w1195 <= w1187 and w1194;
w1196 <= not w430 and w1195;
w1197 <= not w231 and w1196;
w1198 <= not w896 and w1197;
w1199 <= not w502 and w1198;
w1200 <= w179 and not w915;
w1201 <= not w472 and w1200;
w1202 <= not w105 and w1201;
w1203 <= not w21 and w1202;
w1204 <= not w362 and not w384;
w1205 <= not w264 and w1204;
w1206 <= not w819 and w1205;
w1207 <= not w89 and not w449;
w1208 <= w468 and not w552;
w1209 <= not w333 and w1208;
w1210 <= w1207 and w1209;
w1211 <= w1206 and w1210;
w1212 <= w1038 and w1211;
w1213 <= w1203 and w1212;
w1214 <= w1199 and w1213;
w1215 <= w1186 and w1214;
w1216 <= w170 and w1215;
w1217 <= w220 and w1216;
w1218 <= w1183 and w1217;
w1219 <= w1182 and w1218;
w1220 <= not w1181 and w1219;
w1221 <= not w361 and w1220;
w1222 <= not w124 and w1221;
w1223 <= not w395 and w1222;
w1224 <= not w222 and w1223;
w1225 <= not w867 and w1224;
w1226 <= not w504 and w1225;
w1227 <= not w493 and not w738;
w1228 <= not w310 and not w574;
w1229 <= not w208 and w1228;
w1230 <= w670 and w1229;
w1231 <= w294 and w1230;
w1232 <= not w444 and w1231;
w1233 <= not w125 and w1232;
w1234 <= not w396 and w1233;
w1235 <= not w536 and w1234;
w1236 <= not w126 and w1235;
w1237 <= not w371 and w1236;
w1238 <= not w60 and w1237;
w1239 <= not w16 and w1238;
w1240 <= not w568 and w1239;
w1241 <= w13 and w45;
w1242 <= not w330 and not w624;
w1243 <= not w388 and w1242;
w1244 <= not w1241 and w1243;
w1245 <= not w554 and w1244;
w1246 <= not w225 and w1245;
w1247 <= not w266 and w1246;
w1248 <= not w205 and w1247;
w1249 <= not w329 and not w331;
w1250 <= not w386 and w1249;
w1251 <= w1074 and w1250;
w1252 <= not w265 and w1251;
w1253 <= not w274 and w1252;
w1254 <= not w81 and w1253;
w1255 <= not w427 and w1254;
w1256 <= not w649 and w1255;
w1257 <= not w239 and w1256;
w1258 <= not w272 and w1257;
w1259 <= not w453 and not w503;
w1260 <= not w92 and w1259;
w1261 <= not w405 and w1260;
w1262 <= not w592 and w1261;
w1263 <= not w363 and w1262;
w1264 <= not w84 and not w537;
w1265 <= not w782 and not w821;
w1266 <= not w172 and w1265;
w1267 <= not w135 and not w234;
w1268 <= not w96 and w1267;
w1269 <= w1266 and w1268;
w1270 <= w1264 and w1269;
w1271 <= w1263 and w1270;
w1272 <= w1258 and w1271;
w1273 <= w666 and w1272;
w1274 <= w1248 and w1273;
w1275 <= not w681 and w1274;
w1276 <= not w216 and w1275;
w1277 <= not w270 and w1276;
w1278 <= not w50 and w1277;
w1279 <= not w174 and w1278;
w1280 <= not w161 and w1279;
w1281 <= not w53 and not w289;
w1282 <= not w302 and not w335;
w1283 <= w1281 and w1282;
w1284 <= w765 and w1283;
w1285 <= w1280 and w1284;
w1286 <= w1240 and w1285;
w1287 <= w1227 and w1286;
w1288 <= w1226 and w1287;
w1289 <= w1180 and w1288;
w1290 <= w872 and w1289;
w1291 <= w1172 and w1290;
w1292 <= not w129 and w1291;
w1293 <= not w263 and w1292;
w1294 <= not w110 and w1293;
w1295 <= not w572 and w1294;
w1296 <= not w357 and w1295;
w1297 <= not w403 and w1296;
w1298 <= not w466 and w1297;
w1299 <= not w301 and w1298;
w1300 <= not w1170 and not w1299;
w1301 <= not w160 and not w536;
w1302 <= not w105 and not w208;
w1303 <= not w126 and not w287;
w1304 <= not w207 and w1303;
w1305 <= not w240 and not w441;
w1306 <= not w181 and w1305;
w1307 <= not w647 and w1306;
w1308 <= w1304 and w1307;
w1309 <= w1302 and w1308;
w1310 <= not w46 and w1309;
w1311 <= not w82 and w1310;
w1312 <= not w819 and w1311;
w1313 <= not w237 and w1312;
w1314 <= not w466 and not w1241;
w1315 <= not w264 and not w409;
w1316 <= not w164 and w1315;
w1317 <= not w289 and w1316;
w1318 <= not w231 and w1317;
w1319 <= not w524 and w1318;
w1320 <= not w265 and not w738;
w1321 <= not w726 and w1320;
w1322 <= not w307 and w1321;
w1323 <= not w266 and not w867;
w1324 <= not w138 and not w396;
w1325 <= not w555 and w1324;
w1326 <= not w454 and w1325;
w1327 <= not w210 and not w310;
w1328 <= not w338 and not w1037;
w1329 <= not w135 and w1328;
w1330 <= w1327 and w1329;
w1331 <= w781 and w1330;
w1332 <= w1326 and w1331;
w1333 <= w1323 and w1332;
w1334 <= w1322 and w1333;
w1335 <= w1319 and w1334;
w1336 <= w1314 and w1335;
w1337 <= w1115 and w1336;
w1338 <= w1063 and w1337;
w1339 <= not w397 and w1338;
w1340 <= not w167 and w1339;
w1341 <= not w158 and w1340;
w1342 <= not w558 and w1341;
w1343 <= not w42 and not w650;
w1344 <= not w568 and not w896;
w1345 <= w1343 and w1344;
w1346 <= w724 and w1345;
w1347 <= not w687 and w1346;
w1348 <= not w213 and w1347;
w1349 <= not w261 and w1348;
w1350 <= not w425 and w1349;
w1351 <= not w80 and w1350;
w1352 <= not w34 and w1351;
w1353 <= not w607 and w1352;
w1354 <= not w206 and w1353;
w1355 <= not w302 and not w431;
w1356 <= not w608 and w1355;
w1357 <= not w21 and w1356;
w1358 <= not w26 and not w99;
w1359 <= not w100 and not w430;
w1360 <= not w554 and not w706;
w1361 <= not w211 and not w527;
w1362 <= not w624 and w1361;
w1363 <= not w364 and w1362;
w1364 <= w1360 and w1363;
w1365 <= w1154 and w1364;
w1366 <= w1359 and w1365;
w1367 <= w998 and w1366;
w1368 <= not w462 and w1367;
w1369 <= not w37 and w1368;
w1370 <= not w166 and w1369;
w1371 <= not w330 and not w506;
w1372 <= not w760 and w1371;
w1373 <= not w224 and not w997;
w1374 <= not w537 and not w576;
w1375 <= not w85 and w1374;
w1376 <= w1000 and w1375;
w1377 <= w1373 and w1376;
w1378 <= w1372 and w1377;
w1379 <= w539 and w1378;
w1380 <= w1370 and w1379;
w1381 <= w1074 and w1380;
w1382 <= w831 and w1381;
w1383 <= w762 and w1382;
w1384 <= w1172 and w1383;
w1385 <= not w782 and w1384;
w1386 <= not w352 and w1385;
w1387 <= not w163 and w1386;
w1388 <= not w108 and w1387;
w1389 <= not w30 and w1388;
w1390 <= w389 and w1389;
w1391 <= not w574 and w1390;
w1392 <= not w87 and not w502;
w1393 <= not w96 and w1392;
w1394 <= w1391 and w1393;
w1395 <= w1358 and w1394;
w1396 <= w1357 and w1395;
w1397 <= w1354 and w1396;
w1398 <= w1342 and w1397;
w1399 <= w1313 and w1398;
w1400 <= w1301 and w1399;
w1401 <= w1204 and w1400;
w1402 <= not w493 and w1401;
w1403 <= not w444 and w1402;
w1404 <= not w84 and w1403;
w1405 <= not w337 and w1404;
w1406 <= not w712 and w1405;
w1407 <= not w67 and w1406;
w1408 <= not w1299 and not w1407;
w1409 <= not w362 and not w503;
w1410 <= not w218 and w1409;
w1411 <= not w167 and not w267;
w1412 <= not w330 and not w351;
w1413 <= not w309 and w1412;
w1414 <= not w431 and not w681;
w1415 <= not w184 and not w590;
w1416 <= w188 and w1319;
w1417 <= not w219 and w1416;
w1418 <= not w650 and w1417;
w1419 <= not w329 and w1418;
w1420 <= not w67 and w1419;
w1421 <= not w405 and w1420;
w1422 <= not w945 and w1421;
w1423 <= not w93 and w1422;
w1424 <= not w42 and not w946;
w1425 <= not w105 and w1424;
w1426 <= not w370 and w1425;
w1427 <= not w819 and w1426;
w1428 <= not w266 and w1427;
w1429 <= not w92 and w1428;
w1430 <= not w230 and w1429;
w1431 <= not w62 and w1430;
w1432 <= not w90 and not w744;
w1433 <= not w448 and not w687;
w1434 <= not w360 and w1433;
w1435 <= w1432 and w1434;
w1436 <= w1431 and w1435;
w1437 <= w1423 and w1436;
w1438 <= w1415 and w1437;
w1439 <= w1414 and w1438;
w1440 <= w1413 and w1439;
w1441 <= not w537 and w1440;
w1442 <= not w269 and w1441;
w1443 <= not w108 and w1442;
w1444 <= not w592 and w1443;
w1445 <= not w504 and w1444;
w1446 <= not w205 and w1445;
w1447 <= not w299 and w895;
w1448 <= not w58 and w1447;
w1449 <= not w648 and w1448;
w1450 <= not w262 and w1449;
w1451 <= not w112 and w1450;
w1452 <= not w210 and w1451;
w1453 <= not w760 and w1452;
w1454 <= not w175 and w1453;
w1455 <= not w207 and w1454;
w1456 <= not w706 and w1455;
w1457 <= not w158 and not w497;
w1458 <= not w84 and not w233;
w1459 <= not w81 and not w430;
w1460 <= not w102 and w1459;
w1461 <= not w538 and w1460;
w1462 <= not w424 and w1461;
w1463 <= not w288 and not w331;
w1464 <= not w261 and w1463;
w1465 <= not w384 and w1464;
w1466 <= not w228 and not w601;
w1467 <= w1064 and w1466;
w1468 <= not w651 and w1467;
w1469 <= w1266 and w1468;
w1470 <= w1465 and w1469;
w1471 <= w658 and w1470;
w1472 <= w374 and w1471;
w1473 <= w1462 and w1472;
w1474 <= w1040 and w1473;
w1475 <= w1240 and w1474;
w1476 <= w1458 and w1475;
w1477 <= w1361 and w1476;
w1478 <= w525 and w1477;
w1479 <= w1457 and w1478;
w1480 <= not w274 and w1479;
w1481 <= not w440 and w1480;
w1482 <= not w241 and w1481;
w1483 <= not w239 and w1482;
w1484 <= not w460 and w1483;
w1485 <= not w209 and not w493;
w1486 <= w137 and w217;
w1487 <= w1485 and w1486;
w1488 <= not w915 and w1487;
w1489 <= not w388 and w1488;
w1490 <= not w212 and w1489;
w1491 <= not w65 and not w301;
w1492 <= not w206 and not w397;
w1493 <= w1491 and w1492;
w1494 <= w1490 and w1493;
w1495 <= w1484 and w1494;
w1496 <= w1456 and w1495;
w1497 <= w566 and w1496;
w1498 <= w1446 and w1497;
w1499 <= w1411 and w1498;
w1500 <= w1410 and w1499;
w1501 <= w223 and w1500;
w1502 <= w1314 and w1501;
w1503 <= not w359 and w1502;
w1504 <= not w140 and w1503;
w1505 <= not w472 and w1504;
w1506 <= not w96 and w1505;
w1507 <= not w364 and w1506;
w1508 <= not w1407 and not w1507;
w1509 <= not w219 and not w467;
w1510 <= not w105 and not w263;
w1511 <= not w77 and not w649;
w1512 <= not w207 and not w1138;
w1513 <= not w387 and w707;
w1514 <= w1512 and w1513;
w1515 <= w1116 and w1514;
w1516 <= w808 and w1515;
w1517 <= w170 and w1516;
w1518 <= not w552 and w1517;
w1519 <= not w210 and w1518;
w1520 <= not w21 and w1519;
w1521 <= not w574 and not w592;
w1522 <= not w209 and not w439;
w1523 <= not w136 and w1522;
w1524 <= w1363 and w1523;
w1525 <= w1521 and w1524;
w1526 <= w1520 and w1525;
w1527 <= w1415 and w1526;
w1528 <= w55 and w1527;
w1529 <= w1511 and w1528;
w1530 <= w666 and w1529;
w1531 <= w91 and w1530;
w1532 <= not w189 and w1531;
w1533 <= not w576 and w1532;
w1534 <= not w106 and w1533;
w1535 <= not w222 and w1534;
w1536 <= not w112 and not w171;
w1537 <= not w96 and not w289;
w1538 <= not w125 and not w215;
w1539 <= not w538 and not w946;
w1540 <= w1538 and w1539;
w1541 <= w229 and w1540;
w1542 <= not w335 and w1541;
w1543 <= not w37 and w1542;
w1544 <= not w431 and w1543;
w1545 <= not w181 and w1544;
w1546 <= not w427 and not w945;
w1547 <= not w1181 and w1546;
w1548 <= not w262 and w1547;
w1549 <= not w572 and w1548;
w1550 <= not w373 and w1549;
w1551 <= not w46 and not w536;
w1552 <= not w607 and w1551;
w1553 <= not w264 and not w555;
w1554 <= not w915 and w1553;
w1555 <= not w272 and w1554;
w1556 <= not w384 and w1555;
w1557 <= w1552 and w1556;
w1558 <= w1550 and w1557;
w1559 <= w1545 and w1558;
w1560 <= w1537 and w1559;
w1561 <= not w236 and w1560;
w1562 <= not w493 and w1561;
w1563 <= not w396 and w1562;
w1564 <= not w26 and w1563;
w1565 <= not w351 and w1564;
w1566 <= not w303 and w1565;
w1567 <= not w403 and w1566;
w1568 <= not w558 and w1567;
w1569 <= not w212 and w1568;
w1570 <= not w424 and w1569;
w1571 <= not w359 and not w1241;
w1572 <= not w213 and w1571;
w1573 <= not w554 and w1572;
w1574 <= not w309 and w1573;
w1575 <= not w186 and w1574;
w1576 <= not w274 and not w362;
w1577 <= not w208 and w1576;
w1578 <= not w647 and w1577;
w1579 <= not w163 and not w712;
w1580 <= not w158 and w1189;
w1581 <= not w266 and w1580;
w1582 <= w1579 and w1581;
w1583 <= w1578 and w1582;
w1584 <= w1575 and w1583;
w1585 <= w1570 and w1584;
w1586 <= w1536 and w1585;
w1587 <= w1535 and w1586;
w1588 <= w1510 and w1587;
w1589 <= w358 and w1588;
w1590 <= w680 and w1589;
w1591 <= w1183 and w1590;
w1592 <= w1509 and w1591;
w1593 <= w294 and w1592;
w1594 <= not w86 and w1593;
w1595 <= not w261 and w1594;
w1596 <= not w503 and w1595;
w1597 <= not w221 and w1596;
w1598 <= not w502 and w1597;
w1599 <= not w1039 and w1598;
w1600 <= not w206 and w1599;
w1601 <= not w1507 and not w1600;
w1602 <= not w67 and not w184;
w1603 <= not w26 and not w397;
w1604 <= not w363 and w723;
w1605 <= w784 and w1604;
w1606 <= w868 and w1605;
w1607 <= w1410 and w1606;
w1608 <= w1603 and w1607;
w1609 <= not w46 and w1608;
w1610 <= not w651 and w1609;
w1611 <= not w360 and w1610;
w1612 <= not w524 and w1611;
w1613 <= not w466 and w1612;
w1614 <= not w166 and w1613;
w1615 <= not w649 and not w1039;
w1616 <= not w568 and w1615;
w1617 <= w238 and w1616;
w1618 <= w725 and w1617;
w1619 <= not w299 and w1618;
w1620 <= not w529 and w1619;
w1621 <= not w370 and w1620;
w1622 <= not w225 and w1621;
w1623 <= not w104 and not w124;
w1624 <= not w330 and w1623;
w1625 <= not w536 and w1624;
w1626 <= not w328 and w1625;
w1627 <= not w364 and not w453;
w1628 <= not w71 and not w234;
w1629 <= not w183 and w1628;
w1630 <= not w409 and w1629;
w1631 <= not w90 and not w303;
w1632 <= not w298 and w1631;
w1633 <= w1630 and w1632;
w1634 <= w713 and w1633;
w1635 <= w1627 and w1634;
w1636 <= w1626 and w1635;
w1637 <= w1622 and w1636;
w1638 <= w1614 and w1637;
w1639 <= w1602 and w1638;
w1640 <= not w103 and w1639;
w1641 <= not w222 and w1640;
w1642 <= not w307 and w1641;
w1643 <= not w275 and w1642;
w1644 <= not w401 and not w471;
w1645 <= w1264 and w1644;
w1646 <= w1643 and w1645;
w1647 <= w1096 and w1646;
w1648 <= not w87 and w1647;
w1649 <= not w224 and w1648;
w1650 <= not w81 and w1649;
w1651 <= not w650 and w1650;
w1652 <= not w141 and w1651;
w1653 <= not w180 and w1652;
w1654 <= not w93 and w1653;
w1655 <= not w135 and not w387;
w1656 <= not w454 and w1655;
w1657 <= w1229 and w1656;
w1658 <= not w58 and w1657;
w1659 <= not w1181 and w1658;
w1660 <= not w290 and w1659;
w1661 <= not w110 and not w163;
w1662 <= not w30 and not w601;
w1663 <= not w129 and w1662;
w1664 <= not w365 and w1663;
w1665 <= not w209 and w1664;
w1666 <= not w424 and w1665;
w1667 <= not w288 and not w1007;
w1668 <= not w332 and w1667;
w1669 <= not w98 and w1668;
w1670 <= not w384 and w1669;
w1671 <= not w425 and w1538;
w1672 <= not w186 and w1671;
w1673 <= not w178 and not w572;
w1674 <= not w42 and not w818;
w1675 <= not w54 and not w430;
w1676 <= w1674 and w1675;
w1677 <= w1673 and w1676;
w1678 <= w1672 and w1677;
w1679 <= w1307 and w1678;
w1680 <= w1670 and w1679;
w1681 <= w1666 and w1680;
w1682 <= w1661 and w1681;
w1683 <= w162 and w1682;
w1684 <= not w265 and w1683;
w1685 <= not w361 and w1684;
w1686 <= not w106 and w1685;
w1687 <= not w1036 and w1686;
w1688 <= not w112 and w1687;
w1689 <= not w502 and w1688;
w1690 <= not w168 and not w687;
w1691 <= not w79 and w1690;
w1692 <= not w726 and w1691;
w1693 <= not w607 and w1692;
w1694 <= not w590 and w1693;
w1695 <= not w167 and not w213;
w1696 <= not w359 and not w624;
w1697 <= not w404 and w1696;
w1698 <= not w159 and w1697;
w1699 <= w1695 and w1698;
w1700 <= w629 and w1699;
w1701 <= w1694 and w1700;
w1702 <= w1689 and w1701;
w1703 <= w709 and w1702;
w1704 <= w1660 and w1703;
w1705 <= w1654 and w1704;
w1706 <= w1117 and w1705;
w1707 <= w525 and w1706;
w1708 <= not w70 and w1707;
w1709 <= not w335 and w1708;
w1710 <= not w498 and w1709;
w1711 <= not w439 and w1710;
w1712 <= not w99 and w1711;
w1713 <= not w260 and w1712;
w1714 <= not w810 and w1713;
w1715 <= not w1600 and not w1714;
w1716 <= not w590 and not w760;
w1717 <= not w124 and not w527;
w1718 <= not w89 and not w234;
w1719 <= not w1037 and w1718;
w1720 <= not w98 and not w1138;
w1721 <= w1719 and w1720;
w1722 <= w831 and w1721;
w1723 <= w1717 and w1722;
w1724 <= not w441 and w1723;
w1725 <= w1690 and w1724;
w1726 <= not w395 and w1725;
w1727 <= not w462 and w1726;
w1728 <= not w266 and w1727;
w1729 <= not w624 and w1728;
w1730 <= not w287 and not w449;
w1731 <= not w158 and w1730;
w1732 <= not w448 and w1731;
w1733 <= not w298 and w1732;
w1734 <= not w270 and not w554;
w1735 <= not w373 and w1734;
w1736 <= w1343 and w1735;
w1737 <= w429 and w1736;
w1738 <= w1733 and w1737;
w1739 <= w955 and w1738;
w1740 <= w450 and w1739;
w1741 <= w128 and w1740;
w1742 <= not w71 and w1741;
w1743 <= not w106 and w1742;
w1744 <= not w352 and w1743;
w1745 <= not w231 and w1744;
w1746 <= not w209 and w1745;
w1747 <= not w307 and w1746;
w1748 <= not w821 and w1747;
w1749 <= not w123 and w1748;
w1750 <= not w404 and not w576;
w1751 <= not w138 and w1750;
w1752 <= not w240 and w1751;
w1753 <= not w206 and w1752;
w1754 <= not w810 and w1753;
w1755 <= w389 and w443;
w1756 <= not w498 and w1755;
w1757 <= not w1039 and w1756;
w1758 <= not w30 and w1757;
w1759 <= not w60 and not w93;
w1760 <= not w338 and not w537;
w1761 <= not w166 and not w439;
w1762 <= not w401 and not w712;
w1763 <= not w161 and not w1036;
w1764 <= w1602 and w1763;
w1765 <= w1762 and w1764;
w1766 <= w526 and w1765;
w1767 <= not w997 and w1766;
w1768 <= not w225 and w1767;
w1769 <= not w440 and w1768;
w1770 <= not w466 and w1769;
w1771 <= not w306 and w1770;
w1772 <= not w504 and w1771;
w1773 <= not w272 and w1772;
w1774 <= not w56 and not w471;
w1775 <= w897 and w1774;
w1776 <= not w290 and w1775;
w1777 <= not w85 and w1776;
w1778 <= not w354 and w1777;
w1779 <= not w538 and w1778;
w1780 <= w1773 and w1779;
w1781 <= w1761 and w1780;
w1782 <= w455 and w1781;
w1783 <= w1511 and w1782;
w1784 <= w761 and w1783;
w1785 <= w1760 and w1784;
w1786 <= w1759 and w1785;
w1787 <= not w782 and w1786;
w1788 <= not w264 and w1787;
w1789 <= not w738 and w1788;
w1790 <= not w506 and w1789;
w1791 <= not w430 and w1790;
w1792 <= not w135 and w1791;
w1793 <= not w574 and w1792;
w1794 <= not w427 and w1793;
w1795 <= not w164 and not w302;
w1796 <= not w409 and w1795;
w1797 <= w1794 and w1796;
w1798 <= w711 and w1797;
w1799 <= w1758 and w1798;
w1800 <= w1754 and w1799;
w1801 <= w1749 and w1800;
w1802 <= w1729 and w1801;
w1803 <= w1466 and w1802;
w1804 <= w1716 and w1803;
w1805 <= w468 and w1804;
w1806 <= w217 and w1805;
w1807 <= w334 and w1806;
w1808 <= w975 and w1807;
w1809 <= not w87 and w1808;
w1810 <= not w174 and w1809;
w1811 <= not w222 and w1810;
w1812 <= not w186 and w1811;
w1813 <= not w1714 and not w1812;
w1814 <= not w100 and not w387;
w1815 <= w1373 and w1814;
w1816 <= w1182 and w1815;
w1817 <= not w333 and w1816;
w1818 <= not w34 and w1817;
w1819 <= not w647 and w1818;
w1820 <= not w213 and not w744;
w1821 <= not w819 and w1820;
w1822 <= not w180 and w1821;
w1823 <= not w712 and w1822;
w1824 <= not w218 and w1823;
w1825 <= not w62 and w1824;
w1826 <= not w71 and not w222;
w1827 <= not w233 and w1826;
w1828 <= not w136 and w1827;
w1829 <= not w215 and not w602;
w1830 <= w553 and w1829;
w1831 <= not w82 and w1830;
w1832 <= not w93 and not w446;
w1833 <= not w228 and w1832;
w1834 <= w1831 and w1833;
w1835 <= w1632 and w1834;
w1836 <= w1280 and w1835;
w1837 <= w1146 and w1836;
w1838 <= w974 and w1837;
w1839 <= w1536 and w1838;
w1840 <= w1411 and w1839;
w1841 <= w1828 and w1840;
w1842 <= w1825 and w1841;
w1843 <= w1819 and w1842;
w1844 <= not w1037 and w1843;
w1845 <= not w529 and w1844;
w1846 <= not w354 and w1845;
w1847 <= not w650 and w1846;
w1848 <= not w527 and w1847;
w1849 <= not w1812 and not w1848;
w1850 <= not w159 and not w466;
w1851 <= not w174 and not w462;
w1852 <= not w506 and not w558;
w1853 <= not w648 and not w1007;
w1854 <= not w264 and w1853;
w1855 <= not w744 and w1854;
w1856 <= not w237 and w1855;
w1857 <= not w651 and w1856;
w1858 <= not w67 and w1857;
w1859 <= not w187 and w1858;
w1860 <= not w239 and w1859;
w1861 <= not w167 and not w687;
w1862 <= not w1037 and w1861;
w1863 <= not w608 and w1862;
w1864 <= w179 and not w361;
w1865 <= not w396 and w1864;
w1866 <= not w307 and w1865;
w1867 <= w1492 and w1866;
w1868 <= w809 and w1867;
w1869 <= w1361 and w1868;
w1870 <= not w576 and w1869;
w1871 <= not w449 and w1870;
w1872 <= not w274 and w1871;
w1873 <= not w208 and w1872;
w1874 <= not w212 and w1873;
w1875 <= not w260 and w1874;
w1876 <= not w236 and not w819;
w1877 <= not w309 and w1876;
w1878 <= not w65 and not w234;
w1879 <= not w1039 and w1878;
w1880 <= w924 and w1879;
w1881 <= w1877 and w1880;
w1882 <= w1875 and w1881;
w1883 <= w1863 and w1882;
w1884 <= w912 and w1883;
w1885 <= w473 and w1884;
w1886 <= not w53 and w1885;
w1887 <= not w175 and w1886;
w1888 <= not w218 and w1887;
w1889 <= not w726 and w1888;
w1890 <= not w1138 and w1889;
w1891 <= not w945 and w1890;
w1892 <= not w16 and w1891;
w1893 <= not w157 and w1892;
w1894 <= not w404 and not w574;
w1895 <= not w54 and w1894;
w1896 <= w707 and w1895;
w1897 <= w447 and w1896;
w1898 <= w1118 and w1897;
w1899 <= w831 and w1898;
w1900 <= not w552 and w1899;
w1901 <= not w302 and w1900;
w1902 <= not w330 and w1901;
w1903 <= not w460 and w1902;
w1904 <= not w293 and w1903;
w1905 <= not w56 and w156;
w1906 <= not w428 and w1905;
w1907 <= w353 and w1183;
w1908 <= not w30 and w1907;
w1909 <= w1906 and w1908;
w1910 <= w593 and w1909;
w1911 <= w812 and w1910;
w1912 <= w1904 and w1911;
w1913 <= w1893 and w1912;
w1914 <= w1860 and w1913;
w1915 <= w1852 and w1914;
w1916 <= w1851 and w1915;
w1917 <= w1850 and w1916;
w1918 <= w450 and w1917;
w1919 <= w1509 and w1918;
w1920 <= not w493 and w1919;
w1921 <= not w215 and w1920;
w1922 <= not w351 and w1921;
w1923 <= not w231 and w1922;
w1924 <= not w440 and w1923;
w1925 <= not w359 and w1924;
w1926 <= not w228 and w1925;
w1927 <= not w205 and w1926;
w1928 <= not w1848 and not w1927;
w1929 <= not w237 and not w1037;
w1930 <= not w103 and not w332;
w1931 <= not w524 and w1930;
w1932 <= w1833 and w1931;
w1933 <= w728 and w1932;
w1934 <= w232 and w1933;
w1935 <= w1929 and w1934;
w1936 <= not w1036 and w1935;
w1937 <= not w140 and w1936;
w1938 <= not w126 and w1937;
w1939 <= not w1062 and w1938;
w1940 <= not w424 and w1939;
w1941 <= not w810 and w1940;
w1942 <= not w427 and not w472;
w1943 <= not w602 and w1942;
w1944 <= not w395 and w1943;
w1945 <= not w65 and w1944;
w1946 <= w271 and w914;
w1947 <= not w307 and w1946;
w1948 <= not w275 and not w946;
w1949 <= not w100 and not w175;
w1950 <= w1948 and w1949;
w1951 <= w1040 and w1950;
w1952 <= not w388 and w1951;
w1953 <= not w290 and not w444;
w1954 <= not w82 and w1953;
w1955 <= not w306 and w1954;
w1956 <= not w98 and not w651;
w1957 <= not w30 and not w681;
w1958 <= not w141 and not w299;
w1959 <= not w357 and w1958;
w1960 <= not w301 and w1959;
w1961 <= not w157 and not w373;
w1962 <= w1264 and w1961;
w1963 <= w464 and w1962;
w1964 <= w1960 and w1963;
w1965 <= w1626 and w1964;
w1966 <= w1957 and w1965;
w1967 <= w1956 and w1966;
w1968 <= w1265 and w1967;
w1969 <= w1603 and w1968;
w1970 <= w944 and w1969;
w1971 <= not w554 and w1970;
w1972 <= not w127 and w1971;
w1973 <= not w403 and w1972;
w1974 <= not w371 and w1973;
w1975 <= not w504 and w1974;
w1976 <= w1955 and w1975;
w1977 <= w1952 and w1976;
w1978 <= w1535 and w1977;
w1979 <= w1947 and w1978;
w1980 <= w1118 and w1979;
w1981 <= w1945 and w1980;
w1982 <= w1941 and w1981;
w1983 <= w655 and w1982;
w1984 <= not w493 and w1983;
w1985 <= not w219 and w1984;
w1986 <= not w138 and w1985;
w1987 <= w1730 and w1986;
w1988 <= not w225 and w1987;
w1989 <= not w37 and w1988;
w1990 <= not w359 and w1989;
w1991 <= not w405 and w1990;
w1992 <= not w497 and w1991;
w1993 <= not w1927 and not w1992;
w1994 <= not w87 and not w125;
w1995 <= w670 and w1994;
w1996 <= w526 and w1995;
w1997 <= not w167 and w1996;
w1998 <= not w744 and w1997;
w1999 <= not w431 and w1998;
w2000 <= not w79 and w1999;
w2001 <= not w233 and w2000;
w2002 <= not w272 and w2001;
w2003 <= not w568 and w2002;
w2004 <= w1183 and w1187;
w2005 <= not w224 and w2004;
w2006 <= not w190 and w2005;
w2007 <= not w424 and w2006;
w2008 <= not w104 and not w572;
w2009 <= not w183 and w2008;
w2010 <= not w1039 and w2009;
w2011 <= w1719 and w2010;
w2012 <= w747 and w2011;
w2013 <= w1067 and w2012;
w2014 <= w142 and w2013;
w2015 <= w1020 and w2014;
w2016 <= w853 and w2015;
w2017 <= w2007 and w2016;
w2018 <= w2003 and w2017;
w2019 <= w450 and w2018;
w2020 <= not w492 and w2019;
w2021 <= not w354 and w2020;
w2022 <= not w331 and w2021;
w2023 <= not w536 and w2022;
w2024 <= not w299 and w1064;
w2025 <= not w77 and not w576;
w2026 <= not w298 and not w493;
w2027 <= not w102 and not w441;
w2028 <= not w34 and not w158;
w2029 <= w2027 and w2028;
w2030 <= w2026 and w2029;
w2031 <= w2025 and w2030;
w2032 <= w2024 and w2031;
w2033 <= not w264 and w2032;
w2034 <= not w85 and w2033;
w2035 <= not w819 and w2034;
w2036 <= not w99 and w2035;
w2037 <= not w307 and w2036;
w2038 <= not w328 and w2037;
w2039 <= not w460 and w2038;
w2040 <= not w449 and not w648;
w2041 <= not w164 and not w602;
w2042 <= not w361 and w2041;
w2043 <= not w537 and w2042;
w2044 <= not w50 and w2043;
w2045 <= not w269 and w2044;
w2046 <= not w181 and w2045;
w2047 <= not w105 and w2046;
w2048 <= not w161 and not w444;
w2049 <= not w1007 and w1063;
w2050 <= not w81 and w2049;
w2051 <= w2048 and w2050;
w2052 <= w1578 and w2051;
w2053 <= w1814 and w2052;
w2054 <= w947 and w2053;
w2055 <= w2047 and w2054;
w2056 <= w1956 and w2055;
w2057 <= w998 and w2056;
w2058 <= w43 and w2057;
w2059 <= not w138 and w2058;
w2060 <= w2040 and w2059;
w2061 <= not w529 and w2060;
w2062 <= not w222 and w2061;
w2063 <= not w332 and not w462;
w2064 <= not w180 and w2063;
w2065 <= not w502 and w2064;
w2066 <= not w558 and w2065;
w2067 <= not w273 and w2066;
w2068 <= not w448 and not w997;
w2069 <= w410 and w1948;
w2070 <= w2068 and w2069;
w2071 <= w2067 and w2070;
w2072 <= w2062 and w2071;
w2073 <= w2039 and w2072;
w2074 <= w1186 and w2073;
w2075 <= w55 and w2074;
w2076 <= w2023 and w2075;
w2077 <= w291 and w2076;
w2078 <= not w453 and w2077;
w2079 <= not w86 and w2078;
w2080 <= not w90 and w2079;
w2081 <= not w370 and w2080;
w2082 <= not w396 and w2081;
w2083 <= not w261 and w2082;
w2084 <= not w303 and w2083;
w2085 <= not w65 and w2084;
w2086 <= not w504 and w2085;
w2087 <= not w590 and w2086;
w2088 <= not w1992 and not w2087;
w2089 <= not w53 and not w1007;
w2090 <= w1263 and w2089;
w2091 <= w1825 and w2090;
w2092 <= w1314 and w2091;
w2093 <= w1063 and w2092;
w2094 <= w2008 and w2093;
w2095 <= w276 and w2094;
w2096 <= not w129 and w2095;
w2097 <= not w1181 and w2096;
w2098 <= not w738 and w2097;
w2099 <= not w370 and w2098;
w2100 <= not w292 and w2099;
w2101 <= not w77 and w2100;
w2102 <= not w206 and w2101;
w2103 <= not w427 and not w449;
w2104 <= not w460 and w2103;
w2105 <= not w328 and not w915;
w2106 <= w291 and w2105;
w2107 <= not w395 and w2106;
w2108 <= w91 and w1828;
w2109 <= not w110 and w2108;
w2110 <= w682 and w708;
w2111 <= w1076 and w2110;
w2112 <= w1391 and w2111;
w2113 <= w2109 and w2112;
w2114 <= w2107 and w2113;
w2115 <= w692 and w2114;
w2116 <= w606 and w2115;
w2117 <= w2104 and w2116;
w2118 <= w1603 and w2117;
w2119 <= w358 and w2118;
w2120 <= w2102 and w2119;
w2121 <= w1182 and w2120;
w2122 <= w443 and w2121;
w2123 <= not w648 and w2122;
w2124 <= not w178 and w2123;
w2125 <= not w2087 and not w2124;
w2126 <= not w92 and not w211;
w2127 <= not w79 and not w1036;
w2128 <= w2126 and w2127;
w2129 <= w2089 and w2128;
w2130 <= w1760 and w2129;
w2131 <= w1485 and w2130;
w2132 <= w2008 and w2131;
w2133 <= not w125 and w2132;
w2134 <= not w213 and w2133;
w2135 <= not w56 and w2134;
w2136 <= not w210 and w2135;
w2137 <= not w108 and w2136;
w2138 <= w655 and w1466;
w2139 <= not w439 and w2138;
w2140 <= not w206 and w2139;
w2141 <= not w30 and w2140;
w2142 <= not w821 and w2141;
w2143 <= not w293 and w2142;
w2144 <= not w649 and not w896;
w2145 <= not w82 and not w127;
w2146 <= w2144 and w2145;
w2147 <= w822 and w2146;
w2148 <= not w216 and w2147;
w2149 <= not w492 and w2148;
w2150 <= not w506 and w2149;
w2151 <= not w163 and w2150;
w2152 <= not w651 and w2151;
w2153 <= not w129 and not w554;
w2154 <= not w760 and w2153;
w2155 <= not w208 and not w441;
w2156 <= w530 and w2155;
w2157 <= w2028 and w2156;
w2158 <= w1004 and w2157;
w2159 <= not w289 and w2158;
w2160 <= not w738 and w2159;
w2161 <= not w302 and w2160;
w2162 <= not w81 and w2161;
w2163 <= not w221 and w2162;
w2164 <= not w180 and w2163;
w2165 <= not w171 and not w395;
w2166 <= w68 and w2165;
w2167 <= w1877 and w2166;
w2168 <= not w687 and w2167;
w2169 <= not w124 and w2168;
w2170 <= not w352 and w2169;
w2171 <= not w388 and w2170;
w2172 <= not w329 and w2171;
w2173 <= not w287 and not w355;
w2174 <= not w440 and w2173;
w2175 <= not w98 and w2174;
w2176 <= not w42 and not w498;
w2177 <= w1698 and w2176;
w2178 <= w2175 and w2177;
w2179 <= w2172 and w2178;
w2180 <= w743 and w2179;
w2181 <= w2164 and w2180;
w2182 <= w1929 and w2181;
w2183 <= w2154 and w2182;
w2184 <= w51 and w2183;
w2185 <= w1324 and w2184;
w2186 <= not w71 and w2185;
w2187 <= not w648 and w2186;
w2188 <= not w576 and w2187;
w2189 <= not w227 and w2188;
w2190 <= not w331 and w2189;
w2191 <= not w183 and w2190;
w2192 <= not w225 and w2191;
w2193 <= not w502 and w2192;
w2194 <= w553 and w1762;
w2195 <= not w174 and w2194;
w2196 <= not w448 and w2195;
w2197 <= not w364 and w2196;
w2198 <= not w681 and not w744;
w2199 <= not w96 and w137;
w2200 <= not w607 and w2199;
w2201 <= w461 and w667;
w2202 <= not w172 and w2201;
w2203 <= w2200 and w2202;
w2204 <= w470 and w2203;
w2205 <= w1090 and w2204;
w2206 <= not w558 and w2205;
w2207 <= not w647 and w2206;
w2208 <= not w371 and w2207;
w2209 <= not w160 and w2208;
w2210 <= not w93 and w2209;
w2211 <= not w431 and not w536;
w2212 <= not w87 and w2211;
w2213 <= not w292 and w2212;
w2214 <= w2210 and w2213;
w2215 <= w300 and w2214;
w2216 <= w2198 and w2215;
w2217 <= w2197 and w2216;
w2218 <= w1203 and w2217;
w2219 <= w2193 and w2218;
w2220 <= w2152 and w2219;
w2221 <= w2143 and w2220;
w2222 <= w2137 and w2221;
w2223 <= w445 and w2222;
w2224 <= not w290 and w2223;
w2225 <= not w190 and w2224;
w2226 <= not w555 and w2225;
w2227 <= not w2124 and not w2226;
w2228 <= not w178 and not w302;
w2229 <= not w163 and w2228;
w2230 <= not w472 and w2229;
w2231 <= not w405 and w2230;
w2232 <= not w81 and not w395;
w2233 <= w762 and w2232;
w2234 <= not w782 and w2233;
w2235 <= not w85 and w2234;
w2236 <= not w225 and w2235;
w2237 <= w1066 and w1411;
w2238 <= not w681 and w2237;
w2239 <= w960 and w2238;
w2240 <= w1468 and w2239;
w2241 <= w751 and w2240;
w2242 <= w142 and w2241;
w2243 <= w2026 and w2242;
w2244 <= w2236 and w2243;
w2245 <= w2231 and w2244;
w2246 <= w2104 and w2245;
w2247 <= w1760 and w2246;
w2248 <= not w164 and w2247;
w2249 <= not w712 and w2248;
w2250 <= not w222 and w2249;
w2251 <= not w538 and w2250;
w2252 <= not w1039 and w2251;
w2253 <= not w106 and not w289;
w2254 <= not w215 and w2253;
w2255 <= not w210 and w2254;
w2256 <= not w227 and w2255;
w2257 <= not w351 and w2256;
w2258 <= not w127 and w2257;
w2259 <= not w99 and w2258;
w2260 <= not w502 and w2259;
w2261 <= not w236 and w372;
w2262 <= not w274 and w2261;
w2263 <= not w292 and w2262;
w2264 <= not w592 and w2263;
w2265 <= not w123 and w2264;
w2266 <= not w536 and not w602;
w2267 <= not w272 and w2266;
w2268 <= not w102 and not w266;
w2269 <= not w187 and w2268;
w2270 <= w822 and w2269;
w2271 <= w2267 and w2270;
w2272 <= w567 and w2271;
w2273 <= w2265 and w2272;
w2274 <= w173 and w2273;
w2275 <= w2260 and w2274;
w2276 <= w831 and w2275;
w2277 <= not w355 and w2276;
w2278 <= not w288 and w2277;
w2279 <= not w90 and w2278;
w2280 <= not w1062 and w2279;
w2281 <= not w498 and not w608;
w2282 <= not w110 and w2281;
w2283 <= not w403 and not w896;
w2284 <= not w524 and not w1181;
w2285 <= w1571 and w1674;
w2286 <= w2284 and w2285;
w2287 <= w2283 and w2286;
w2288 <= w176 and w2287;
w2289 <= not w1037 and w2288;
w2290 <= w2282 and w2289;
w2291 <= not w262 and w2290;
w2292 <= not w529 and w2291;
w2293 <= not w365 and w2292;
w2294 <= not w1138 and w2293;
w2295 <= not w409 and w2294;
w2296 <= not w237 and not w467;
w2297 <= not w26 and not w453;
w2298 <= not w77 and w2297;
w2299 <= w2296 and w2298;
w2300 <= not w216 and w2299;
w2301 <= not w82 and w2300;
w2302 <= not w726 and w2301;
w2303 <= not w428 and w2302;
w2304 <= not w293 and w2303;
w2305 <= not w810 and w2304;
w2306 <= not w263 and not w504;
w2307 <= w728 and w1774;
w2308 <= w243 and w2307;
w2309 <= w2306 and w2308;
w2310 <= w2305 and w2309;
w2311 <= w2295 and w2310;
w2312 <= w2280 and w2311;
w2313 <= w2252 and w2312;
w2314 <= w1602 and w2313;
w2315 <= w872 and w2314;
w2316 <= w1187 and w2315;
w2317 <= not w397 and w2316;
w2318 <= w956 and w2317;
w2319 <= not w650 and w2318;
w2320 <= not w92 and w2319;
w2321 <= not w260 and w2320;
w2322 <= not w821 and w2321;
w2323 <= not w166 and w2322;
w2324 <= not w2226 and not w2323;
w2325 <= not w108 and not w499;
w2326 <= w297 and w2325;
w2327 <= w1814 and w2326;
w2328 <= w1315 and w2327;
w2329 <= w1696 and w2328;
w2330 <= not w58 and w2329;
w2331 <= w1043 and w2330;
w2332 <= not w446 and w2331;
w2333 <= not w53 and w2332;
w2334 <= not w352 and w2333;
w2335 <= not w225 and w2334;
w2336 <= not w712 and w2335;
w2337 <= not w472 and w2336;
w2338 <= not w135 and w2337;
w2339 <= not w207 and w2338;
w2340 <= not w1062 and w2339;
w2341 <= not w34 and not w386;
w2342 <= not w208 and not w227;
w2343 <= not w818 and w2342;
w2344 <= not w363 and w2343;
w2345 <= not w82 and not w206;
w2346 <= w1259 and w2345;
w2347 <= not w574 and w2346;
w2348 <= not w760 and w2347;
w2349 <= not w80 and w2348;
w2350 <= not w175 and w2349;
w2351 <= not w307 and w2350;
w2352 <= not w524 and w2351;
w2353 <= not w572 and not w1037;
w2354 <= not w140 and w2353;
w2355 <= not w1138 and w2354;
w2356 <= not w405 and w2355;
w2357 <= not w527 and w2356;
w2358 <= not w54 and not w77;
w2359 <= not w158 and not w354;
w2360 <= not w183 and not w997;
w2361 <= not w303 and w2360;
w2362 <= w91 and not w867;
w2363 <= w2361 and w2362;
w2364 <= w2359 and w2363;
w2365 <= w2358 and w2364;
w2366 <= w2357 and w2365;
w2367 <= w1066 and w2366;
w2368 <= w2352 and w2367;
w2369 <= w1182 and w2368;
w2370 <= not w171 and w2369;
w2371 <= not w177 and w2370;
w2372 <= not w219 and w2371;
w2373 <= not w65 and w2372;
w2374 <= not w384 and w2373;
w2375 <= w223 and w2374;
w2376 <= not w364 and w2375;
w2377 <= not w236 and not w647;
w2378 <= not w726 and w2377;
w2379 <= not w360 and w2378;
w2380 <= not w592 and w2379;
w2381 <= w2376 and w2380;
w2382 <= w2344 and w2381;
w2383 <= w725 and w2382;
w2384 <= w1975 and w2383;
w2385 <= w600 and w2384;
w2386 <= w539 and w2385;
w2387 <= w2341 and w2386;
w2388 <= w1602 and w2387;
w2389 <= w334 and w2388;
w2390 <= w2003 and w2389;
w2391 <= w2340 and w2390;
w2392 <= not w648 and w2391;
w2393 <= not w168 and w2392;
w2394 <= not w396 and w2393;
w2395 <= not w92 and w2394;
w2396 <= not w558 and w2395;
w2397 <= not w273 and w2396;
w2398 <= not w467 and w2397;
w2399 <= not w601 and w2398;
w2400 <= not w2323 and not w2399;
w2401 <= not w190 and not w552;
w2402 <= not w240 and not w386;
w2403 <= not w301 and not w624;
w2404 <= w137 and not w430;
w2405 <= not w187 and w2404;
w2406 <= w925 and w2405;
w2407 <= w834 and w2406;
w2408 <= w2403 and w2407;
w2409 <= w2283 and w2408;
w2410 <= w2402 and w2409;
w2411 <= w128 and w2410;
w2412 <= w2401 and w2411;
w2413 <= not w331 and w2412;
w2414 <= not w225 and w2413;
w2415 <= not w218 and w2414;
w2416 <= not w460 and w2415;
w2417 <= not w93 and w2416;
w2418 <= not w590 and w2417;
w2419 <= not w102 and not w365;
w2420 <= not w425 and not w449;
w2421 <= not w309 and w2420;
w2422 <= not w538 and w2421;
w2423 <= w300 and w1139;
w2424 <= w235 and w2423;
w2425 <= w2422 and w2424;
w2426 <= w1850 and w2425;
w2427 <= w556 and w2426;
w2428 <= w831 and w2427;
w2429 <= w820 and w2428;
w2430 <= not w1007 and w2429;
w2431 <= not w46 and w2430;
w2432 <= not w744 and w2431;
w2433 <= not w56 and w2432;
w2434 <= not w945 and w2433;
w2435 <= not w706 and w2434;
w2436 <= not w395 and not w529;
w2437 <= not w141 and w2436;
w2438 <= not w178 and w2437;
w2439 <= not w592 and w2438;
w2440 <= not w96 and w2439;
w2441 <= not w607 and w2440;
w2442 <= not w98 and not w1181;
w2443 <= not w355 and not w439;
w2444 <= w577 and w2443;
w2445 <= not w370 and w2444;
w2446 <= not w227 and w2445;
w2447 <= not w454 and w2446;
w2448 <= not w167 and w217;
w2449 <= not w648 and w2448;
w2450 <= not w166 and w2449;
w2451 <= w286 and w2450;
w2452 <= w2447 and w2451;
w2453 <= w2442 and w2452;
w2454 <= w2374 and w2453;
w2455 <= w2441 and w2454;
w2456 <= w2435 and w2455;
w2457 <= w2419 and w2456;
w2458 <= w655 and w2457;
w2459 <= w2418 and w2458;
w2460 <= not w124 and w2459;
w2461 <= not w174 and w2460;
w2462 <= not w352 and w2461;
w2463 <= not w161 and w2462;
w2464 <= not w373 and w2463;
w2465 <= not w498 and w2464;
w2466 <= not w726 and w2465;
w2467 <= not w230 and w2466;
w2468 <= not w228 and w2467;
w2469 <= not w2399 and not w2468;
w2470 <= not w183 and not w262;
w2471 <= not w26 and w2470;
w2472 <= not w208 and w2471;
w2473 <= w559 and w2472;
w2474 <= not w896 and w2473;
w2475 <= not w65 and w2474;
w2476 <= not w160 and w2475;
w2477 <= not w187 and w2476;
w2478 <= not w30 and w2477;
w2479 <= not w333 and not w529;
w2480 <= not w177 and not w440;
w2481 <= not w92 and w2480;
w2482 <= w2362 and w2481;
w2483 <= w2479 and w2482;
w2484 <= w2105 and w2483;
w2485 <= not w190 and w2484;
w2486 <= not w554 and w2485;
w2487 <= not w222 and w2486;
w2488 <= not w241 and w2487;
w2489 <= not w306 and w2488;
w2490 <= not w166 and w2489;
w2491 <= not w174 and not w568;
w2492 <= w573 and w2491;
w2493 <= w924 and w2492;
w2494 <= w1814 and w2493;
w2495 <= w779 and w2494;
w2496 <= w1137 and w2495;
w2497 <= w2490 and w2496;
w2498 <= w2478 and w2497;
w2499 <= w1314 and w2498;
w2500 <= w1324 and w2499;
w2501 <= not w332 and w2500;
w2502 <= not w687 and w2501;
w2503 <= not w269 and w2502;
w2504 <= not w42 and w2503;
w2505 <= not w651 and w2504;
w2506 <= not w504 and w2505;
w2507 <= not w2468 and not w2506;
w2508 <= not w260 and not w818;
w2509 <= not w362 and not w552;
w2510 <= not w189 and w2509;
w2511 <= not w738 and w2510;
w2512 <= not w163 and w2511;
w2513 <= not w126 and w2512;
w2514 <= not w218 and w2513;
w2515 <= not w301 and w2514;
w2516 <= not w424 and w2515;
w2517 <= not w298 and not w810;
w2518 <= not w444 and not w558;
w2519 <= not w333 and not w403;
w2520 <= w2025 and w2519;
w2521 <= not w782 and w2520;
w2522 <= not w110 and w2521;
w2523 <= not w158 and w2522;
w2524 <= not w503 and w2523;
w2525 <= not w275 and w2524;
w2526 <= not w1062 and w2525;
w2527 <= not w175 and not w180;
w2528 <= not w1138 and w2527;
w2529 <= w808 and w1115;
w2530 <= not w30 and w2529;
w2531 <= w2528 and w2530;
w2532 <= w2284 and w2531;
w2533 <= w1774 and w2532;
w2534 <= w912 and w2533;
w2535 <= not w50 and w2534;
w2536 <= not w449 and w2535;
w2537 <= not w370 and w2536;
w2538 <= not w160 and w2537;
w2539 <= not w467 and w2538;
w2540 <= not w16 and w2539;
w2541 <= not w104 and not w472;
w2542 <= not w460 and w2541;
w2543 <= not w396 and not w439;
w2544 <= w1735 and w2543;
w2545 <= w2542 and w2544;
w2546 <= w530 and w2545;
w2547 <= w725 and w2546;
w2548 <= w2540 and w2547;
w2549 <= w2526 and w2548;
w2550 <= w1537 and w2549;
w2551 <= w2518 and w2550;
w2552 <= w2517 and w2551;
w2553 <= not w299 and w2552;
w2554 <= not w103 and w2553;
w2555 <= not w287 and w2554;
w2556 <= not w53 and w2555;
w2557 <= not w359 and w2556;
w2558 <= not w608 and w2557;
w2559 <= not w446 and w551;
w2560 <= not w65 and w2559;
w2561 <= not w129 and not w493;
w2562 <= not w649 and w2561;
w2563 <= w2560 and w2562;
w2564 <= w2306 and w2563;
w2565 <= not w177 and w2564;
w2566 <= not w292 and w2565;
w2567 <= not w647 and w2566;
w2568 <= not w58 and not w328;
w2569 <= not w112 and not w136;
w2570 <= not w187 and w2569;
w2571 <= not w141 and w2570;
w2572 <= not w293 and w2571;
w2573 <= w1513 and w1763;
w2574 <= w2572 and w2573;
w2575 <= w1673 and w2574;
w2576 <= w1354 and w2575;
w2577 <= w746 and w2576;
w2578 <= w2568 and w2577;
w2579 <= w868 and w2578;
w2580 <= w2419 and w2579;
w2581 <= not w332 and w2580;
w2582 <= not w37 and w2581;
w2583 <= not w172 and w2582;
w2584 <= not w497 and w2583;
w2585 <= not w590 and w2584;
w2586 <= not w26 and not w440;
w2587 <= w217 and w2586;
w2588 <= not w462 and w2587;
w2589 <= not w355 and not w537;
w2590 <= not w108 and w2589;
w2591 <= not w428 and w2590;
w2592 <= w2588 and w2591;
w2593 <= w2585 and w2592;
w2594 <= w2567 and w2593;
w2595 <= w2558 and w2594;
w2596 <= w2516 and w2595;
w2597 <= w2508 and w2596;
w2598 <= w94 and w2597;
w2599 <= w914 and w2598;
w2600 <= w655 and w2599;
w2601 <= not w1007 and w2600;
w2602 <= not w404 and w2601;
w2603 <= not w453 and w2602;
w2604 <= not w915 and w2603;
w2605 <= not w212 and w2604;
w2606 <= not w499 and w2605;
w2607 <= not w306 and w2606;
w2608 <= not w123 and w2607;
w2609 <= not w166 and w2608;
w2610 <= not w2506 and not w2609;
w2611 <= not w290 and not w439;
w2612 <= not w175 and w2611;
w2613 <= not w239 and w2612;
w2614 <= w63 and w1056;
w2615 <= not w538 and w2614;
w2616 <= not w1138 and w2615;
w2617 <= not w466 and w2616;
w2618 <= not w157 and not w222;
w2619 <= not w50 and w2618;
w2620 <= w2325 and w2619;
w2621 <= w2068 and w2620;
w2622 <= w1322 and w2621;
w2623 <= w2617 and w2622;
w2624 <= w2260 and w2623;
w2625 <= w1117 and w2624;
w2626 <= w914 and w2625;
w2627 <= w2518 and w2626;
w2628 <= not w104 and w2627;
w2629 <= not w331 and w2628;
w2630 <= not w1039 and w2629;
w2631 <= not w818 and w2630;
w2632 <= not w30 and w2631;
w2633 <= not w357 and not w460;
w2634 <= not w506 and not w744;
w2635 <= not w449 and w2634;
w2636 <= not w274 and w2635;
w2637 <= not w168 and w2636;
w2638 <= not w183 and w2637;
w2639 <= not w536 and not w810;
w2640 <= not w110 and not w230;
w2641 <= w1571 and w2640;
w2642 <= w2639 and w2641;
w2643 <= w2442 and w2642;
w2644 <= not w946 and w2643;
w2645 <= not w430 and w2644;
w2646 <= not w53 and w2645;
w2647 <= not w335 and w2646;
w2648 <= not w712 and w2647;
w2649 <= not w329 and w2648;
w2650 <= not w821 and w2649;
w2651 <= not w205 and w2650;
w2652 <= not w388 and w1717;
w2653 <= not w241 and w2652;
w2654 <= not w184 and w2653;
w2655 <= not w190 and not w498;
w2656 <= not w21 and w2655;
w2657 <= w2238 and w2656;
w2658 <= w2165 and w2657;
w2659 <= w2654 and w2658;
w2660 <= w2585 and w2659;
w2661 <= w2651 and w2660;
w2662 <= w2638 and w2661;
w2663 <= w2633 and w2662;
w2664 <= w1118 and w2663;
w2665 <= w2632 and w2664;
w2666 <= w2613 and w2665;
w2667 <= w872 and w2666;
w2668 <= not w554 and w2667;
w2669 <= not w574 and w2668;
w2670 <= not w135 and w2669;
w2671 <= not w945 and w2670;
w2672 <= not w2609 and not w2671;
w2673 <= not w164 and not w1181;
w2674 <= not w269 and not w591;
w2675 <= not w86 and not w106;
w2676 <= not w290 and w739;
w2677 <= not w810 and w2676;
w2678 <= w2675 and w2677;
w2679 <= w2674 and w2678;
w2680 <= w1063 and w2679;
w2681 <= not w70 and w2680;
w2682 <= not w744 and w2681;
w2683 <= not w158 and w2682;
w2684 <= not w650 and w2683;
w2685 <= not w373 and w2684;
w2686 <= not w187 and w2685;
w2687 <= not w371 and not w502;
w2688 <= not w335 and w455;
w2689 <= w2687 and w2688;
w2690 <= w2380 and w2689;
w2691 <= w2479 and w2690;
w2692 <= w429 and w2691;
w2693 <= not w87 and not w552;
w2694 <= not w53 and w2693;
w2695 <= w1249 and w2694;
w2696 <= w2692 and w2695;
w2697 <= w2686 and w2696;
w2698 <= w2673 and w2697;
w2699 <= w1188 and w2698;
w2700 <= w2586 and w2699;
w2701 <= w442 and w2700;
w2702 <= not w189 and w2701;
w2703 <= not w263 and w2702;
w2704 <= not w234 and w2703;
w2705 <= not w503 and w2704;
w2706 <= not w178 and w2705;
w2707 <= not w466 and w2706;
w2708 <= not w681 and not w946;
w2709 <= not w337 and w2708;
w2710 <= not w240 and w2709;
w2711 <= not w760 and w2710;
w2712 <= not w607 and w2711;
w2713 <= not w306 and w2712;
w2714 <= w501 and w1662;
w2715 <= not w361 and w2714;
w2716 <= not w302 and w2715;
w2717 <= not w80 and w2716;
w2718 <= w353 and not w427;
w2719 <= not w180 and w2718;
w2720 <= w567 and w2719;
w2721 <= w139 and w2720;
w2722 <= w2717 and w2721;
w2723 <= w2713 and w2722;
w2724 <= w1929 and w2723;
w2725 <= w450 and w2724;
w2726 <= w1172 and w2725;
w2727 <= w569 and w2726;
w2728 <= not w351 and w2727;
w2729 <= not w649 and w2728;
w2730 <= not w328 and w2729;
w2731 <= not w424 and w2730;
w2732 <= w960 and w1537;
w2733 <= w1361 and w2732;
w2734 <= w589 and w2733;
w2735 <= not w1007 and w2734;
w2736 <= not w444 and w2735;
w2737 <= not w82 and w2736;
w2738 <= not w65 and w2737;
w2739 <= not w460 and w2738;
w2740 <= not w62 and w2739;
w2741 <= not w590 and w2740;
w2742 <= not w67 and not w260;
w2743 <= not w129 and not w821;
w2744 <= not w228 and not w307;
w2745 <= not w99 and w2008;
w2746 <= not w212 and w2745;
w2747 <= w1763 and w2746;
w2748 <= w2744 and w2747;
w2749 <= w2743 and w2748;
w2750 <= w2742 and w2749;
w2751 <= w1644 and w2750;
w2752 <= w2741 and w2751;
w2753 <= w2731 and w2752;
w2754 <= w2707 and w2753;
w2755 <= w724 and w2754;
w2756 <= w1512 and w2755;
w2757 <= w1852 and w2756;
w2758 <= w468 and w2757;
w2759 <= w356 and w2758;
w2760 <= w2211 and w2759;
w2761 <= not w219 and w2760;
w2762 <= not w81 and w2761;
w2763 <= not w266 and w2762;
w2764 <= not w209 and w2763;
w2765 <= w2609 and not w2671;
w2766 <= not w2764 and w2765;
w2767 <= not w2672 and not w2766;
w2768 <= w2506 and w2609;
w2769 <= not w2610 and not w2768;
w2770 <= not w2767 and w2769;
w2771 <= not w2610 and not w2770;
w2772 <= w2468 and w2506;
w2773 <= not w2507 and not w2772;
w2774 <= not w2771 and w2773;
w2775 <= not w2507 and not w2774;
w2776 <= w2399 and w2468;
w2777 <= not w2469 and not w2776;
w2778 <= not w2775 and w2777;
w2779 <= not w2469 and not w2778;
w2780 <= w2323 and w2399;
w2781 <= not w2400 and not w2780;
w2782 <= not w2779 and w2781;
w2783 <= not w2400 and not w2782;
w2784 <= w2226 and w2323;
w2785 <= not w2324 and not w2784;
w2786 <= not w2783 and w2785;
w2787 <= not w2324 and not w2786;
w2788 <= w2124 and w2226;
w2789 <= not w2227 and not w2788;
w2790 <= not w2787 and w2789;
w2791 <= not w2227 and not w2790;
w2792 <= w2087 and w2124;
w2793 <= not w2125 and not w2792;
w2794 <= not w2791 and w2793;
w2795 <= not w2125 and not w2794;
w2796 <= w1992 and w2087;
w2797 <= not w2088 and not w2796;
w2798 <= not w2795 and w2797;
w2799 <= not w2088 and not w2798;
w2800 <= w1927 and w1992;
w2801 <= not w1993 and not w2800;
w2802 <= not w2799 and w2801;
w2803 <= not w1993 and not w2802;
w2804 <= w1848 and w1927;
w2805 <= not w1928 and not w2804;
w2806 <= not w2803 and w2805;
w2807 <= not w1928 and not w2806;
w2808 <= w1812 and w1848;
w2809 <= not w1849 and not w2808;
w2810 <= not w2807 and w2809;
w2811 <= not w1849 and not w2810;
w2812 <= w1714 and w1812;
w2813 <= not w1813 and not w2812;
w2814 <= not w2811 and w2813;
w2815 <= not w1813 and not w2814;
w2816 <= w1600 and w1714;
w2817 <= not w1715 and not w2816;
w2818 <= not w2815 and w2817;
w2819 <= not w1715 and not w2818;
w2820 <= w1507 and w1600;
w2821 <= not w1601 and not w2820;
w2822 <= not w2819 and w2821;
w2823 <= not w1601 and not w2822;
w2824 <= w1407 and w1507;
w2825 <= not w1508 and not w2824;
w2826 <= not w2823 and w2825;
w2827 <= not w1508 and not w2826;
w2828 <= w1299 and w1407;
w2829 <= not w1408 and not w2828;
w2830 <= not w2827 and w2829;
w2831 <= not w1408 and not w2830;
w2832 <= w1170 and w1299;
w2833 <= not w1300 and not w2832;
w2834 <= not w2831 and w2833;
w2835 <= not w1300 and not w2834;
w2836 <= w1113 and w1170;
w2837 <= not w1171 and not w2836;
w2838 <= not w2835 and w2837;
w2839 <= not w1171 and not w2838;
w2840 <= w995 and w1113;
w2841 <= not w1114 and not w2840;
w2842 <= not w2839 and w2841;
w2843 <= not w1114 and not w2842;
w2844 <= w893 and w995;
w2845 <= not w996 and not w2844;
w2846 <= not w2843 and w2845;
w2847 <= not w996 and not w2846;
w2848 <= w802 and w893;
w2849 <= not w894 and not w2848;
w2850 <= not w2847 and w2849;
w2851 <= not w894 and not w2850;
w2852 <= w645 and w802;
w2853 <= not w803 and not w2852;
w2854 <= not w2851 and w2853;
w2855 <= not w803 and not w2854;
w2856 <= w522 and w645;
w2857 <= not w646 and not w2856;
w2858 <= not w2855 and w2857;
w2859 <= not w646 and not w2858;
w2860 <= w327 and w522;
w2861 <= not w523 and not w2860;
w2862 <= not w2859 and w2861;
w2863 <= not w523 and not w2862;
w2864 <= not w141 and not w262;
w2865 <= not w403 and w2864;
w2866 <= not w590 and w2865;
w2867 <= w2025 and w2866;
w2868 <= not w1007 and w2867;
w2869 <= not w492 and w2868;
w2870 <= not w361 and w2869;
w2871 <= not w572 and w2870;
w2872 <= not w241 and w2871;
w2873 <= not w607 and w2872;
w2874 <= not w272 and w2873;
w2875 <= not w706 and w2874;
w2876 <= not w84 and w1491;
w2877 <= not w503 and w2876;
w2878 <= not w34 and w2877;
w2879 <= w925 and w1343;
w2880 <= w2878 and w2879;
w2881 <= w2875 and w2880;
w2882 <= w2154 and w2881;
w2883 <= w1115 and w2882;
w2884 <= not w236 and w2883;
w2885 <= not w211 and w2884;
w2886 <= not w290 and w2885;
w2887 <= not w270 and w2886;
w2888 <= not w574 and w2887;
w2889 <= not w649 and w2888;
w2890 <= not w209 and w2889;
w2891 <= not w175 and w2890;
w2892 <= not w212 and w2891;
w2893 <= not w260 and w2892;
w2894 <= w2198 and w2687;
w2895 <= not w397 and w2894;
w2896 <= not w915 and w2895;
w2897 <= not w648 and w1695;
w2898 <= not w216 and w2897;
w2899 <= w767 and w1358;
w2900 <= w2165 and w2899;
w2901 <= w2898 and w2900;
w2902 <= w2896 and w2901;
w2903 <= w1851 and w2902;
w2904 <= w1956 and w2903;
w2905 <= w223 and w2904;
w2906 <= w468 and w2905;
w2907 <= w1760 and w2906;
w2908 <= w2401 and w2907;
w2909 <= not w529 and w2908;
w2910 <= not w405 and w2909;
w2911 <= not w527 and w2910;
w2912 <= not w601 and w2911;
w2913 <= not w424 and w2912;
w2914 <= not w184 and w2913;
w2915 <= not w106 and w2344;
w2916 <= not w240 and w2915;
w2917 <= not w37 and w2916;
w2918 <= not w266 and w2917;
w2919 <= not w218 and w2918;
w2920 <= not w307 and w2919;
w2921 <= not w945 and w2920;
w2922 <= not w454 and w2921;
w2923 <= w569 and w944;
w2924 <= not w224 and w2923;
w2925 <= not w466 and w2924;
w2926 <= not w287 and w356;
w2927 <= not w273 and w2926;
w2928 <= not w56 and not w112;
w2929 <= not w333 and w2928;
w2930 <= not w50 and w2929;
w2931 <= w2048 and w2930;
w2932 <= w2927 and w2931;
w2933 <= w2925 and w2932;
w2934 <= w1758 and w2933;
w2935 <= w2922 and w2934;
w2936 <= w2914 and w2935;
w2937 <= w179 and w2936;
w2938 <= w2893 and w2937;
w2939 <= w525 and w2938;
w2940 <= w1324 and w2939;
w2941 <= not w71 and w2940;
w2942 <= not w441 and w2941;
w2943 <= not w292 and w2942;
w2944 <= not w261 and w2943;
w2945 <= not w1138 and w2944;
w2946 <= not w135 and w2945;
w2947 <= not w306 and w2946;
w2948 <= not w327 and not w2947;
w2949 <= w327 and w2947;
w2950 <= not w2948 and not w2949;
w2951 <= not w2863 and w2950;
w2952 <= w2863 and not w2950;
w2953 <= not w2951 and not w2952;
w2954 <= w10 and w2953;
w2955 <= not a(31) and not w9;
w2956 <= not w2947 and w2955;
w2957 <= a(30) and w9;
w2958 <= a(31) and w2957;
w2959 <= not w522 and w2958;
w2960 <= a(30) and not a(31);
w2961 <= not a(30) and a(31);
w2962 <= not w2960 and not w2961;
w2963 <= w9 and not w2962;
w2964 <= not w327 and w2963;
w2965 <= not w2959 and not w2964;
w2966 <= not w2956 and w2965;
w2967 <= not w2954 and w2966;
w2968 <= not w210 and w2695;
w2969 <= not w227 and w2968;
w2970 <= not w292 and w2969;
w2971 <= not w209 and w2970;
w2972 <= not w180 and w2971;
w2973 <= not w558 and w2972;
w2974 <= not w424 and w2973;
w2975 <= not w221 and not w388;
w2976 <= not w260 and not w1062;
w2977 <= not w123 and not w591;
w2978 <= not w125 and not w462;
w2979 <= not w335 and not w648;
w2980 <= not w126 and w2979;
w2981 <= w2978 and w2980;
w2982 <= w2977 and w2981;
w2983 <= w2976 and w2982;
w2984 <= w2975 and w2983;
w2985 <= w1716 and w2984;
w2986 <= w220 and w2985;
w2987 <= w2974 and w2986;
w2988 <= w468 and w2987;
w2989 <= w1076 and w2988;
w2990 <= not w444 and w2989;
w2991 <= not w602 and w2990;
w2992 <= not w498 and w2991;
w2993 <= not w576 and not w687;
w2994 <= not w572 and w2993;
w2995 <= not w211 and w2994;
w2996 <= not w332 and w2995;
w2997 <= not w425 and w2996;
w2998 <= not w135 and w2997;
w2999 <= not w96 and w2998;
w3000 <= not w945 and w2999;
w3001 <= not w1181 and w2568;
w3002 <= not w70 and w3001;
w3003 <= not w497 and w3002;
w3004 <= w308 and w508;
w3005 <= w1373 and w3004;
w3006 <= w3003 and w3005;
w3007 <= w429 and w3006;
w3008 <= w866 and w3007;
w3009 <= w2252 and w3008;
w3010 <= w2586 and w3009;
w3011 <= w3000 and w3010;
w3012 <= w2992 and w3011;
w3013 <= w739 and w3012;
w3014 <= not w362 and w3013;
w3015 <= not w288 and w3014;
w3016 <= not w1037 and w3015;
w3017 <= not w138 and w3016;
w3018 <= not w175 and w3017;
w3019 <= not w138 and not w726;
w3020 <= not w467 and w3019;
w3021 <= w658 and w3020;
w3022 <= w550 and w3021;
w3023 <= not w1181 and w3022;
w3024 <= not w70 and w3023;
w3025 <= not w263 and w3024;
w3026 <= not w225 and w3025;
w3027 <= not w896 and w3026;
w3028 <= not w77 and w3027;
w3029 <= not w293 and w3028;
w3030 <= w432 and w2994;
w3031 <= w3029 and w3030;
w3032 <= w2633 and w3031;
w3033 <= w2508 and w3032;
w3034 <= w1762 and w3033;
w3035 <= w1819 and w3034;
w3036 <= not w71 and w3035;
w3037 <= not w112 and w3036;
w3038 <= not w53 and w3037;
w3039 <= not w163 and w3038;
w3040 <= not w222 and w3039;
w3041 <= not w440 and w3040;
w3042 <= not w105 and w3041;
w3043 <= not w601 and w3042;
w3044 <= not w397 and w2126;
w3045 <= not w648 and w3044;
w3046 <= not w216 and w3045;
w3047 <= not w108 and w3046;
w3048 <= not w1138 and w3047;
w3049 <= not w210 and w2282;
w3050 <= not w103 and w903;
w3051 <= w1268 and w3050;
w3052 <= w3049 and w3051;
w3053 <= w1067 and w3052;
w3054 <= w3048 and w3053;
w3055 <= w1852 and w3054;
w3056 <= w2613 and w3055;
w3057 <= w1716 and w3056;
w3058 <= w1301 and w3057;
w3059 <= w1183 and w3058;
w3060 <= not w177 and w3059;
w3061 <= not w126 and w3060;
w3062 <= not w62 and w3061;
w3063 <= w553 and not w782;
w3064 <= w832 and w3063;
w3065 <= w374 and w3064;
w3066 <= w625 and w3065;
w3067 <= w2026 and w3066;
w3068 <= w1061 and w3067;
w3069 <= w1423 and w3068;
w3070 <= w3062 and w3069;
w3071 <= w447 and w3070;
w3072 <= w3043 and w3071;
w3073 <= w1929 and w3072;
w3074 <= w1172 and w3073;
w3075 <= w276 and w3074;
w3076 <= not w1241 and w3075;
w3077 <= not w396 and w3076;
w3078 <= not w338 and w3077;
w3079 <= not w427 and w3078;
w3080 <= not w98 and w3079;
w3081 <= not w206 and w3080;
w3082 <= not w269 and not w397;
w3083 <= not w466 and w3082;
w3084 <= w63 and w3083;
w3085 <= w2402 and w3084;
w3086 <= not w440 and w3085;
w3087 <= not w401 and w3086;
w3088 <= not w454 and w3087;
w3089 <= not w186 and w3088;
w3090 <= not w298 and w3089;
w3091 <= w811 and w2743;
w3092 <= not w337 and w3091;
w3093 <= not w395 and w3092;
w3094 <= not w233 and w3093;
w3095 <= not w260 and not w738;
w3096 <= not w647 and w682;
w3097 <= not w945 and w3096;
w3098 <= not w103 and not w360;
w3099 <= not w409 and w3098;
w3100 <= not w157 and w3099;
w3101 <= w2284 and w3100;
w3102 <= w3097 and w3101;
w3103 <= w3095 and w3102;
w3104 <= w600 and w3103;
w3105 <= w2568 and w3104;
w3106 <= w998 and w3105;
w3107 <= w1074 and w3106;
w3108 <= w739 and w3107;
w3109 <= w3094 and w3108;
w3110 <= w745 and w3109;
w3111 <= w276 and w3110;
w3112 <= not w71 and w3111;
w3113 <= not w190 and w3112;
w3114 <= not w591 and w3113;
w3115 <= not w352 and w3114;
w3116 <= w336 and w445;
w3117 <= w128 and w3116;
w3118 <= not w46 and w3117;
w3119 <= not w138 and w3118;
w3120 <= not w303 and w3119;
w3121 <= not w98 and w3120;
w3122 <= not w208 and w3121;
w3123 <= not w172 and w3122;
w3124 <= not w160 and w3123;
w3125 <= not w230 and w3124;
w3126 <= not w205 and w3125;
w3127 <= w442 and not w946;
w3128 <= not w211 and not w265;
w3129 <= not w87 and w3128;
w3130 <= w3127 and w3129;
w3131 <= w1358 and w3130;
w3132 <= w1490 and w3131;
w3133 <= w3126 and w3132;
w3134 <= w1760 and w3133;
w3135 <= w666 and w3134;
w3136 <= w1187 and w3135;
w3137 <= not w449 and w3136;
w3138 <= not w262 and w3137;
w3139 <= not w77 and w3138;
w3140 <= not w34 and w3139;
w3141 <= not w159 and not w264;
w3142 <= not w552 and w3141;
w3143 <= not w171 and w3142;
w3144 <= not w355 and w3143;
w3145 <= not w687 and w3144;
w3146 <= not w1036 and w3145;
w3147 <= not w183 and w3146;
w3148 <= not w37 and w3147;
w3149 <= not w760 and w3148;
w3150 <= not w102 and w3149;
w3151 <= not w726 and w3150;
w3152 <= not w273 and w3151;
w3153 <= not w527 and w3152;
w3154 <= not w123 and w3153;
w3155 <= w609 and w1466;
w3156 <= not w65 and w3155;
w3157 <= not w403 and w3156;
w3158 <= not w1062 and w3157;
w3159 <= not w30 and w3158;
w3160 <= not w364 and w3159;
w3161 <= not w168 and not w330;
w3162 <= w2267 and w3161;
w3163 <= w3160 and w3162;
w3164 <= w3154 and w3163;
w3165 <= w3140 and w3164;
w3166 <= w3115 and w3165;
w3167 <= w3090 and w3166;
w3168 <= w55 and w3167;
w3169 <= w556 and w3168;
w3170 <= w1509 and w3169;
w3171 <= not w648 and w3170;
w3172 <= not w293 and w3171;
w3173 <= not w93 and w3172;
w3174 <= not w184 and w3173;
w3175 <= not w3081 and not w3174;
w3176 <= w3081 and w3174;
w3177 <= not w3175 and not w3176;
w3178 <= not a(20) and w3177;
w3179 <= not w3175 and not w3178;
w3180 <= w3018 and not w3179;
w3181 <= not w3018 and w3179;
w3182 <= not w3180 and not w3181;
w3183 <= not w2967 and w3182;
w3184 <= not w2967 and not w3183;
w3185 <= w3182 and not w3183;
w3186 <= not w3184 and not w3185;
w3187 <= not w108 and not w161;
w3188 <= not w333 and w2640;
w3189 <= not w89 and w3188;
w3190 <= not w216 and w3189;
w3191 <= not w591 and w3190;
w3192 <= not w572 and w3191;
w3193 <= not w127 and w3192;
w3194 <= not w726 and w3193;
w3195 <= not w190 and w1329;
w3196 <= not w208 and w3195;
w3197 <= not w289 and w474;
w3198 <= not w159 and w3197;
w3199 <= not w601 and w3198;
w3200 <= not w206 and w406;
w3201 <= not w298 and w3200;
w3202 <= w998 and w1063;
w3203 <= not w160 and w3202;
w3204 <= w3201 and w3203;
w3205 <= w3199 and w3204;
w3206 <= w2866 and w3205;
w3207 <= w947 and w3206;
w3208 <= w3196 and w3207;
w3209 <= w3194 and w3208;
w3210 <= w708 and w3209;
w3211 <= w226 and w3210;
w3212 <= not w288 and w3211;
w3213 <= not w576 and w3212;
w3214 <= not w287 and w3213;
w3215 <= not w498 and w3214;
w3216 <= not w568 and w3215;
w3217 <= not w123 and w3216;
w3218 <= not w492 and not w1181;
w3219 <= not w738 and w3218;
w3220 <= not w269 and w3219;
w3221 <= not w234 and w3220;
w3222 <= not w462 and w3221;
w3223 <= not w574 and w3222;
w3224 <= not w460 and w3223;
w3225 <= not w205 and w3224;
w3226 <= not w215 and w655;
w3227 <= not w650 and w3226;
w3228 <= not w896 and w3227;
w3229 <= not w77 and w3228;
w3230 <= not w867 and w3229;
w3231 <= not w466 and w3230;
w3232 <= not w140 and w2586;
w3233 <= not w157 and w3232;
w3234 <= not w330 and not w387;
w3235 <= not w424 and w3234;
w3236 <= w3233 and w3235;
w3237 <= w3231 and w3236;
w3238 <= w1458 and w3237;
w3239 <= w3225 and w3238;
w3240 <= w1414 and w3239;
w3241 <= w63 and w3240;
w3242 <= w358 and w3241;
w3243 <= w666 and w3242;
w3244 <= w442 and w3243;
w3245 <= not w328 and w3244;
w3246 <= not w386 and w3245;
w3247 <= not w166 and w3246;
w3248 <= not w332 and not w370;
w3249 <= not w373 and w3248;
w3250 <= w1006 and w3249;
w3251 <= w1866 and w3250;
w3252 <= w459 and w3251;
w3253 <= w2172 and w3252;
w3254 <= w3247 and w3253;
w3255 <= w3217 and w3254;
w3256 <= w807 and w3255;
w3257 <= w3187 and w3256;
w3258 <= w739 and w3257;
w3259 <= w505 and w3258;
w3260 <= not w168 and w3259;
w3261 <= not w529 and w3260;
w3262 <= not w93 and w3261;
w3263 <= w3081 and not w3262;
w3264 <= not w3081 and w3262;
w3265 <= w2855 and not w2857;
w3266 <= not w2858 and not w3265;
w3267 <= w10 and w3266;
w3268 <= not w522 and w2955;
w3269 <= not w802 and w2958;
w3270 <= not w645 and w2963;
w3271 <= not w3269 and not w3270;
w3272 <= not w3268 and w3271;
w3273 <= not w3267 and w3272;
w3274 <= not w3263 and not w3273;
w3275 <= not w3264 and w3274;
w3276 <= not w3263 and not w3275;
w3277 <= not a(20) and not w3178;
w3278 <= not w3176 and w3179;
w3279 <= not w3277 and not w3278;
w3280 <= not w3276 and not w3279;
w3281 <= w2859 and not w2861;
w3282 <= not w2862 and not w3281;
w3283 <= w10 and w3282;
w3284 <= not w327 and w2955;
w3285 <= not w645 and w2958;
w3286 <= not w522 and w2963;
w3287 <= not w3285 and not w3286;
w3288 <= not w3284 and w3287;
w3289 <= not w3283 and w3288;
w3290 <= w3276 and w3279;
w3291 <= not w3280 and not w3290;
w3292 <= not w3289 and w3291;
w3293 <= not w3280 and not w3292;
w3294 <= not w3186 and not w3293;
w3295 <= w3186 and w3293;
w3296 <= not w3294 and not w3295;
w3297 <= a(28) and not a(29);
w3298 <= not a(28) and a(29);
w3299 <= not w3297 and not w3298;
w3300 <= a(26) and not a(27);
w3301 <= not a(26) and a(27);
w3302 <= not w3300 and not w3301;
w3303 <= not w3299 and not w3302;
w3304 <= not w404 and not w591;
w3305 <= not w945 and w3304;
w3306 <= w2361 and w3305;
w3307 <= w2296 and w3306;
w3308 <= not w129 and w3307;
w3309 <= not w681 and w3308;
w3310 <= not w274 and w3309;
w3311 <= not w80 and w3310;
w3312 <= not w502 and w3311;
w3313 <= not w328 and w3312;
w3314 <= not w81 and not w471;
w3315 <= not w363 and w3314;
w3316 <= not w236 and w3315;
w3317 <= not w446 and w3316;
w3318 <= not w396 and w3317;
w3319 <= not w498 and w3318;
w3320 <= not w624 and w3319;
w3321 <= not w135 and w3320;
w3322 <= not w1241 and w2443;
w3323 <= not w89 and w3322;
w3324 <= not w352 and w3323;
w3325 <= not w307 and not w362;
w3326 <= not w267 and w3325;
w3327 <= w872 and w1116;
w3328 <= not w576 and w3327;
w3329 <= w1327 and w1674;
w3330 <= w3328 and w3329;
w3331 <= w3326 and w3330;
w3332 <= w3324 and w3331;
w3333 <= w3321 and w3332;
w3334 <= w226 and w3333;
w3335 <= not w552 and w3334;
w3336 <= not w70 and w3335;
w3337 <= not w395 and w3336;
w3338 <= not w386 and w3337;
w3339 <= not w272 and w3338;
w3340 <= not w810 and w3339;
w3341 <= not w602 and w2008;
w3342 <= not w687 and w3341;
w3343 <= not w53 and w3342;
w3344 <= not w189 and not w270;
w3345 <= w235 and w897;
w3346 <= w3344 and w3345;
w3347 <= not w1007 and w3346;
w3348 <= not w448 and w3347;
w3349 <= not w126 and w3348;
w3350 <= not w647 and w3349;
w3351 <= w51 and w450;
w3352 <= w980 and w3351;
w3353 <= w3201 and w3352;
w3354 <= w1323 and w3353;
w3355 <= w1067 and w3354;
w3356 <= w3350 and w3355;
w3357 <= w3343 and w3356;
w3358 <= w1463 and w3357;
w3359 <= w808 and w3358;
w3360 <= w1117 and w3359;
w3361 <= w655 and w3360;
w3362 <= not w56 and w3361;
w3363 <= not w240 and w3362;
w3364 <= not w161 and w3363;
w3365 <= not w338 and w3364;
w3366 <= not w141 and w3365;
w3367 <= not w427 and w3366;
w3368 <= not w287 and w1076;
w3369 <= not w472 and w3368;
w3370 <= not w538 and w3369;
w3371 <= not w503 and not w651;
w3372 <= not w77 and w3371;
w3373 <= not w21 and not w175;
w3374 <= w3372 and w3373;
w3375 <= w3370 and w3374;
w3376 <= w3160 and w3375;
w3377 <= w3367 and w3376;
w3378 <= w3340 and w3377;
w3379 <= w2675 and w3378;
w3380 <= w3313 and w3379;
w3381 <= w182 and w3380;
w3382 <= w1852 and w3381;
w3383 <= w426 and w3382;
w3384 <= w913 and w3383;
w3385 <= w745 and w3384;
w3386 <= not w397 and w3385;
w3387 <= not w712 and w3386;
w3388 <= not w160 and w3387;
w3389 <= not w239 and w3388;
w3390 <= not w230 and w3389;
w3391 <= not w454 and w3390;
w3392 <= w3299 and not w3302;
w3393 <= not w3391 and w3392;
w3394 <= not w54 and not w206;
w3395 <= not w189 and w3394;
w3396 <= not w431 and w3395;
w3397 <= not w471 and w3396;
w3398 <= not w647 and w3397;
w3399 <= not w945 and w3398;
w3400 <= w727 and w2026;
w3401 <= not w1036 and w3400;
w3402 <= not w231 and w3401;
w3403 <= not w915 and w3402;
w3404 <= not w558 and w3403;
w3405 <= not w460 and w3404;
w3406 <= not w266 and w2040;
w3407 <= not w388 and w3406;
w3408 <= w353 and not w404;
w3409 <= not w409 and w3408;
w3410 <= w689 and w3161;
w3411 <= w3409 and w3410;
w3412 <= w2491 and w3411;
w3413 <= w528 and w3412;
w3414 <= w372 and w3413;
w3415 <= w1536 and w3414;
w3416 <= w3407 and w3415;
w3417 <= w550 and w3416;
w3418 <= w981 and w3417;
w3419 <= w3405 and w3418;
w3420 <= w1511 and w3419;
w3421 <= w505 and w3420;
w3422 <= not w265 and w3421;
w3423 <= not w237 and w3422;
w3424 <= not w99 and w3423;
w3425 <= not w92 and not w506;
w3426 <= w336 and w2048;
w3427 <= w1466 and w3426;
w3428 <= not w290 and w3427;
w3429 <= not w219 and w3428;
w3430 <= not w712 and w3429;
w3431 <= not w141 and w3430;
w3432 <= not w172 and w3431;
w3433 <= w876 and w1190;
w3434 <= w2155 and w3433;
w3435 <= w1942 and w3434;
w3436 <= w3432 and w3435;
w3437 <= w549 and w3436;
w3438 <= w1956 and w3437;
w3439 <= w226 and w3438;
w3440 <= w1204 and w3439;
w3441 <= not w552 and w3440;
w3442 <= not w159 and w3441;
w3443 <= not w354 and w3442;
w3444 <= w3425 and w3443;
w3445 <= not w301 and w3444;
w3446 <= not w183 and not w361;
w3447 <= not w650 and w3446;
w3448 <= w903 and not w997;
w3449 <= not w360 and w3448;
w3450 <= w107 and w3449;
w3451 <= w3447 and w3450;
w3452 <= w1957 and w3451;
w3453 <= w3445 and w3452;
w3454 <= not w782 and w3453;
w3455 <= not w896 and w3454;
w3456 <= not w180 and w3455;
w3457 <= not w56 and not w80;
w3458 <= not w273 and w3457;
w3459 <= not w221 and not w267;
w3460 <= w3233 and w3459;
w3461 <= w3458 and w3460;
w3462 <= w465 and w3461;
w3463 <= w1521 and w3462;
w3464 <= w400 and w3463;
w3465 <= w3456 and w3464;
w3466 <= w3424 and w3465;
w3467 <= w3399 and w3466;
w3468 <= w964 and w3467;
w3469 <= w1463 and w3468;
w3470 <= w1189 and w3469;
w3471 <= w526 and w3470;
w3472 <= not w269 and w3471;
w3473 <= not w127 and w3472;
w3474 <= not w306 and w3473;
w3475 <= not w14 and not w17;
w3476 <= not w3299 and w3302;
w3477 <= not w3475 and w3476;
w3478 <= not w3474 and w3477;
w3479 <= not w168 and not w819;
w3480 <= not w648 and not w726;
w3481 <= not w310 and w3480;
w3482 <= not w267 and w3481;
w3483 <= not w504 and w3482;
w3484 <= not w161 and not w1062;
w3485 <= w1895 and w3484;
w3486 <= w3483 and w3485;
w3487 <= w1945 and w3486;
w3488 <= w1414 and w3487;
w3489 <= w3479 and w3488;
w3490 <= w1509 and w3489;
w3491 <= w356 and w3490;
w3492 <= not w289 and w3491;
w3493 <= not w269 and w3492;
w3494 <= not w558 and w3493;
w3495 <= w51 and not w1241;
w3496 <= not w441 and w3495;
w3497 <= not w261 and w3496;
w3498 <= not w503 and w3497;
w3499 <= not w365 and w3498;
w3500 <= not w357 and w3499;
w3501 <= not w430 and not w554;
w3502 <= not w292 and w3501;
w3503 <= not w712 and w3502;
w3504 <= not w425 and w3503;
w3505 <= not w363 and w2517;
w3506 <= w2202 and w3505;
w3507 <= w1948 and w3506;
w3508 <= w2283 and w3507;
w3509 <= w3504 and w3508;
w3510 <= not w397 and w3509;
w3511 <= not w498 and w3510;
w3512 <= not w471 and w3511;
w3513 <= not w67 and w3512;
w3514 <= not w273 and w3513;
w3515 <= not w272 and w3514;
w3516 <= not w290 and not w361;
w3517 <= not w331 and w3516;
w3518 <= not w405 and w3517;
w3519 <= w1265 and w1761;
w3520 <= not w333 and w3519;
w3521 <= not w30 and w3520;
w3522 <= not w293 and w3521;
w3523 <= w3518 and w3522;
w3524 <= w3515 and w3523;
w3525 <= w1863 and w3524;
w3526 <= w3500 and w3525;
w3527 <= w156 and w3526;
w3528 <= w1622 and w3527;
w3529 <= w3494 and w3528;
w3530 <= not w171 and w3529;
w3531 <= not w70 and w3530;
w3532 <= not w215 and w3531;
w3533 <= not w1036 and w3532;
w3534 <= not w449 and w3533;
w3535 <= not w240 and w3534;
w3536 <= not w624 and w3535;
w3537 <= not w239 and w3536;
w3538 <= not w21 and w3537;
w3539 <= not w424 and w3538;
w3540 <= not w706 and w3539;
w3541 <= w3302 and w3475;
w3542 <= not w3540 and w3541;
w3543 <= not w3478 and not w3542;
w3544 <= not w3393 and w3543;
w3545 <= not w3303 and w3544;
w3546 <= not w3474 and not w3540;
w3547 <= not w2947 and not w3474;
w3548 <= not w2948 and not w2951;
w3549 <= w2947 and w3474;
w3550 <= not w3547 and not w3549;
w3551 <= not w3548 and w3550;
w3552 <= not w3547 and not w3551;
w3553 <= w3474 and w3540;
w3554 <= not w3546 and not w3553;
w3555 <= not w3552 and w3554;
w3556 <= not w3546 and not w3555;
w3557 <= not w3391 and not w3540;
w3558 <= w3391 and w3540;
w3559 <= not w3557 and not w3558;
w3560 <= not w3556 and w3559;
w3561 <= w3556 and not w3559;
w3562 <= not w3560 and not w3561;
w3563 <= w3544 and not w3562;
w3564 <= not w3545 and not w3563;
w3565 <= a(29) and not w3564;
w3566 <= not a(29) and w3564;
w3567 <= not w3565 and not w3566;
w3568 <= w3296 and not w3567;
w3569 <= not w3294 and not w3568;
w3570 <= not w3180 and not w3183;
w3571 <= not w554 and w1466;
w3572 <= not w444 and w3161;
w3573 <= not w446 and w3572;
w3574 <= not w997 and w3573;
w3575 <= not w591 and w3574;
w3576 <= not w84 and w3575;
w3577 <= not w302 and w3576;
w3578 <= not w180 and w3577;
w3579 <= not w16 and w3578;
w3580 <= not w67 and not w98;
w3581 <= w137 and w3580;
w3582 <= not w492 and w3581;
w3583 <= not w288 and w3582;
w3584 <= not w110 and w3583;
w3585 <= not w178 and w3584;
w3586 <= not w504 and w3585;
w3587 <= w1343 and w1393;
w3588 <= w3407 and w3587;
w3589 <= w3187 and w3588;
w3590 <= not w333 and w3589;
w3591 <= not w167 and w3590;
w3592 <= not w106 and w3591;
w3593 <= not w234 and w3592;
w3594 <= not w292 and w3593;
w3595 <= not w309 and w3594;
w3596 <= not w303 and w3595;
w3597 <= not w30 and w3596;
w3598 <= not w568 and w3597;
w3599 <= w3586 and w3598;
w3600 <= w2516 and w3599;
w3601 <= w3579 and w3600;
w3602 <= w176 and w3601;
w3603 <= not w71 and w3602;
w3604 <= w3571 and w3603;
w3605 <= not w360 and w3604;
w3606 <= not w209 and w3605;
w3607 <= not w401 and w3606;
w3608 <= not w357 and w3607;
w3609 <= not w273 and w3608;
w3610 <= not w590 and w3609;
w3611 <= not w164 and not w1007;
w3612 <= not w210 and w3611;
w3613 <= not w396 and w3612;
w3614 <= not w351 and w3613;
w3615 <= not w1138 and w3614;
w3616 <= not w187 and w3615;
w3617 <= not w439 and not w576;
w3618 <= not w241 and w3617;
w3619 <= not w207 and w3618;
w3620 <= not w157 and w3619;
w3621 <= not w428 and w1315;
w3622 <= not w945 and w3621;
w3623 <= w2362 and w3622;
w3624 <= w658 and w3623;
w3625 <= w3620 and w3624;
w3626 <= w1258 and w3625;
w3627 <= w3616 and w3626;
w3628 <= w3610 and w3627;
w3629 <= w1850 and w3628;
w3630 <= w981 and w3629;
w3631 <= w1301 and w3630;
w3632 <= not w104 and w3631;
w3633 <= not w782 and w3632;
w3634 <= not w86 and w3633;
w3635 <= not w53 and w3634;
w3636 <= not w141 and w3635;
w3637 <= not w387 and w3636;
w3638 <= w3018 and not w3637;
w3639 <= not w3018 and w3637;
w3640 <= not w3570 and not w3639;
w3641 <= not w3638 and w3640;
w3642 <= not w3570 and not w3641;
w3643 <= not w3639 and not w3641;
w3644 <= not w3638 and w3643;
w3645 <= not w3642 and not w3644;
w3646 <= w2955 and not w3474;
w3647 <= not w2947 and w2963;
w3648 <= not w327 and w2958;
w3649 <= w3548 and not w3550;
w3650 <= not w3551 and not w3649;
w3651 <= w10 and w3650;
w3652 <= not w3648 and not w3651;
w3653 <= not w3647 and w3652;
w3654 <= not w3646 and w3653;
w3655 <= not w3645 and not w3654;
w3656 <= not w3645 and not w3655;
w3657 <= not w3654 and not w3655;
w3658 <= not w3656 and not w3657;
w3659 <= not w3569 and not w3658;
w3660 <= not w3569 and not w3659;
w3661 <= not w3658 and not w3659;
w3662 <= not w3660 and not w3661;
w3663 <= not w124 and not w215;
w3664 <= not w50 and w3663;
w3665 <= not w104 and w3664;
w3666 <= not w84 and w3665;
w3667 <= not w425 and w3666;
w3668 <= not w502 and w3667;
w3669 <= not w493 and w1774;
w3670 <= not w602 and w3669;
w3671 <= not w687 and w3670;
w3672 <= not w492 and w3671;
w3673 <= not w158 and w3672;
w3674 <= not w558 and w3673;
w3675 <= w575 and w830;
w3676 <= not w58 and w3675;
w3677 <= not w85 and w3676;
w3678 <= not w166 and w3677;
w3679 <= w336 and w2491;
w3680 <= w3678 and w3679;
w3681 <= w3674 and w3680;
w3682 <= w3668 and w3681;
w3683 <= w2517 and w3682;
w3684 <= w655 and w3683;
w3685 <= w1076 and w3684;
w3686 <= w450 and w3685;
w3687 <= w1302 and w3686;
w3688 <= not w738 and w3687;
w3689 <= not w446 and w3688;
w3690 <= not w112 and w3689;
w3691 <= not w82 and w3690;
w3692 <= not w360 and w3691;
w3693 <= not w555 and w2228;
w3694 <= not w140 and w3693;
w3695 <= not w96 and w3694;
w3696 <= not w409 and w3695;
w3697 <= not w275 and w3696;
w3698 <= not w371 and w3697;
w3699 <= not w499 and w3698;
w3700 <= w1327 and w3050;
w3701 <= w525 and w3700;
w3702 <= not w53 and w3701;
w3703 <= not w462 and w3702;
w3704 <= not w357 and w682;
w3705 <= not w945 and w3704;
w3706 <= not w504 and w3705;
w3707 <= w1719 and w3706;
w3708 <= w3703 and w3707;
w3709 <= w2447 and w3708;
w3710 <= w807 and w3709;
w3711 <= not w211 and w3710;
w3712 <= not w537 and w3711;
w3713 <= not w819 and w3712;
w3714 <= not w329 and w3713;
w3715 <= not w260 and w3714;
w3716 <= not w206 and w3715;
w3717 <= not w363 and w3716;
w3718 <= w1323 and w1512;
w3719 <= not w498 and w3718;
w3720 <= not w67 and w3719;
w3721 <= not w160 and w3720;
w3722 <= not w466 and w3721;
w3723 <= not w592 and w3722;
w3724 <= not w1039 and w3723;
w3725 <= not w21 and w3724;
w3726 <= not w79 and not w401;
w3727 <= not w126 and w3726;
w3728 <= w2975 and w3727;
w3729 <= w3725 and w3728;
w3730 <= w3717 and w3729;
w3731 <= w3699 and w3730;
w3732 <= w2675 and w3731;
w3733 <= w872 and w3732;
w3734 <= w3692 and w3733;
w3735 <= w1696 and w3734;
w3736 <= w473 and w3735;
w3737 <= not w397 and w3736;
w3738 <= not w337 and w3737;
w3739 <= not w212 and w3738;
w3740 <= not w228 and w3739;
w3741 <= w3392 and not w3740;
w3742 <= w3477 and not w3540;
w3743 <= not w3391 and w3541;
w3744 <= not w3742 and not w3743;
w3745 <= not w3741 and w3744;
w3746 <= not w3303 and w3745;
w3747 <= not w3557 and not w3560;
w3748 <= not w3391 and not w3740;
w3749 <= w3391 and w3740;
w3750 <= not w3748 and not w3749;
w3751 <= not w3747 and w3750;
w3752 <= w3747 and not w3750;
w3753 <= not w3751 and not w3752;
w3754 <= w3745 and not w3753;
w3755 <= not w3746 and not w3754;
w3756 <= a(29) and not w3755;
w3757 <= not a(29) and w3755;
w3758 <= not w3756 and not w3757;
w3759 <= w3662 and w3758;
w3760 <= not w3662 and not w3758;
w3761 <= not w3759 and not w3760;
w3762 <= not w221 and not w373;
w3763 <= w3372 and w3762;
w3764 <= not w180 and w3763;
w3765 <= not w726 and w3764;
w3766 <= not w357 and w3765;
w3767 <= not w233 and not w896;
w3768 <= w3766 and w3767;
w3769 <= w600 and w3768;
w3770 <= w474 and w3769;
w3771 <= w389 and w3770;
w3772 <= w128 and w3771;
w3773 <= not w34 and w3772;
w3774 <= not w307 and w3773;
w3775 <= w707 and w1040;
w3776 <= w406 and w3775;
w3777 <= w762 and w3776;
w3778 <= not w592 and w3777;
w3779 <= not w187 and w3778;
w3780 <= not w527 and w3779;
w3781 <= not w212 and w3780;
w3782 <= not w267 and w3781;
w3783 <= not w1062 and w3782;
w3784 <= w2143 and w2508;
w3785 <= w63 and w3784;
w3786 <= not w424 and w3785;
w3787 <= not w54 and w3786;
w3788 <= w2210 and w3787;
w3789 <= w3783 and w3788;
w3790 <= not w21 and w3789;
w3791 <= not w504 and w3790;
w3792 <= not w364 and w525;
w3793 <= not w166 and w3792;
w3794 <= w559 and w3141;
w3795 <= w2898 and w3794;
w3796 <= w1189 and w3795;
w3797 <= w914 and w3796;
w3798 <= w291 and w3797;
w3799 <= not w224 and w3798;
w3800 <= not w219 and w3799;
w3801 <= not w492 and w3800;
w3802 <= w3793 and w3801;
w3803 <= not w568 and w3802;
w3804 <= not w205 and w3803;
w3805 <= w3505 and w3804;
w3806 <= w1415 and w3805;
w3807 <= w903 and w3806;
w3808 <= not w384 and w3807;
w3809 <= w3791 and w3808;
w3810 <= w3774 and w3809;
w3811 <= not w263 and w3810;
w3812 <= not w231 and w3811;
w3813 <= a(23) and not a(24);
w3814 <= not a(23) and a(24);
w3815 <= not w3813 and not w3814;
w3816 <= a(25) and not a(26);
w3817 <= not a(25) and a(26);
w3818 <= not w3816 and not w3817;
w3819 <= not w3815 and w3818;
w3820 <= not w3812 and w3819;
w3821 <= not w62 and not w212;
w3822 <= w2325 and w2976;
w3823 <= w2568 and w3822;
w3824 <= w1414 and w3823;
w3825 <= w1759 and w3824;
w3826 <= w3821 and w3825;
w3827 <= not w125 and w3826;
w3828 <= not w782 and w3827;
w3829 <= not w712 and w3828;
w3830 <= not w427 and w3829;
w3831 <= not w98 and w3830;
w3832 <= not w105 and w3831;
w3833 <= not w275 and w3832;
w3834 <= not w607 and w3833;
w3835 <= not w371 and w3834;
w3836 <= not w293 and w3835;
w3837 <= not w46 and not w440;
w3838 <= not w329 and w3837;
w3839 <= not w310 and w3838;
w3840 <= not w818 and w3839;
w3841 <= w682 and w913;
w3842 <= not w171 and not w236;
w3843 <= not w71 and w3842;
w3844 <= not w404 and w3843;
w3845 <= not w1241 and w3844;
w3846 <= not w332 and w3845;
w3847 <= not w333 and w3846;
w3848 <= w710 and w3847;
w3849 <= not w1007 and w3848;
w3850 <= w452 and w3849;
w3851 <= w3841 and w3850;
w3852 <= w667 and w3851;
w3853 <= w3840 and w3852;
w3854 <= w3836 and w3853;
w3855 <= w1666 and w3854;
w3856 <= not w552 and w3855;
w3857 <= not w425 and w3856;
w3858 <= not w360 and w3857;
w3859 <= not w403 and w3858;
w3860 <= not w208 and w3859;
w3861 <= not w230 and w3860;
w3862 <= not w467 and w3861;
w3863 <= not w821 and w3862;
w3864 <= not w504 and w3863;
w3865 <= not w265 and w2673;
w3866 <= not w177 and w3865;
w3867 <= w2633 and w3866;
w3868 <= not w439 and w3867;
w3869 <= not w180 and w3868;
w3870 <= not w77 and w3869;
w3871 <= not w726 and w3870;
w3872 <= not w502 and w3871;
w3873 <= not w206 and w3872;
w3874 <= not w706 and w3873;
w3875 <= w1375 and w3664;
w3876 <= w3344 and w3875;
w3877 <= w1227 and w3876;
w3878 <= not w211 and w3877;
w3879 <= not w103 and w3878;
w3880 <= not w361 and w3879;
w3881 <= not w1037 and w3880;
w3882 <= not w446 and w3881;
w3883 <= not w307 and w1415;
w3884 <= not w384 and w3883;
w3885 <= w1090 and w3884;
w3886 <= w3882 and w3885;
w3887 <= w2675 and w3886;
w3888 <= w3874 and w3887;
w3889 <= w3864 and w3888;
w3890 <= w981 and w3889;
w3891 <= w455 and w3890;
w3892 <= w2518 and w3891;
w3893 <= w655 and w3892;
w3894 <= not w946 and w3893;
w3895 <= not w915 and w3894;
w3896 <= not w387 and w3895;
w3897 <= not w471 and w3896;
w3898 <= not w218 and w3897;
w3899 <= not w273 and w3898;
w3900 <= not w11 and not w19;
w3901 <= w3815 and not w3818;
w3902 <= not w3900 and w3901;
w3903 <= not w3899 and w3902;
w3904 <= not w427 and not w431;
w3905 <= not w365 and w3904;
w3906 <= not w440 and w3905;
w3907 <= not w360 and w3906;
w3908 <= w2405 and w3767;
w3909 <= not w554 and w3908;
w3910 <= not w172 and w3909;
w3911 <= not w647 and w3910;
w3912 <= not w386 and w3911;
w3913 <= not w527 and w3912;
w3914 <= w1413 and w1661;
w3915 <= not w262 and w3914;
w3916 <= not w26 and w3915;
w3917 <= not w650 and w3916;
w3918 <= not w37 and w3917;
w3919 <= not w222 and w3918;
w3920 <= not w225 and not w819;
w3921 <= not w82 and w3920;
w3922 <= not w338 and w3921;
w3923 <= w1282 and w3922;
w3924 <= not w90 and w3923;
w3925 <= not w331 and w3924;
w3926 <= w1851 and w2232;
w3927 <= not w84 and w3926;
w3928 <= not w529 and w3927;
w3929 <= not w158 and w3928;
w3930 <= not w337 and w3929;
w3931 <= not w240 and w3930;
w3932 <= not w161 and w3931;
w3933 <= w3925 and w3932;
w3934 <= w473 and w3933;
w3935 <= not w370 and w3934;
w3936 <= not w227 and w3935;
w3937 <= not w218 and w3936;
w3938 <= not w307 and w3937;
w3939 <= w2068 and w2638;
w3940 <= w2674 and w3939;
w3941 <= w1183 and w3940;
w3942 <= w1324 and w3941;
w3943 <= not w441 and w3942;
w3944 <= not w42 and w3943;
w3945 <= not w210 and w2928;
w3946 <= not w352 and w3945;
w3947 <= w3343 and w3946;
w3948 <= w3944 and w3947;
w3949 <= w3938 and w3948;
w3950 <= w1718 and w3949;
w3951 <= w356 and w3950;
w3952 <= not w388 and w3951;
w3953 <= w3849 and w3866;
w3954 <= w3063 and w3953;
w3955 <= w3882 and w3954;
w3956 <= not w58 and w3955;
w3957 <= not w129 and w3956;
w3958 <= not w46 and w3957;
w3959 <= not w681 and w3958;
w3960 <= not w397 and w3959;
w3961 <= not w444 and w3960;
w3962 <= not w946 and w3961;
w3963 <= not w125 and w3962;
w3964 <= not w453 and w3963;
w3965 <= not w86 and w3964;
w3966 <= w3952 and w3965;
w3967 <= w3919 and w3966;
w3968 <= not w760 and w3967;
w3969 <= not w34 and w3968;
w3970 <= w1139 and w3787;
w3971 <= w3725 and w3970;
w3972 <= w539 and w3971;
w3973 <= w981 and w3972;
w3974 <= w94 and w3973;
w3975 <= not w65 and w3974;
w3976 <= w3969 and w3975;
w3977 <= w3913 and w3976;
w3978 <= w3907 and w3977;
w3979 <= w406 and w3978;
w3980 <= not w524 and w3979;
w3981 <= w3815 and w3900;
w3982 <= not w3980 and w3981;
w3983 <= not w3903 and not w3982;
w3984 <= not w3820 and w3983;
w3985 <= not w3815 and not w3818;
w3986 <= not w3899 and not w3980;
w3987 <= not w3740 and not w3899;
w3988 <= not w3748 and not w3751;
w3989 <= w3740 and w3899;
w3990 <= not w3987 and not w3989;
w3991 <= not w3988 and w3990;
w3992 <= not w3987 and not w3991;
w3993 <= w3899 and w3980;
w3994 <= not w3986 and not w3993;
w3995 <= not w3992 and w3994;
w3996 <= not w3986 and not w3995;
w3997 <= not w3812 and not w3980;
w3998 <= w3812 and w3980;
w3999 <= not w3997 and not w3998;
w4000 <= not w3996 and w3999;
w4001 <= w3996 and not w3999;
w4002 <= not w4000 and not w4001;
w4003 <= w3985 and w4002;
w4004 <= w3984 and not w4003;
w4005 <= a(26) and not w4004;
w4006 <= a(26) and not w4005;
w4007 <= not w4004 and not w4005;
w4008 <= not w4006 and not w4007;
w4009 <= w3761 and not w4008;
w4010 <= w3761 and not w4009;
w4011 <= not w4008 and not w4009;
w4012 <= not w4010 and not w4011;
w4013 <= w3392 and not w3540;
w4014 <= not w2947 and w3477;
w4015 <= not w3474 and w3541;
w4016 <= not w4014 and not w4015;
w4017 <= not w4013 and w4016;
w4018 <= w3552 and not w3554;
w4019 <= not w3555 and not w4018;
w4020 <= w3303 and w4019;
w4021 <= w4017 and not w4020;
w4022 <= a(29) and not w4021;
w4023 <= not w4021 and not w4022;
w4024 <= a(29) and not w4022;
w4025 <= not w4023 and not w4024;
w4026 <= not w3289 and not w3292;
w4027 <= w3291 and not w3292;
w4028 <= not w4026 and not w4027;
w4029 <= not w4025 and not w4028;
w4030 <= not w4025 and not w4029;
w4031 <= not w4028 and not w4029;
w4032 <= not w4030 and not w4031;
w4033 <= not w3273 and not w3275;
w4034 <= not w3264 and w3276;
w4035 <= not w4033 and not w4034;
w4036 <= not w330 and not w529;
w4037 <= not w289 and not w946;
w4038 <= not w112 and w4037;
w4039 <= not w302 and w4038;
w4040 <= w185 and w1695;
w4041 <= w727 and w4040;
w4042 <= w2127 and w4041;
w4043 <= w4039 and w4042;
w4044 <= w2878 and w4043;
w4045 <= w812 and w4044;
w4046 <= w2152 and w4045;
w4047 <= w3340 and w4046;
w4048 <= w3836 and w4047;
w4049 <= w2435 and w4048;
w4050 <= w1118 and w4049;
w4051 <= w442 and w4050;
w4052 <= w4036 and w4051;
w4053 <= not w262 and w4052;
w4054 <= not w227 and w4053;
w4055 <= not w221 and w4054;
w4056 <= not w1039 and w4055;
w4057 <= not w330 and w1008;
w4058 <= not w915 and w4057;
w4059 <= not w100 and w4058;
w4060 <= not w867 and w4059;
w4061 <= not w310 and w4060;
w4062 <= not w21 and w4061;
w4063 <= w1074 and w1716;
w4064 <= not w177 and w4063;
w4065 <= not w497 and w4064;
w4066 <= not w337 and w1116;
w4067 <= not w351 and w4066;
w4068 <= w980 and w4067;
w4069 <= w747 and w4068;
w4070 <= w1627 and w4069;
w4071 <= w4065 and w4070;
w4072 <= w4062 and w4071;
w4073 <= w426 and w4072;
w4074 <= w1186 and w4073;
w4075 <= w1076 and w4074;
w4076 <= not w58 and w4075;
w4077 <= not w269 and w4076;
w4078 <= not w1036 and w4077;
w4079 <= not w529 and w4078;
w4080 <= not w462 and w4079;
w4081 <= not w624 and w4080;
w4082 <= not w135 and w4081;
w4083 <= not w1039 and w4082;
w4084 <= not w103 and not w1138;
w4085 <= not w821 and w4084;
w4086 <= not w123 and w4085;
w4087 <= w214 and not w524;
w4088 <= not w329 and w4087;
w4089 <= w4086 and w4088;
w4090 <= w2306 and w4089;
w4091 <= w3456 and w4090;
w4092 <= w4083 and w4091;
w4093 <= w3343 and w4092;
w4094 <= w708 and w4093;
w4095 <= w170 and w4094;
w4096 <= w389 and w4095;
w4097 <= w975 and w4096;
w4098 <= not w332 and w4097;
w4099 <= not w289 and w4098;
w4100 <= not w1037 and w4099;
w4101 <= not w262 and w4100;
w4102 <= not w338 and w4101;
w4103 <= w1459 and w4102;
w4104 <= not w261 and w4103;
w4105 <= not w373 and w4104;
w4106 <= not w136 and w4105;
w4107 <= not w4056 and not w4106;
w4108 <= w4056 and w4106;
w4109 <= not w4107 and not w4108;
w4110 <= not a(17) and w4109;
w4111 <= not w4107 and not w4110;
w4112 <= w3081 and not w4111;
w4113 <= w2851 and not w2853;
w4114 <= not w2854 and not w4113;
w4115 <= w10 and w4114;
w4116 <= not w645 and w2955;
w4117 <= not w893 and w2958;
w4118 <= not w802 and w2963;
w4119 <= not w4117 and not w4118;
w4120 <= not w4116 and w4119;
w4121 <= not w4115 and w4120;
w4122 <= not w3081 and w4111;
w4123 <= not w4112 and not w4122;
w4124 <= not w4121 and w4123;
w4125 <= not w4112 and not w4124;
w4126 <= not w4035 and not w4125;
w4127 <= w4035 and w4125;
w4128 <= not w4126 and not w4127;
w4129 <= not w4121 and not w4124;
w4130 <= w4123 and not w4124;
w4131 <= not w4129 and not w4130;
w4132 <= not a(17) and not w4110;
w4133 <= not w4108 and w4111;
w4134 <= not w4132 and not w4133;
w4135 <= not w802 and w2955;
w4136 <= not w893 and w2963;
w4137 <= not w995 and w2958;
w4138 <= w2847 and not w2849;
w4139 <= not w2850 and not w4138;
w4140 <= w10 and w4139;
w4141 <= not w4137 and not w4140;
w4142 <= not w4136 and w4141;
w4143 <= not w4135 and w4142;
w4144 <= not w4134 and not w4143;
w4145 <= w2283 and w2450;
w4146 <= w912 and w4145;
w4147 <= w2025 and w4146;
w4148 <= not w30 and w4147;
w4149 <= not w298 and w4148;
w4150 <= not w384 and w4149;
w4151 <= not w331 and not w365;
w4152 <= not w171 and not w1062;
w4153 <= not w810 and w4152;
w4154 <= w3020 and w4153;
w4155 <= w4151 and w4154;
w4156 <= w2067 and w4155;
w4157 <= w2236 and w4156;
w4158 <= w2137 and w4157;
w4159 <= w740 and w4158;
w4160 <= w334 and w4159;
w4161 <= w162 and w4160;
w4162 <= w820 and w4161;
w4163 <= not w71 and w4162;
w4164 <= not w602 and w4163;
w4165 <= not w1037 and w4164;
w4166 <= not w124 and w4165;
w4167 <= not w647 and w4166;
w4168 <= not w431 and w2403;
w4169 <= not w818 and w4168;
w4170 <= w3762 and w4169;
w4171 <= w713 and w4170;
w4172 <= w1952 and w4171;
w4173 <= w2675 and w4172;
w4174 <= w91 and w4173;
w4175 <= not w58 and w4174;
w4176 <= not w288 and w4175;
w4177 <= not w50 and w4176;
w4178 <= not w168 and w4177;
w4179 <= not w574 and w4178;
w4180 <= not w360 and w4179;
w4181 <= not w34 and w4180;
w4182 <= not w241 and w4181;
w4183 <= w476 and w2176;
w4184 <= w2265 and w4183;
w4185 <= w2442 and w4184;
w4186 <= w4182 and w4185;
w4187 <= w4167 and w4186;
w4188 <= w4150 and w4187;
w4189 <= w2570 and w4188;
w4190 <= w2617 and w4189;
w4191 <= w1716 and w4190;
w4192 <= not w362 and w4191;
w4193 <= not w396 and w4192;
w4194 <= not w163 and w4193;
w4195 <= not w261 and w4194;
w4196 <= not w330 and w4195;
w4197 <= not w649 and w4196;
w4198 <= not w239 and w4197;
w4199 <= not w601 and w4198;
w4200 <= not w821 and w4199;
w4201 <= not w706 and w4200;
w4202 <= w4056 and not w4201;
w4203 <= not w4056 and w4201;
w4204 <= not w85 and not w90;
w4205 <= w185 and w4204;
w4206 <= not w687 and w4205;
w4207 <= not w337 and w4206;
w4208 <= not w365 and w4207;
w4209 <= not w363 and w4208;
w4210 <= not w211 and not w354;
w4211 <= not w338 and w4210;
w4212 <= not w359 and w4211;
w4213 <= not w105 and w4212;
w4214 <= not w818 and w4213;
w4215 <= w1879 and w2619;
w4216 <= w4214 and w4215;
w4217 <= w4150 and w4216;
w4218 <= w4209 and w4217;
w4219 <= w1852 and w4218;
w4220 <= w708 and w4219;
w4221 <= w1172 and w4220;
w4222 <= not w213 and w4221;
w4223 <= not w240 and w4222;
w4224 <= not w81 and w4223;
w4225 <= not w37 and w4224;
w4226 <= not w867 and w4225;
w4227 <= not w135 and w4226;
w4228 <= not w306 and w4227;
w4229 <= not w274 and not w309;
w4230 <= not w273 and w4229;
w4231 <= not w34 and not w265;
w4232 <= not w92 and w4231;
w4233 <= not w405 and w4232;
w4234 <= w982 and w2572;
w4235 <= w4153 and w4234;
w4236 <= w4233 and w4235;
w4237 <= w3399 and w4236;
w4238 <= w2673 and w4237;
w4239 <= w4230 and w4238;
w4240 <= not w58 and w4239;
w4241 <= not w493 and w4240;
w4242 <= not w84 and w4241;
w4243 <= not w462 and w4242;
w4244 <= not w439 and w4243;
w4245 <= not w208 and w4244;
w4246 <= not w499 and w4245;
w4247 <= not w70 and not w387;
w4248 <= not w218 and w4247;
w4249 <= w876 and w4248;
w4250 <= w1537 and w4249;
w4251 <= not w89 and w4250;
w4252 <= not w554 and w4251;
w4253 <= not w56 and w4252;
w4254 <= not w529 and w4253;
w4255 <= not w331 and w4254;
w4256 <= not w712 and w4255;
w4257 <= not w261 and w4256;
w4258 <= not w360 and w4257;
w4259 <= not w233 and w4258;
w4260 <= not w726 and w4259;
w4261 <= not w209 and not w361;
w4262 <= not w568 and w4261;
w4263 <= w2306 and w4262;
w4264 <= w2008 and w4263;
w4265 <= not w446 and w4264;
w4266 <= not w591 and w4265;
w4267 <= not w592 and w4266;
w4268 <= not w127 and not w444;
w4269 <= not w275 and w4268;
w4270 <= not w168 and not w650;
w4271 <= w3049 and w4270;
w4272 <= w4269 and w4271;
w4273 <= w4267 and w4272;
w4274 <= w2675 and w4273;
w4275 <= w2104 and w4274;
w4276 <= w4260 and w4275;
w4277 <= w4246 and w4276;
w4278 <= w4228 and w4277;
w4279 <= w426 and w4278;
w4280 <= w1117 and w4279;
w4281 <= not w53 and w4280;
w4282 <= not w624 and w4281;
w4283 <= not w212 and w4282;
w4284 <= not w607 and w4283;
w4285 <= not w21 and w4284;
w4286 <= not w123 and w4285;
w4287 <= not w1181 and w1604;
w4288 <= not w224 and w4287;
w4289 <= not w396 and w4288;
w4290 <= not w298 and w4289;
w4291 <= not w497 and w4290;
w4292 <= not w608 and not w1241;
w4293 <= w1070 and w2269;
w4294 <= w4292 and w4293;
w4295 <= w975 and w4294;
w4296 <= not w167 and w4295;
w4297 <= not w190 and w4296;
w4298 <= not w138 and w4297;
w4299 <= not w744 and w4298;
w4300 <= not w174 and w4299;
w4301 <= not w307 and w4300;
w4302 <= not w37 and not w228;
w4303 <= w811 and w2145;
w4304 <= w4088 and w4303;
w4305 <= w1948 and w4304;
w4306 <= w2742 and w4305;
w4307 <= w4302 and w4306;
w4308 <= not w104 and w4307;
w4309 <= not w125 and w4308;
w4310 <= not w370 and w4309;
w4311 <= w1207 and w4169;
w4312 <= w374 and w4311;
w4313 <= w4310 and w4312;
w4314 <= w3313 and w4313;
w4315 <= w1485 and w4314;
w4316 <= not w362 and w4315;
w4317 <= not w355 and w4316;
w4318 <= not w81 and w4317;
w4319 <= not w231 and w4318;
w4320 <= not w915 and w4319;
w4321 <= not w136 and w4320;
w4322 <= not w206 and w4321;
w4323 <= not w184 and w4322;
w4324 <= w728 and w3231;
w4325 <= w2231 and w4324;
w4326 <= w550 and w4325;
w4327 <= w1265 and w4326;
w4328 <= w762 and w4327;
w4329 <= w913 and w4328;
w4330 <= w525 and w4329;
w4331 <= not w602 and w4330;
w4332 <= not w290 and w4331;
w4333 <= not w87 and w4332;
w4334 <= not w446 and w4333;
w4335 <= not w529 and w4334;
w4336 <= not w572 and w4335;
w4337 <= not w42 and w4336;
w4338 <= not w536 and w4337;
w4339 <= not w538 and w4338;
w4340 <= not w273 and w4339;
w4341 <= w1949 and w3351;
w4342 <= w1281 and w4341;
w4343 <= w927 and w4342;
w4344 <= w1720 and w4343;
w4345 <= w4340 and w4344;
w4346 <= w4323 and w4345;
w4347 <= w4301 and w4346;
w4348 <= w4291 and w4347;
w4349 <= w709 and w4348;
w4350 <= w2633 and w4349;
w4351 <= w220 and w4350;
w4352 <= not w171 and w4351;
w4353 <= not w332 and w4352;
w4354 <= not w270 and w4353;
w4355 <= not w498 and w4354;
w4356 <= not w424 and w4355;
w4357 <= not w4286 and not w4356;
w4358 <= w4286 and w4356;
w4359 <= not w4357 and not w4358;
w4360 <= not a(14) and w4359;
w4361 <= not w4357 and not w4360;
w4362 <= w4201 and not w4361;
w4363 <= w2839 and not w2841;
w4364 <= not w2842 and not w4363;
w4365 <= w10 and w4364;
w4366 <= not w995 and w2955;
w4367 <= not w1170 and w2958;
w4368 <= not w1113 and w2963;
w4369 <= not w4367 and not w4368;
w4370 <= not w4366 and w4369;
w4371 <= not w4365 and w4370;
w4372 <= not w4201 and w4361;
w4373 <= not w4362 and not w4372;
w4374 <= not w4371 and w4373;
w4375 <= not w4362 and not w4374;
w4376 <= not w4202 and not w4375;
w4377 <= not w4203 and w4376;
w4378 <= not w4202 and not w4377;
w4379 <= w4134 and w4143;
w4380 <= not w4144 and not w4379;
w4381 <= not w4378 and w4380;
w4382 <= not w4144 and not w4381;
w4383 <= not w4131 and not w4382;
w4384 <= w4131 and w4382;
w4385 <= not w4383 and not w4384;
w4386 <= not w2947 and w3392;
w4387 <= not w522 and w3477;
w4388 <= not w327 and w3541;
w4389 <= not w4387 and not w4388;
w4390 <= not w4386 and w4389;
w4391 <= not w3303 and w4390;
w4392 <= not w2953 and w4390;
w4393 <= not w4391 and not w4392;
w4394 <= a(29) and not w4393;
w4395 <= not a(29) and w4393;
w4396 <= not w4394 and not w4395;
w4397 <= w4385 and not w4396;
w4398 <= not w4383 and not w4397;
w4399 <= w4128 and not w4398;
w4400 <= not w4126 and not w4399;
w4401 <= not w4032 and not w4400;
w4402 <= not w4029 and not w4401;
w4403 <= not w3296 and w3567;
w4404 <= not w3568 and not w4403;
w4405 <= not w4402 and w4404;
w4406 <= w3819 and not w3980;
w4407 <= not w3740 and w3902;
w4408 <= not w3899 and w3981;
w4409 <= not w4407 and not w4408;
w4410 <= not w4406 and w4409;
w4411 <= w3992 and not w3994;
w4412 <= not w3995 and not w4411;
w4413 <= w3985 and w4412;
w4414 <= w4410 and not w4413;
w4415 <= a(26) and not w4414;
w4416 <= not w4414 and not w4415;
w4417 <= a(26) and not w4415;
w4418 <= not w4416 and not w4417;
w4419 <= not w4402 and not w4405;
w4420 <= w4404 and not w4405;
w4421 <= not w4419 and not w4420;
w4422 <= not w4418 and not w4421;
w4423 <= not w4405 and not w4422;
w4424 <= not w649 and w1949;
w4425 <= not w178 and w4424;
w4426 <= not w80 and w4425;
w4427 <= not w401 and w4426;
w4428 <= not w140 and w4427;
w4429 <= w1323 and w1720;
w4430 <= w539 and w4429;
w4431 <= w2105 and w4430;
w4432 <= not w108 and w4431;
w4433 <= not w79 and w4432;
w4434 <= not w329 and w4433;
w4435 <= not w241 and w4434;
w4436 <= not w92 and w4435;
w4437 <= not w310 and w4436;
w4438 <= w68 and w4437;
w4439 <= w4428 and w4438;
w4440 <= w2281 and w4439;
w4441 <= w981 and w4440;
w4442 <= w1696 and w4441;
w4443 <= w1302 and w4442;
w4444 <= not w209 and w4443;
w4445 <= not w524 and w4444;
w4446 <= not w403 and w4445;
w4447 <= w3907 and w4446;
w4448 <= not w231 and w4447;
w4449 <= not w536 and w4448;
w4450 <= w3774 and w4449;
w4451 <= not w3997 and not w4000;
w4452 <= not w3812 and not w4450;
w4453 <= w3812 and w4450;
w4454 <= not w4452 and not w4453;
w4455 <= not w4451 and w4454;
w4456 <= w3812 and not w4455;
w4457 <= not w4450 and not w4456;
w4458 <= not a(21) and a(22);
w4459 <= a(21) and not a(22);
w4460 <= not w4458 and not w4459;
w4461 <= a(20) and not a(21);
w4462 <= not a(20) and a(21);
w4463 <= not w4461 and not w4462;
w4464 <= not a(22) and a(23);
w4465 <= a(22) and not a(23);
w4466 <= not w4464 and not w4465;
w4467 <= w4463 and not w4466;
w4468 <= w4460 and w4467;
w4469 <= not w4450 and w4468;
w4470 <= not w4457 and not w4469;
w4471 <= not w4463 and not w4466;
w4472 <= not w4469 and not w4471;
w4473 <= not w4470 and not w4472;
w4474 <= a(23) and not w4473;
w4475 <= not a(23) and w4473;
w4476 <= not w4474 and not w4475;
w4477 <= not w4423 and not w4476;
w4478 <= w4423 and w4476;
w4479 <= not w4477 and not w4478;
w4480 <= not w4012 and w4479;
w4481 <= not w4012 and not w4480;
w4482 <= w4479 and not w4480;
w4483 <= not w4481 and not w4482;
w4484 <= w4032 and w4400;
w4485 <= not w4401 and not w4484;
w4486 <= w3819 and not w3899;
w4487 <= not w3391 and w3902;
w4488 <= not w3740 and w3981;
w4489 <= not w4487 and not w4488;
w4490 <= not w4486 and w4489;
w4491 <= not w3985 and w4490;
w4492 <= w3988 and not w3990;
w4493 <= not w3991 and not w4492;
w4494 <= w4490 and not w4493;
w4495 <= not w4491 and not w4494;
w4496 <= a(26) and not w4495;
w4497 <= not a(26) and w4495;
w4498 <= not w4496 and not w4497;
w4499 <= w4485 and not w4498;
w4500 <= not w3740 and w3819;
w4501 <= not w3540 and w3902;
w4502 <= not w3391 and w3981;
w4503 <= not w4501 and not w4502;
w4504 <= not w4500 and w4503;
w4505 <= w3753 and w3985;
w4506 <= w4504 and not w4505;
w4507 <= a(26) and not w4506;
w4508 <= a(26) and not w4507;
w4509 <= not w4506 and not w4507;
w4510 <= not w4508 and not w4509;
w4511 <= not w4128 and w4398;
w4512 <= not w4399 and not w4511;
w4513 <= w3392 and not w3474;
w4514 <= not w327 and w3477;
w4515 <= not w2947 and w3541;
w4516 <= not w4514 and not w4515;
w4517 <= not w4513 and w4516;
w4518 <= not w3303 and w4517;
w4519 <= not w3650 and w4517;
w4520 <= not w4518 and not w4519;
w4521 <= a(29) and not w4520;
w4522 <= not a(29) and w4520;
w4523 <= not w4521 and not w4522;
w4524 <= w4512 and not w4523;
w4525 <= not w4512 and w4523;
w4526 <= not w4524 and not w4525;
w4527 <= not w4510 and w4526;
w4528 <= not w4524 and not w4527;
w4529 <= w4485 and not w4499;
w4530 <= not w4498 and not w4499;
w4531 <= not w4529 and not w4530;
w4532 <= not w4528 and not w4531;
w4533 <= not w4499 and not w4532;
w4534 <= w4418 and not w4420;
w4535 <= not w4419 and w4534;
w4536 <= not w4422 and not w4535;
w4537 <= not w4533 and w4536;
w4538 <= not w3812 and w4468;
w4539 <= not w4460 and w4463;
w4540 <= not w4450 and w4539;
w4541 <= not w4538 and not w4540;
w4542 <= not w4452 and not w4455;
w4543 <= w4450 and w4542;
w4544 <= not w4457 and not w4543;
w4545 <= w4471 and w4544;
w4546 <= w4541 and not w4545;
w4547 <= a(23) and not w4546;
w4548 <= not w4546 and not w4547;
w4549 <= a(23) and not w4547;
w4550 <= not w4548 and not w4549;
w4551 <= w4533 and not w4536;
w4552 <= not w4537 and not w4551;
w4553 <= not w4550 and w4552;
w4554 <= not w4537 and not w4553;
w4555 <= w4483 and w4554;
w4556 <= not w4483 and not w4554;
w4557 <= not w4555 and not w4556;
w4558 <= w4526 and not w4527;
w4559 <= not w4510 and not w4527;
w4560 <= not w4558 and not w4559;
w4561 <= not w4375 and not w4377;
w4562 <= not w4203 and w4378;
w4563 <= not w4561 and not w4562;
w4564 <= not w893 and w2955;
w4565 <= not w995 and w2963;
w4566 <= not w1113 and w2958;
w4567 <= w2843 and not w2845;
w4568 <= not w2846 and not w4567;
w4569 <= w10 and w4568;
w4570 <= not w4566 and not w4569;
w4571 <= not w4565 and w4570;
w4572 <= not w4564 and w4571;
w4573 <= not w4563 and not w4572;
w4574 <= not w522 and w3392;
w4575 <= not w802 and w3477;
w4576 <= not w645 and w3541;
w4577 <= not w4575 and not w4576;
w4578 <= not w4574 and w4577;
w4579 <= w3266 and w3303;
w4580 <= w4578 and not w4579;
w4581 <= a(29) and not w4580;
w4582 <= not w4580 and not w4581;
w4583 <= a(29) and not w4581;
w4584 <= not w4582 and not w4583;
w4585 <= not w4563 and not w4573;
w4586 <= not w4572 and not w4573;
w4587 <= not w4585 and not w4586;
w4588 <= not w4584 and not w4587;
w4589 <= not w4573 and not w4588;
w4590 <= w4378 and not w4380;
w4591 <= not w4381 and not w4590;
w4592 <= not w4589 and w4591;
w4593 <= not w327 and w3392;
w4594 <= not w645 and w3477;
w4595 <= not w522 and w3541;
w4596 <= not w4594 and not w4595;
w4597 <= not w4593 and w4596;
w4598 <= w3282 and w3303;
w4599 <= w4597 and not w4598;
w4600 <= a(29) and not w4599;
w4601 <= a(29) and not w4600;
w4602 <= not w4599 and not w4600;
w4603 <= not w4601 and not w4602;
w4604 <= w4589 and not w4591;
w4605 <= not w4592 and not w4604;
w4606 <= not w4603 and w4605;
w4607 <= not w4592 and not w4606;
w4608 <= not w4385 and w4396;
w4609 <= not w4397 and not w4608;
w4610 <= not w4607 and w4609;
w4611 <= w4607 and not w4609;
w4612 <= not w4610 and not w4611;
w4613 <= not w3391 and w3819;
w4614 <= not w3474 and w3902;
w4615 <= not w3540 and w3981;
w4616 <= not w4614 and not w4615;
w4617 <= not w4613 and w4616;
w4618 <= w3562 and w3985;
w4619 <= w4617 and not w4618;
w4620 <= a(26) and not w4619;
w4621 <= a(26) and not w4620;
w4622 <= not w4619 and not w4620;
w4623 <= not w4621 and not w4622;
w4624 <= w4612 and not w4623;
w4625 <= not w4610 and not w4624;
w4626 <= not w4560 and not w4625;
w4627 <= w4560 and w4625;
w4628 <= not w4626 and not w4627;
w4629 <= not w4463 and w4466;
w4630 <= not w3812 and w4629;
w4631 <= not w3899 and w4468;
w4632 <= not w3980 and w4539;
w4633 <= not w4631 and not w4632;
w4634 <= not w4630 and w4633;
w4635 <= w4002 and w4471;
w4636 <= w4634 and not w4635;
w4637 <= a(23) and not w4636;
w4638 <= a(23) and not w4637;
w4639 <= not w4636 and not w4637;
w4640 <= not w4638 and not w4639;
w4641 <= w4628 and not w4640;
w4642 <= not w4626 and not w4641;
w4643 <= not w4450 and w4629;
w4644 <= not w3980 and w4468;
w4645 <= not w3812 and w4539;
w4646 <= not w4644 and not w4645;
w4647 <= not w4643 and w4646;
w4648 <= not w4471 and w4647;
w4649 <= w4451 and not w4454;
w4650 <= not w4455 and not w4649;
w4651 <= w4647 and not w4650;
w4652 <= not w4648 and not w4651;
w4653 <= a(23) and not w4652;
w4654 <= not a(23) and w4652;
w4655 <= not w4653 and not w4654;
w4656 <= not w4642 and not w4655;
w4657 <= w4642 and w4655;
w4658 <= not w4656 and not w4657;
w4659 <= not w4528 and not w4532;
w4660 <= not w4531 and not w4532;
w4661 <= not w4659 and not w4660;
w4662 <= w4658 and not w4661;
w4663 <= not w4656 and not w4662;
w4664 <= w4550 and not w4552;
w4665 <= not w4553 and not w4664;
w4666 <= not w4663 and w4665;
w4667 <= w4658 and not w4662;
w4668 <= not w4661 and not w4662;
w4669 <= not w4667 and not w4668;
w4670 <= w4612 and not w4624;
w4671 <= not w4623 and not w4624;
w4672 <= not w4670 and not w4671;
w4673 <= w4605 and not w4606;
w4674 <= not w4603 and not w4606;
w4675 <= not w4673 and not w4674;
w4676 <= not w3540 and w3819;
w4677 <= not w2947 and w3902;
w4678 <= not w3474 and w3981;
w4679 <= not w4677 and not w4678;
w4680 <= not w4676 and w4679;
w4681 <= not w3985 and w4680;
w4682 <= not w4019 and w4680;
w4683 <= not w4681 and not w4682;
w4684 <= a(26) and not w4683;
w4685 <= not a(26) and w4683;
w4686 <= not w4684 and not w4685;
w4687 <= not w4675 and not w4686;
w4688 <= not w4584 and not w4588;
w4689 <= not w4587 and not w4588;
w4690 <= not w4688 and not w4689;
w4691 <= not w4371 and not w4374;
w4692 <= w4373 and not w4374;
w4693 <= not w4691 and not w4692;
w4694 <= not a(14) and not w4360;
w4695 <= not w4358 and w4361;
w4696 <= not w4694 and not w4695;
w4697 <= not w552 and w2978;
w4698 <= not w89 and w4697;
w4699 <= not w576 and w4698;
w4700 <= not w263 and w4699;
w4701 <= not w329 and w4700;
w4702 <= not w601 and w4701;
w4703 <= not w499 and w3425;
w4704 <= not w821 and w4703;
w4705 <= w268 and w1324;
w4706 <= not w384 and w4705;
w4707 <= w2296 and w4706;
w4708 <= w4704 and w4707;
w4709 <= w76 and w4708;
w4710 <= w1116 and w4709;
w4711 <= w809 and w4710;
w4712 <= w903 and w4711;
w4713 <= w3187 and w4712;
w4714 <= w1762 and w4713;
w4715 <= w2518 and w4714;
w4716 <= w4036 and w4715;
w4717 <= not w104 and w4716;
w4718 <= not w221 and w4717;
w4719 <= not w524 and w4718;
w4720 <= not w187 and w4719;
w4721 <= not w270 and not w302;
w4722 <= not w310 and not w446;
w4723 <= not w239 and w4722;
w4724 <= w2089 and w4723;
w4725 <= not w1241 and w4724;
w4726 <= not w332 and w4725;
w4727 <= not w124 and w4726;
w4728 <= not w168 and w4727;
w4729 <= not w96 and w4728;
w4730 <= not w140 and not w210;
w4731 <= not w896 and w4730;
w4732 <= not w184 and w4731;
w4733 <= w1696 and w4302;
w4734 <= not w650 and w4733;
w4735 <= w4732 and w4734;
w4736 <= w232 and w4735;
w4737 <= w374 and w4736;
w4738 <= w4729 and w4737;
w4739 <= w4721 and w4738;
w4740 <= w868 and w4739;
w4741 <= w2154 and w4740;
w4742 <= w276 and w4741;
w4743 <= not w404 and w4742;
w4744 <= not w211 and w4743;
w4745 <= not w492 and w4744;
w4746 <= not w537 and w4745;
w4747 <= not w85 and w4746;
w4748 <= not w351 and w4747;
w4749 <= not w126 and w4748;
w4750 <= not w726 and w4749;
w4751 <= not w99 and not w493;
w4752 <= not w472 and w4751;
w4753 <= not w135 and w4752;
w4754 <= not w607 and w4753;
w4755 <= w2519 and w2656;
w4756 <= w4754 and w4755;
w4757 <= w1661 and w4756;
w4758 <= w505 and w4757;
w4759 <= not w946 and w4758;
w4760 <= not w225 and w4759;
w4761 <= not w181 and w4760;
w4762 <= not w328 and w4761;
w4763 <= not w431 and not w819;
w4764 <= w1908 and w4763;
w4765 <= w4762 and w4764;
w4766 <= w4750 and w4765;
w4767 <= w1863 and w4766;
w4768 <= w4720 and w4767;
w4769 <= w4702 and w4768;
w4770 <= w1511 and w4769;
w4771 <= w358 and w4770;
w4772 <= w2402 and w4771;
w4773 <= not w602 and w4772;
w4774 <= not w26 and w4773;
w4775 <= not w178 and w4774;
w4776 <= not w471 and w4775;
w4777 <= not w218 and w4776;
w4778 <= not w172 and w4777;
w4779 <= not w206 and w4778;
w4780 <= w4286 and not w4779;
w4781 <= not w4286 and w4779;
w4782 <= w2831 and not w2833;
w4783 <= not w2834 and not w4782;
w4784 <= w10 and w4783;
w4785 <= not w1170 and w2955;
w4786 <= not w1407 and w2958;
w4787 <= not w1299 and w2963;
w4788 <= not w4786 and not w4787;
w4789 <= not w4785 and w4788;
w4790 <= not w4784 and w4789;
w4791 <= not w4780 and not w4790;
w4792 <= not w4781 and w4791;
w4793 <= not w4780 and not w4792;
w4794 <= not w4696 and not w4793;
w4795 <= w2835 and not w2837;
w4796 <= not w2838 and not w4795;
w4797 <= w10 and w4796;
w4798 <= not w1113 and w2955;
w4799 <= not w1299 and w2958;
w4800 <= not w1170 and w2963;
w4801 <= not w4799 and not w4800;
w4802 <= not w4798 and w4801;
w4803 <= not w4797 and w4802;
w4804 <= w4696 and w4793;
w4805 <= not w4794 and not w4804;
w4806 <= not w4803 and w4805;
w4807 <= not w4794 and not w4806;
w4808 <= not w4693 and not w4807;
w4809 <= w4693 and w4807;
w4810 <= not w4808 and not w4809;
w4811 <= not w645 and w3392;
w4812 <= not w893 and w3477;
w4813 <= not w802 and w3541;
w4814 <= not w4812 and not w4813;
w4815 <= not w4811 and w4814;
w4816 <= not w3303 and w4815;
w4817 <= not w4114 and w4815;
w4818 <= not w4816 and not w4817;
w4819 <= a(29) and not w4818;
w4820 <= not a(29) and w4818;
w4821 <= not w4819 and not w4820;
w4822 <= w4810 and not w4821;
w4823 <= not w4808 and not w4822;
w4824 <= not w4690 and not w4823;
w4825 <= w4690 and w4823;
w4826 <= not w4824 and not w4825;
w4827 <= not w3474 and w3819;
w4828 <= not w327 and w3902;
w4829 <= not w2947 and w3981;
w4830 <= not w4828 and not w4829;
w4831 <= not w4827 and w4830;
w4832 <= w3650 and w3985;
w4833 <= w4831 and not w4832;
w4834 <= a(26) and not w4833;
w4835 <= a(26) and not w4834;
w4836 <= not w4833 and not w4834;
w4837 <= not w4835 and not w4836;
w4838 <= w4826 and not w4837;
w4839 <= not w4824 and not w4838;
w4840 <= w4675 and w4686;
w4841 <= not w4687 and not w4840;
w4842 <= not w4839 and w4841;
w4843 <= not w4687 and not w4842;
w4844 <= not w4672 and not w4843;
w4845 <= w4672 and w4843;
w4846 <= not w4844 and not w4845;
w4847 <= not w3980 and w4629;
w4848 <= not w3740 and w4468;
w4849 <= not w3899 and w4539;
w4850 <= not w4848 and not w4849;
w4851 <= not w4847 and w4850;
w4852 <= w4412 and w4471;
w4853 <= w4851 and not w4852;
w4854 <= a(23) and not w4853;
w4855 <= a(23) and not w4854;
w4856 <= not w4853 and not w4854;
w4857 <= not w4855 and not w4856;
w4858 <= w4846 and not w4857;
w4859 <= not w4844 and not w4858;
w4860 <= not a(18) and a(19);
w4861 <= a(18) and not a(19);
w4862 <= not w4860 and not w4861;
w4863 <= a(19) and not a(20);
w4864 <= not a(19) and a(20);
w4865 <= not w4863 and not w4864;
w4866 <= a(17) and not a(18);
w4867 <= not a(17) and a(18);
w4868 <= not w4866 and not w4867;
w4869 <= not w4865 and w4868;
w4870 <= w4862 and w4869;
w4871 <= not w4450 and w4870;
w4872 <= not w4457 and not w4871;
w4873 <= not w4865 and not w4868;
w4874 <= not w4871 and not w4873;
w4875 <= not w4872 and not w4874;
w4876 <= a(20) and not w4875;
w4877 <= not a(20) and w4875;
w4878 <= not w4876 and not w4877;
w4879 <= not w4859 and not w4878;
w4880 <= w4628 and not w4641;
w4881 <= not w4640 and not w4641;
w4882 <= not w4880 and not w4881;
w4883 <= w4859 and w4878;
w4884 <= not w4879 and not w4883;
w4885 <= not w4882 and w4884;
w4886 <= not w4879 and not w4885;
w4887 <= not w4669 and not w4886;
w4888 <= w4669 and w4886;
w4889 <= not w4887 and not w4888;
w4890 <= not w4882 and not w4885;
w4891 <= w4884 and not w4885;
w4892 <= not w4890 and not w4891;
w4893 <= w4846 and not w4858;
w4894 <= not w4857 and not w4858;
w4895 <= not w4893 and not w4894;
w4896 <= not w3899 and w4629;
w4897 <= not w3391 and w4468;
w4898 <= not w3740 and w4539;
w4899 <= not w4897 and not w4898;
w4900 <= not w4896 and w4899;
w4901 <= w4471 and w4493;
w4902 <= w4900 and not w4901;
w4903 <= a(23) and not w4902;
w4904 <= not w4902 and not w4903;
w4905 <= a(23) and not w4903;
w4906 <= not w4904 and not w4905;
w4907 <= w4839 and not w4841;
w4908 <= not w4842 and not w4907;
w4909 <= not w4906 and w4908;
w4910 <= not w4906 and not w4909;
w4911 <= w4908 and not w4909;
w4912 <= not w4910 and not w4911;
w4913 <= w4826 and not w4838;
w4914 <= not w4837 and not w4838;
w4915 <= not w4913 and not w4914;
w4916 <= not w802 and w3392;
w4917 <= not w995 and w3477;
w4918 <= not w893 and w3541;
w4919 <= not w4917 and not w4918;
w4920 <= not w4916 and w4919;
w4921 <= w3303 and w4139;
w4922 <= w4920 and not w4921;
w4923 <= a(29) and not w4922;
w4924 <= not w4922 and not w4923;
w4925 <= a(29) and not w4923;
w4926 <= not w4924 and not w4925;
w4927 <= not w4803 and not w4806;
w4928 <= w4805 and not w4806;
w4929 <= not w4927 and not w4928;
w4930 <= not w4926 and not w4929;
w4931 <= not w4926 and not w4930;
w4932 <= not w4929 and not w4930;
w4933 <= not w4931 and not w4932;
w4934 <= not w4790 and not w4792;
w4935 <= not w4781 and w4793;
w4936 <= not w4934 and not w4935;
w4937 <= not w329 and not w997;
w4938 <= w2481 and w4937;
w4939 <= w4292 and w4938;
w4940 <= w3373 and w4939;
w4941 <= w3821 and w4940;
w4942 <= w356 and w4941;
w4943 <= w1172 and w4942;
w4944 <= not w240 and w4943;
w4945 <= not w237 and w4944;
w4946 <= not w524 and w4945;
w4947 <= not w403 and w4946;
w4948 <= not w818 and w4947;
w4949 <= not w299 and w1644;
w4950 <= not w56 and w4949;
w4951 <= not w357 and w4950;
w4952 <= not w65 and w4951;
w4953 <= not w260 and w4952;
w4954 <= not w93 and w4953;
w4955 <= not w105 and not w760;
w4956 <= not w454 and w4955;
w4957 <= w1266 and w1796;
w4958 <= w4956 and w4957;
w4959 <= w746 and w4958;
w4960 <= w4954 and w4959;
w4961 <= w3098 and w4960;
w4962 <= not w89 and w4961;
w4963 <= not w70 and w4962;
w4964 <= not w1037 and w4963;
w4965 <= not w337 and w4964;
w4966 <= not w225 and w4965;
w4967 <= not w309 and w4966;
w4968 <= not w624 and w4967;
w4969 <= not w166 and w4968;
w4970 <= not w239 and not w448;
w4971 <= not w186 and w4970;
w4972 <= not w274 and not w333;
w4973 <= not w218 and w4972;
w4974 <= w914 and w2341;
w4975 <= not w1007 and w4974;
w4976 <= w747 and w4975;
w4977 <= w4973 and w4976;
w4978 <= w4971 and w4977;
w4979 <= w4151 and w4978;
w4980 <= w4267 and w4979;
w4981 <= w1545 and w4980;
w4982 <= w2914 and w4981;
w4983 <= w4969 and w4982;
w4984 <= w4948 and w4983;
w4985 <= not w687 and w4984;
w4986 <= not w1036 and w4985;
w4987 <= not w136 and w4986;
w4988 <= not w497 and w4987;
w4989 <= not w446 and not w681;
w4990 <= not w218 and w4989;
w4991 <= not w497 and w4990;
w4992 <= w2543 and w2978;
w4993 <= w4991 and w4992;
w4994 <= w556 and w4993;
w4995 <= w831 and w4994;
w4996 <= not w338 and w4995;
w4997 <= not w351 and w4996;
w4998 <= not w79 and w4997;
w4999 <= not w160 and not w651;
w5000 <= not w215 and not w782;
w5001 <= not w337 and w5000;
w5002 <= w4999 and w5001;
w5003 <= w1184 and w5002;
w5004 <= w4998 and w5003;
w5005 <= w599 and w5004;
w5006 <= w1603 and w5005;
w5007 <= w1602 and w5006;
w5008 <= w291 and w5007;
w5009 <= w975 and w5008;
w5010 <= not w552 and w5009;
w5011 <= not w104 and w5010;
w5012 <= not w264 and w5011;
w5013 <= not w270 and w5012;
w5014 <= not w738 and w5013;
w5015 <= not w1138 and w5014;
w5016 <= not w310 and w5015;
w5017 <= not w93 and w5016;
w5018 <= not w233 and not w760;
w5019 <= not w65 and w5018;
w5020 <= not w428 and w5019;
w5021 <= w947 and w1042;
w5022 <= w3598 and w5021;
w5023 <= w724 and w5022;
w5024 <= w746 and w5023;
w5025 <= w3029 and w5024;
w5026 <= w5020 and w5025;
w5027 <= w2105 and w5026;
w5028 <= w5017 and w5027;
w5029 <= w4948 and w5028;
w5030 <= w443 and w5029;
w5031 <= w51 and w5030;
w5032 <= w353 and w5031;
w5033 <= not w213 and w5032;
w5034 <= not w441 and w5033;
w5035 <= not w529 and w5034;
w5036 <= not w221 and w5035;
w5037 <= not w359 and w5036;
w5038 <= not w867 and w5037;
w5039 <= not w275 and w5038;
w5040 <= not w272 and w5039;
w5041 <= not w364 and w5040;
w5042 <= not w4988 and not w5041;
w5043 <= w4988 and w5041;
w5044 <= not w5042 and not w5043;
w5045 <= not a(11) and w5044;
w5046 <= not w5042 and not w5045;
w5047 <= w4286 and not w5046;
w5048 <= w2827 and not w2829;
w5049 <= not w2830 and not w5048;
w5050 <= w10 and w5049;
w5051 <= not w1299 and w2955;
w5052 <= not w1507 and w2958;
w5053 <= not w1407 and w2963;
w5054 <= not w5052 and not w5053;
w5055 <= not w5051 and w5054;
w5056 <= not w5050 and w5055;
w5057 <= not w4286 and w5046;
w5058 <= not w5047 and not w5057;
w5059 <= not w5056 and w5058;
w5060 <= not w5047 and not w5059;
w5061 <= not w4936 and not w5060;
w5062 <= w4936 and w5060;
w5063 <= not w5061 and not w5062;
w5064 <= not w5056 and not w5059;
w5065 <= w5058 and not w5059;
w5066 <= not w5064 and not w5065;
w5067 <= not a(11) and not w5045;
w5068 <= not w5043 and w5046;
w5069 <= not w5067 and not w5068;
w5070 <= not w1407 and w2955;
w5071 <= not w1507 and w2963;
w5072 <= not w1600 and w2958;
w5073 <= w2823 and not w2825;
w5074 <= not w2826 and not w5073;
w5075 <= w10 and w5074;
w5076 <= not w5072 and not w5075;
w5077 <= not w5071 and w5076;
w5078 <= not w5070 and w5077;
w5079 <= not w5069 and not w5078;
w5080 <= not w50 and w1118;
w5081 <= not w42 and w5080;
w5082 <= not w140 and w5081;
w5083 <= not w499 and w5082;
w5084 <= not w363 and w1458;
w5085 <= not w205 and w5084;
w5086 <= not w103 and w1265;
w5087 <= not w187 and w5086;
w5088 <= w5085 and w5087;
w5089 <= w856 and w5088;
w5090 <= w5083 and w5089;
w5091 <= w1570 and w5090;
w5092 <= w3586 and w5091;
w5093 <= w1520 and w5092;
w5094 <= w1850 and w5093;
w5095 <= w2419 and w5094;
w5096 <= w705 and w5095;
w5097 <= not w1007 and w5096;
w5098 <= not w449 and w5097;
w5099 <= not w225 and w5098;
w5100 <= not w760 and w5099;
w5101 <= not w608 and w5100;
w5102 <= not w472 and w5101;
w5103 <= not w260 and w5102;
w5104 <= w4988 and not w5103;
w5105 <= not w4988 and w5103;
w5106 <= not w648 and not w1036;
w5107 <= not w263 and w1063;
w5108 <= not w222 and w5107;
w5109 <= w2213 and w5108;
w5110 <= w832 and w5109;
w5111 <= w4291 and w5110;
w5112 <= w447 and w5111;
w5113 <= w589 and w5112;
w5114 <= w291 and w5113;
w5115 <= w3098 and w5114;
w5116 <= not w506 and w5115;
w5117 <= not w331 and w5116;
w5118 <= not w161 and w5117;
w5119 <= not w574 and w5118;
w5120 <= not w915 and w5119;
w5121 <= not w135 and w5120;
w5122 <= not w207 and w5121;
w5123 <= not w230 and w5122;
w5124 <= not w104 and not w397;
w5125 <= not w221 and w5124;
w5126 <= w2358 and w5125;
w5127 <= not w946 and w5126;
w5128 <= not w262 and w5127;
w5129 <= not w261 and w2175;
w5130 <= not w608 and w5129;
w5131 <= not w896 and w5130;
w5132 <= not w538 and w5131;
w5133 <= not w301 and w5132;
w5134 <= not w821 and w5133;
w5135 <= not w110 and not w388;
w5136 <= not w384 and w5135;
w5137 <= not w171 and w5136;
w5138 <= not w681 and w5137;
w5139 <= not w164 and w5138;
w5140 <= not w85 and w5139;
w5141 <= not w373 and w5140;
w5142 <= not w178 and w5141;
w5143 <= not w307 and w5142;
w5144 <= not w590 and w5143;
w5145 <= w2232 and w4248;
w5146 <= w528 and w5145;
w5147 <= w959 and w5146;
w5148 <= w1066 and w5147;
w5149 <= w5144 and w5148;
w5150 <= w5134 and w5149;
w5151 <= not w46 and w5150;
w5152 <= not w555 and w5151;
w5153 <= not w352 and w5152;
w5154 <= not w102 and w5153;
w5155 <= not w108 and w5154;
w5156 <= not w558 and w5155;
w5157 <= not w1039 and w5156;
w5158 <= not w409 and w5157;
w5159 <= not w504 and w5158;
w5160 <= w1020 and w2687;
w5161 <= w1090 and w5160;
w5162 <= w1302 and w5161;
w5163 <= not w265 and w5162;
w5164 <= not w233 and w5163;
w5165 <= not w65 and w5164;
w5166 <= not w647 and w5165;
w5167 <= not w467 and w5166;
w5168 <= not w16 and w5167;
w5169 <= w1667 and w2068;
w5170 <= not w167 and w5169;
w5171 <= not w190 and w5170;
w5172 <= not w234 and w5171;
w5173 <= not w462 and w5172;
w5174 <= not w93 and w5173;
w5175 <= w571 and w5001;
w5176 <= w1754 and w5175;
w5177 <= w5174 and w5176;
w5178 <= w5168 and w5177;
w5179 <= w5159 and w5178;
w5180 <= w5128 and w5179;
w5181 <= w5123 and w5180;
w5182 <= not w537 and w5181;
w5183 <= w5106 and w5182;
w5184 <= not w274 and w5183;
w5185 <= not w80 and w5184;
w5186 <= not w136 and w5185;
w5187 <= not w601 and w5186;
w5188 <= not w272 and w5187;
w5189 <= not w364 and w5188;
w5190 <= w2359 and w2975;
w5191 <= w1956 and w5190;
w5192 <= not w299 and w5191;
w5193 <= not w290 and w5192;
w5194 <= not w87 and w5193;
w5195 <= not w50 and w5194;
w5196 <= not w819 and w5195;
w5197 <= not w126 and w5196;
w5198 <= not w1039 and w5197;
w5199 <= not w384 and w5198;
w5200 <= w569 and w872;
w5201 <= not w210 and w5200;
w5202 <= not w175 and w5201;
w5203 <= not w123 and w5202;
w5204 <= not w184 and w5203;
w5205 <= w137 and not w448;
w5206 <= not w363 and w5205;
w5207 <= w3203 and w5206;
w5208 <= w528 and w5207;
w5209 <= w5204 and w5208;
w5210 <= w5199 and w5209;
w5211 <= w808 and w5210;
w5212 <= w807 and w5211;
w5213 <= w2281 and w5212;
w5214 <= w1510 and w5213;
w5215 <= w556 and w5214;
w5216 <= not w1241 and w5215;
w5217 <= not w219 and w5216;
w5218 <= not w360 and w5217;
w5219 <= not w241 and w5218;
w5220 <= not w92 and w5219;
w5221 <= not w454 and w5220;
w5222 <= w1539 and w2443;
w5223 <= w1038 and w5222;
w5224 <= w600 and w5223;
w5225 <= not w58 and w5224;
w5226 <= not w42 and w5225;
w5227 <= not w240 and w5226;
w5228 <= not w222 and w5227;
w5229 <= not w425 and w5228;
w5230 <= not w310 and w5229;
w5231 <= not w212 and w5230;
w5232 <= not w89 and w1183;
w5233 <= not w602 and w5232;
w5234 <= not w213 and w5233;
w5235 <= not w524 and w5234;
w5236 <= not w647 and w5235;
w5237 <= not w273 and w5236;
w5238 <= not w499 and w5237;
w5239 <= not w293 and w5238;
w5240 <= w2562 and w3199;
w5241 <= w3247 and w5240;
w5242 <= w5239 and w5241;
w5243 <= w1512 and w5242;
w5244 <= w182 and w5243;
w5245 <= w5231 and w5244;
w5246 <= w1189 and w5245;
w5247 <= w550 and w5246;
w5248 <= w5221 and w5247;
w5249 <= w35 and w5248;
w5250 <= not w270 and w5249;
w5251 <= not w337 and w5250;
w5252 <= not w760 and w5251;
w5253 <= not w231 and w5252;
w5254 <= not w127 and w5253;
w5255 <= not w364 and w5254;
w5256 <= not w5189 and not w5255;
w5257 <= w5189 and w5255;
w5258 <= not w5256 and not w5257;
w5259 <= not a(8) and w5258;
w5260 <= not w5256 and not w5259;
w5261 <= w4988 and not w5260;
w5262 <= w2815 and not w2817;
w5263 <= not w2818 and not w5262;
w5264 <= w10 and w5263;
w5265 <= not w1600 and w2955;
w5266 <= not w1812 and w2958;
w5267 <= not w1714 and w2963;
w5268 <= not w5266 and not w5267;
w5269 <= not w5265 and w5268;
w5270 <= not w5264 and w5269;
w5271 <= not w4988 and w5260;
w5272 <= not w5261 and not w5271;
w5273 <= not w5270 and w5272;
w5274 <= not w5261 and not w5273;
w5275 <= not w5104 and not w5274;
w5276 <= not w5105 and w5275;
w5277 <= not w5104 and not w5276;
w5278 <= w5069 and w5078;
w5279 <= not w5079 and not w5278;
w5280 <= not w5277 and w5279;
w5281 <= not w5079 and not w5280;
w5282 <= not w5066 and not w5281;
w5283 <= w5066 and w5281;
w5284 <= not w5282 and not w5283;
w5285 <= not w995 and w3392;
w5286 <= not w1170 and w3477;
w5287 <= not w1113 and w3541;
w5288 <= not w5286 and not w5287;
w5289 <= not w5285 and w5288;
w5290 <= not w3303 and w5289;
w5291 <= not w4364 and w5289;
w5292 <= not w5290 and not w5291;
w5293 <= a(29) and not w5292;
w5294 <= not a(29) and w5292;
w5295 <= not w5293 and not w5294;
w5296 <= w5284 and not w5295;
w5297 <= not w5282 and not w5296;
w5298 <= w5063 and not w5297;
w5299 <= not w5061 and not w5298;
w5300 <= not w4933 and not w5299;
w5301 <= not w4930 and not w5300;
w5302 <= not w4810 and w4821;
w5303 <= not w4822 and not w5302;
w5304 <= not w5301 and w5303;
w5305 <= w5301 and not w5303;
w5306 <= not w5304 and not w5305;
w5307 <= not w2947 and w3819;
w5308 <= not w522 and w3902;
w5309 <= not w327 and w3981;
w5310 <= not w5308 and not w5309;
w5311 <= not w5307 and w5310;
w5312 <= w2953 and w3985;
w5313 <= w5311 and not w5312;
w5314 <= a(26) and not w5313;
w5315 <= a(26) and not w5314;
w5316 <= not w5313 and not w5314;
w5317 <= not w5315 and not w5316;
w5318 <= w5306 and not w5317;
w5319 <= not w5304 and not w5318;
w5320 <= not w4915 and not w5319;
w5321 <= w4915 and w5319;
w5322 <= not w5320 and not w5321;
w5323 <= not w3740 and w4629;
w5324 <= not w3540 and w4468;
w5325 <= not w3391 and w4539;
w5326 <= not w5324 and not w5325;
w5327 <= not w5323 and w5326;
w5328 <= w3753 and w4471;
w5329 <= w5327 and not w5328;
w5330 <= a(23) and not w5329;
w5331 <= a(23) and not w5330;
w5332 <= not w5329 and not w5330;
w5333 <= not w5331 and not w5332;
w5334 <= w5322 and not w5333;
w5335 <= not w5320 and not w5334;
w5336 <= not w4912 and not w5335;
w5337 <= not w4909 and not w5336;
w5338 <= not w4895 and not w5337;
w5339 <= w4895 and w5337;
w5340 <= not w5338 and not w5339;
w5341 <= not w3812 and w4870;
w5342 <= not w4862 and w4868;
w5343 <= not w4450 and w5342;
w5344 <= not w5341 and not w5343;
w5345 <= w4544 and w4873;
w5346 <= w5344 and not w5345;
w5347 <= a(20) and not w5346;
w5348 <= a(20) and not w5347;
w5349 <= not w5346 and not w5347;
w5350 <= not w5348 and not w5349;
w5351 <= w5340 and not w5350;
w5352 <= not w5338 and not w5351;
w5353 <= not w4892 and not w5352;
w5354 <= w4892 and w5352;
w5355 <= not w5353 and not w5354;
w5356 <= w5340 and not w5351;
w5357 <= not w5350 and not w5351;
w5358 <= not w5356 and not w5357;
w5359 <= w5322 and not w5334;
w5360 <= not w5333 and not w5334;
w5361 <= not w5359 and not w5360;
w5362 <= w5306 and not w5318;
w5363 <= not w5317 and not w5318;
w5364 <= not w5362 and not w5363;
w5365 <= w4933 and w5299;
w5366 <= not w5300 and not w5365;
w5367 <= not w327 and w3819;
w5368 <= not w645 and w3902;
w5369 <= not w522 and w3981;
w5370 <= not w5368 and not w5369;
w5371 <= not w5367 and w5370;
w5372 <= not w3985 and w5371;
w5373 <= not w3282 and w5371;
w5374 <= not w5372 and not w5373;
w5375 <= a(26) and not w5374;
w5376 <= not a(26) and w5374;
w5377 <= not w5375 and not w5376;
w5378 <= w5366 and not w5377;
w5379 <= not w522 and w3819;
w5380 <= not w802 and w3902;
w5381 <= not w645 and w3981;
w5382 <= not w5380 and not w5381;
w5383 <= not w5379 and w5382;
w5384 <= w3266 and w3985;
w5385 <= w5383 and not w5384;
w5386 <= a(26) and not w5385;
w5387 <= a(26) and not w5386;
w5388 <= not w5385 and not w5386;
w5389 <= not w5387 and not w5388;
w5390 <= not w5063 and w5297;
w5391 <= not w5298 and not w5390;
w5392 <= not w893 and w3392;
w5393 <= not w1113 and w3477;
w5394 <= not w995 and w3541;
w5395 <= not w5393 and not w5394;
w5396 <= not w5392 and w5395;
w5397 <= not w3303 and w5396;
w5398 <= not w4568 and w5396;
w5399 <= not w5397 and not w5398;
w5400 <= a(29) and not w5399;
w5401 <= not a(29) and w5399;
w5402 <= not w5400 and not w5401;
w5403 <= w5391 and not w5402;
w5404 <= not w5391 and w5402;
w5405 <= not w5403 and not w5404;
w5406 <= not w5389 and w5405;
w5407 <= not w5403 and not w5406;
w5408 <= not w5366 and w5377;
w5409 <= not w5378 and not w5408;
w5410 <= not w5407 and w5409;
w5411 <= not w5378 and not w5410;
w5412 <= not w5364 and not w5411;
w5413 <= w5364 and w5411;
w5414 <= not w5412 and not w5413;
w5415 <= not w3391 and w4629;
w5416 <= not w3474 and w4468;
w5417 <= not w3540 and w4539;
w5418 <= not w5416 and not w5417;
w5419 <= not w5415 and w5418;
w5420 <= w3562 and w4471;
w5421 <= w5419 and not w5420;
w5422 <= a(23) and not w5421;
w5423 <= a(23) and not w5422;
w5424 <= not w5421 and not w5422;
w5425 <= not w5423 and not w5424;
w5426 <= w5414 and not w5425;
w5427 <= not w5412 and not w5426;
w5428 <= not w5361 and not w5427;
w5429 <= w5361 and w5427;
w5430 <= not w5428 and not w5429;
w5431 <= w4865 and not w4868;
w5432 <= not w3812 and w5431;
w5433 <= not w3899 and w4870;
w5434 <= not w3980 and w5342;
w5435 <= not w5433 and not w5434;
w5436 <= not w5432 and w5435;
w5437 <= w4002 and w4873;
w5438 <= w5436 and not w5437;
w5439 <= a(20) and not w5438;
w5440 <= a(20) and not w5439;
w5441 <= not w5438 and not w5439;
w5442 <= not w5440 and not w5441;
w5443 <= w5430 and not w5442;
w5444 <= not w5428 and not w5443;
w5445 <= not w4450 and w5431;
w5446 <= not w3980 and w4870;
w5447 <= not w3812 and w5342;
w5448 <= not w5446 and not w5447;
w5449 <= not w5445 and w5448;
w5450 <= not w4873 and w5449;
w5451 <= not w4650 and w5449;
w5452 <= not w5450 and not w5451;
w5453 <= a(20) and not w5452;
w5454 <= not a(20) and w5452;
w5455 <= not w5453 and not w5454;
w5456 <= not w5444 and not w5455;
w5457 <= w4912 and w5335;
w5458 <= not w5336 and not w5457;
w5459 <= w5444 and w5455;
w5460 <= not w5456 and not w5459;
w5461 <= w5458 and w5460;
w5462 <= not w5456 and not w5461;
w5463 <= not w5358 and not w5462;
w5464 <= w5358 and w5462;
w5465 <= not w5463 and not w5464;
w5466 <= w5414 and not w5426;
w5467 <= not w5425 and not w5426;
w5468 <= not w5466 and not w5467;
w5469 <= not w3540 and w4629;
w5470 <= not w2947 and w4468;
w5471 <= not w3474 and w4539;
w5472 <= not w5470 and not w5471;
w5473 <= not w5469 and w5472;
w5474 <= w4019 and w4471;
w5475 <= w5473 and not w5474;
w5476 <= a(23) and not w5475;
w5477 <= not w5475 and not w5476;
w5478 <= a(23) and not w5476;
w5479 <= not w5477 and not w5478;
w5480 <= w5407 and not w5409;
w5481 <= not w5410 and not w5480;
w5482 <= not w5479 and w5481;
w5483 <= not w5479 and not w5482;
w5484 <= w5481 and not w5482;
w5485 <= not w5483 and not w5484;
w5486 <= w5405 and not w5406;
w5487 <= not w5389 and not w5406;
w5488 <= not w5486 and not w5487;
w5489 <= not w5274 and not w5276;
w5490 <= not w5105 and w5277;
w5491 <= not w5489 and not w5490;
w5492 <= not w1507 and w2955;
w5493 <= not w1600 and w2963;
w5494 <= not w1714 and w2958;
w5495 <= w2819 and not w2821;
w5496 <= not w2822 and not w5495;
w5497 <= w10 and w5496;
w5498 <= not w5494 and not w5497;
w5499 <= not w5493 and w5498;
w5500 <= not w5492 and w5499;
w5501 <= not w5491 and not w5500;
w5502 <= not w1170 and w3392;
w5503 <= not w1407 and w3477;
w5504 <= not w1299 and w3541;
w5505 <= not w5503 and not w5504;
w5506 <= not w5502 and w5505;
w5507 <= w3303 and w4783;
w5508 <= w5506 and not w5507;
w5509 <= a(29) and not w5508;
w5510 <= not w5508 and not w5509;
w5511 <= a(29) and not w5509;
w5512 <= not w5510 and not w5511;
w5513 <= not w5491 and not w5501;
w5514 <= not w5500 and not w5501;
w5515 <= not w5513 and not w5514;
w5516 <= not w5512 and not w5515;
w5517 <= not w5501 and not w5516;
w5518 <= w5277 and not w5279;
w5519 <= not w5280 and not w5518;
w5520 <= not w5517 and w5519;
w5521 <= not w1113 and w3392;
w5522 <= not w1299 and w3477;
w5523 <= not w1170 and w3541;
w5524 <= not w5522 and not w5523;
w5525 <= not w5521 and w5524;
w5526 <= w3303 and w4796;
w5527 <= w5525 and not w5526;
w5528 <= a(29) and not w5527;
w5529 <= a(29) and not w5528;
w5530 <= not w5527 and not w5528;
w5531 <= not w5529 and not w5530;
w5532 <= w5517 and not w5519;
w5533 <= not w5520 and not w5532;
w5534 <= not w5531 and w5533;
w5535 <= not w5520 and not w5534;
w5536 <= not w5284 and w5295;
w5537 <= not w5296 and not w5536;
w5538 <= not w5535 and w5537;
w5539 <= w5535 and not w5537;
w5540 <= not w5538 and not w5539;
w5541 <= not w645 and w3819;
w5542 <= not w893 and w3902;
w5543 <= not w802 and w3981;
w5544 <= not w5542 and not w5543;
w5545 <= not w5541 and w5544;
w5546 <= w3985 and w4114;
w5547 <= w5545 and not w5546;
w5548 <= a(26) and not w5547;
w5549 <= a(26) and not w5548;
w5550 <= not w5547 and not w5548;
w5551 <= not w5549 and not w5550;
w5552 <= w5540 and not w5551;
w5553 <= not w5538 and not w5552;
w5554 <= not w5488 and not w5553;
w5555 <= w5488 and w5553;
w5556 <= not w5554 and not w5555;
w5557 <= not w3474 and w4629;
w5558 <= not w327 and w4468;
w5559 <= not w2947 and w4539;
w5560 <= not w5558 and not w5559;
w5561 <= not w5557 and w5560;
w5562 <= w3650 and w4471;
w5563 <= w5561 and not w5562;
w5564 <= a(23) and not w5563;
w5565 <= a(23) and not w5564;
w5566 <= not w5563 and not w5564;
w5567 <= not w5565 and not w5566;
w5568 <= w5556 and not w5567;
w5569 <= not w5554 and not w5568;
w5570 <= not w5485 and not w5569;
w5571 <= not w5482 and not w5570;
w5572 <= not w5468 and not w5571;
w5573 <= w5468 and w5571;
w5574 <= not w5572 and not w5573;
w5575 <= not w3980 and w5431;
w5576 <= not w3740 and w4870;
w5577 <= not w3899 and w5342;
w5578 <= not w5576 and not w5577;
w5579 <= not w5575 and w5578;
w5580 <= w4412 and w4873;
w5581 <= w5579 and not w5580;
w5582 <= a(20) and not w5581;
w5583 <= a(20) and not w5582;
w5584 <= not w5581 and not w5582;
w5585 <= not w5583 and not w5584;
w5586 <= w5574 and not w5585;
w5587 <= not w5572 and not w5586;
w5588 <= not a(15) and a(16);
w5589 <= a(15) and not a(16);
w5590 <= not w5588 and not w5589;
w5591 <= a(14) and not a(15);
w5592 <= not a(14) and a(15);
w5593 <= not w5591 and not w5592;
w5594 <= a(16) and not a(17);
w5595 <= not a(16) and a(17);
w5596 <= not w5594 and not w5595;
w5597 <= w5593 and not w5596;
w5598 <= w5590 and w5597;
w5599 <= not w4450 and w5598;
w5600 <= not w4457 and not w5599;
w5601 <= not w5593 and not w5596;
w5602 <= not w5599 and not w5601;
w5603 <= not w5600 and not w5602;
w5604 <= a(17) and not w5603;
w5605 <= not a(17) and w5603;
w5606 <= not w5604 and not w5605;
w5607 <= not w5587 and not w5606;
w5608 <= w5430 and not w5443;
w5609 <= not w5442 and not w5443;
w5610 <= not w5608 and not w5609;
w5611 <= w5587 and w5606;
w5612 <= not w5607 and not w5611;
w5613 <= not w5610 and w5612;
w5614 <= not w5607 and not w5613;
w5615 <= not w5458 and not w5460;
w5616 <= not w5461 and not w5615;
w5617 <= not w5614 and w5616;
w5618 <= not w5610 and not w5613;
w5619 <= w5612 and not w5613;
w5620 <= not w5618 and not w5619;
w5621 <= w5574 and not w5586;
w5622 <= not w5585 and not w5586;
w5623 <= not w5621 and not w5622;
w5624 <= w5485 and w5569;
w5625 <= not w5570 and not w5624;
w5626 <= not w3899 and w5431;
w5627 <= not w3391 and w4870;
w5628 <= not w3740 and w5342;
w5629 <= not w5627 and not w5628;
w5630 <= not w5626 and w5629;
w5631 <= not w4873 and w5630;
w5632 <= not w4493 and w5630;
w5633 <= not w5631 and not w5632;
w5634 <= a(20) and not w5633;
w5635 <= not a(20) and w5633;
w5636 <= not w5634 and not w5635;
w5637 <= w5625 and not w5636;
w5638 <= w5556 and not w5568;
w5639 <= not w5567 and not w5568;
w5640 <= not w5638 and not w5639;
w5641 <= w5540 and not w5552;
w5642 <= not w5551 and not w5552;
w5643 <= not w5641 and not w5642;
w5644 <= w5533 and not w5534;
w5645 <= not w5531 and not w5534;
w5646 <= not w5644 and not w5645;
w5647 <= not w802 and w3819;
w5648 <= not w995 and w3902;
w5649 <= not w893 and w3981;
w5650 <= not w5648 and not w5649;
w5651 <= not w5647 and w5650;
w5652 <= not w3985 and w5651;
w5653 <= not w4139 and w5651;
w5654 <= not w5652 and not w5653;
w5655 <= a(26) and not w5654;
w5656 <= not a(26) and w5654;
w5657 <= not w5655 and not w5656;
w5658 <= not w5646 and not w5657;
w5659 <= not w5512 and not w5516;
w5660 <= not w5515 and not w5516;
w5661 <= not w5659 and not w5660;
w5662 <= not w5270 and not w5273;
w5663 <= w5272 and not w5273;
w5664 <= not w5662 and not w5663;
w5665 <= not a(8) and not w5259;
w5666 <= not w5257 and w5260;
w5667 <= not w5665 and not w5666;
w5668 <= w468 and w526;
w5669 <= not w231 and w5668;
w5670 <= w3622 and w5669;
w5671 <= w3518 and w5670;
w5672 <= w1359 and w5671;
w5673 <= w3095 and w5672;
w5674 <= w912 and w5673;
w5675 <= w1510 and w5674;
w5676 <= not w404 and w5675;
w5677 <= not w819 and w5676;
w5678 <= not w472 and w5677;
w5679 <= not w1138 and w5678;
w5680 <= not w384 and w5679;
w5681 <= not w590 and w5680;
w5682 <= not w224 and not w299;
w5683 <= not w222 and w5682;
w5684 <= w593 and w5683;
w5685 <= w5204 and w5684;
w5686 <= w759 and w5685;
w5687 <= w5174 and w5686;
w5688 <= w3140 and w5687;
w5689 <= w5681 and w5688;
w5690 <= w2568 and w5689;
w5691 <= w43 and w5690;
w5692 <= w505 and w5691;
w5693 <= not w289 and w5692;
w5694 <= not w50 and w5693;
w5695 <= not w112 and w5694;
w5696 <= not w292 and w5695;
w5697 <= not w498 and w5696;
w5698 <= not w108 and w5697;
w5699 <= not w536 and w5698;
w5700 <= not w218 and w5699;
w5701 <= w5189 and not w5700;
w5702 <= not w5189 and w5700;
w5703 <= w1432 and w3459;
w5704 <= not w171 and w5703;
w5705 <= not w439 and w5704;
w5706 <= not w140 and w5705;
w5707 <= not w472 and w5706;
w5708 <= not w601 and w5707;
w5709 <= not w299 and not w365;
w5710 <= not w62 and w5709;
w5711 <= not w216 and not w263;
w5712 <= not w138 and w5711;
w5713 <= w5710 and w5712;
w5714 <= not w177 and w5713;
w5715 <= not w103 and w5714;
w5716 <= not w819 and w5715;
w5717 <= not w222 and w5716;
w5718 <= not w896 and w5717;
w5719 <= not w21 and w5718;
w5720 <= not w93 and w5719;
w5721 <= not w386 and not w867;
w5722 <= not w298 and w5721;
w5723 <= not w71 and w5722;
w5724 <= not w446 and w5723;
w5725 <= not w210 and w5724;
w5726 <= not w163 and w5725;
w5727 <= not w86 and not w537;
w5728 <= not w124 and w5727;
w5729 <= w5726 and w5728;
w5730 <= w5720 and w5729;
w5731 <= w1172 and w5730;
w5732 <= w162 and w5731;
w5733 <= w35 and w5732;
w5734 <= w2693 and w5733;
w5735 <= not w555 and w5734;
w5736 <= not w441 and w5735;
w5737 <= not w56 and w5736;
w5738 <= not w462 and w5737;
w5739 <= not w79 and w5738;
w5740 <= not w428 and w5739;
w5741 <= not w1062 and w5740;
w5742 <= not w265 and not w384;
w5743 <= not w157 and w5742;
w5744 <= w2925 and w5743;
w5745 <= w5741 and w5744;
w5746 <= w4323 and w5745;
w5747 <= w551 and w5746;
w5748 <= w5708 and w5747;
w5749 <= w2586 and w5748;
w5750 <= w2875 and w5749;
w5751 <= w455 and w5750;
w5752 <= not w782 and w5751;
w5753 <= not w648 and w5752;
w5754 <= not w106 and w5753;
w5755 <= not w395 and w5754;
w5756 <= not w266 and w5755;
w5757 <= not w181 and w5756;
w5758 <= not w558 and w5757;
w5759 <= not w16 and w5758;
w5760 <= not w166 and w5759;
w5761 <= not a(2) and not w5760;
w5762 <= a(2) and not w5760;
w5763 <= not a(2) and w5760;
w5764 <= not w5762 and not w5763;
w5765 <= not a(5) and not w5764;
w5766 <= not w5761 and not w5765;
w5767 <= w5189 and not w5766;
w5768 <= w2803 and not w2805;
w5769 <= not w2806 and not w5768;
w5770 <= w10 and w5769;
w5771 <= not w1848 and w2955;
w5772 <= not w1992 and w2958;
w5773 <= not w1927 and w2963;
w5774 <= not w5772 and not w5773;
w5775 <= not w5771 and w5774;
w5776 <= not w5770 and w5775;
w5777 <= not w5189 and w5766;
w5778 <= not w5767 and not w5777;
w5779 <= not w5776 and w5778;
w5780 <= not w5767 and not w5779;
w5781 <= not w5701 and not w5780;
w5782 <= not w5702 and w5781;
w5783 <= not w5701 and not w5782;
w5784 <= not w5667 and not w5783;
w5785 <= w2811 and not w2813;
w5786 <= not w2814 and not w5785;
w5787 <= w10 and w5786;
w5788 <= not w1714 and w2955;
w5789 <= not w1848 and w2958;
w5790 <= not w1812 and w2963;
w5791 <= not w5789 and not w5790;
w5792 <= not w5788 and w5791;
w5793 <= not w5787 and w5792;
w5794 <= w5667 and w5783;
w5795 <= not w5784 and not w5794;
w5796 <= not w5793 and w5795;
w5797 <= not w5784 and not w5796;
w5798 <= not w5664 and not w5797;
w5799 <= w5664 and w5797;
w5800 <= not w5798 and not w5799;
w5801 <= not w1299 and w3392;
w5802 <= not w1507 and w3477;
w5803 <= not w1407 and w3541;
w5804 <= not w5802 and not w5803;
w5805 <= not w5801 and w5804;
w5806 <= not w3303 and w5805;
w5807 <= not w5049 and w5805;
w5808 <= not w5806 and not w5807;
w5809 <= a(29) and not w5808;
w5810 <= not a(29) and w5808;
w5811 <= not w5809 and not w5810;
w5812 <= w5800 and not w5811;
w5813 <= not w5798 and not w5812;
w5814 <= not w5661 and not w5813;
w5815 <= w5661 and w5813;
w5816 <= not w5814 and not w5815;
w5817 <= not w893 and w3819;
w5818 <= not w1113 and w3902;
w5819 <= not w995 and w3981;
w5820 <= not w5818 and not w5819;
w5821 <= not w5817 and w5820;
w5822 <= w3985 and w4568;
w5823 <= w5821 and not w5822;
w5824 <= a(26) and not w5823;
w5825 <= a(26) and not w5824;
w5826 <= not w5823 and not w5824;
w5827 <= not w5825 and not w5826;
w5828 <= w5816 and not w5827;
w5829 <= not w5814 and not w5828;
w5830 <= w5646 and w5657;
w5831 <= not w5658 and not w5830;
w5832 <= not w5829 and w5831;
w5833 <= not w5658 and not w5832;
w5834 <= not w5643 and not w5833;
w5835 <= w5643 and w5833;
w5836 <= not w5834 and not w5835;
w5837 <= not w2947 and w4629;
w5838 <= not w522 and w4468;
w5839 <= not w327 and w4539;
w5840 <= not w5838 and not w5839;
w5841 <= not w5837 and w5840;
w5842 <= w2953 and w4471;
w5843 <= w5841 and not w5842;
w5844 <= a(23) and not w5843;
w5845 <= a(23) and not w5844;
w5846 <= not w5843 and not w5844;
w5847 <= not w5845 and not w5846;
w5848 <= w5836 and not w5847;
w5849 <= not w5834 and not w5848;
w5850 <= not w5640 and not w5849;
w5851 <= w5640 and w5849;
w5852 <= not w5850 and not w5851;
w5853 <= not w3740 and w5431;
w5854 <= not w3540 and w4870;
w5855 <= not w3391 and w5342;
w5856 <= not w5854 and not w5855;
w5857 <= not w5853 and w5856;
w5858 <= w3753 and w4873;
w5859 <= w5857 and not w5858;
w5860 <= a(20) and not w5859;
w5861 <= a(20) and not w5860;
w5862 <= not w5859 and not w5860;
w5863 <= not w5861 and not w5862;
w5864 <= w5852 and not w5863;
w5865 <= not w5850 and not w5864;
w5866 <= not w5625 and w5636;
w5867 <= not w5637 and not w5866;
w5868 <= not w5865 and w5867;
w5869 <= not w5637 and not w5868;
w5870 <= not w5623 and not w5869;
w5871 <= w5623 and w5869;
w5872 <= not w5870 and not w5871;
w5873 <= not w3812 and w5598;
w5874 <= not w5590 and w5593;
w5875 <= not w4450 and w5874;
w5876 <= not w5873 and not w5875;
w5877 <= w4544 and w5601;
w5878 <= w5876 and not w5877;
w5879 <= a(17) and not w5878;
w5880 <= a(17) and not w5879;
w5881 <= not w5878 and not w5879;
w5882 <= not w5880 and not w5881;
w5883 <= w5872 and not w5882;
w5884 <= not w5870 and not w5883;
w5885 <= not w5620 and not w5884;
w5886 <= w5620 and w5884;
w5887 <= not w5885 and not w5886;
w5888 <= w5872 and not w5883;
w5889 <= not w5882 and not w5883;
w5890 <= not w5888 and not w5889;
w5891 <= w5852 and not w5864;
w5892 <= not w5863 and not w5864;
w5893 <= not w5891 and not w5892;
w5894 <= w5836 and not w5848;
w5895 <= not w5847 and not w5848;
w5896 <= not w5894 and not w5895;
w5897 <= not w327 and w4629;
w5898 <= not w645 and w4468;
w5899 <= not w522 and w4539;
w5900 <= not w5898 and not w5899;
w5901 <= not w5897 and w5900;
w5902 <= w3282 and w4471;
w5903 <= w5901 and not w5902;
w5904 <= a(23) and not w5903;
w5905 <= not w5903 and not w5904;
w5906 <= a(23) and not w5904;
w5907 <= not w5905 and not w5906;
w5908 <= w5829 and not w5831;
w5909 <= not w5832 and not w5908;
w5910 <= not w5907 and w5909;
w5911 <= not w5907 and not w5910;
w5912 <= w5909 and not w5910;
w5913 <= not w5911 and not w5912;
w5914 <= w5816 and not w5828;
w5915 <= not w5827 and not w5828;
w5916 <= not w5914 and not w5915;
w5917 <= not w1407 and w3392;
w5918 <= not w1600 and w3477;
w5919 <= not w1507 and w3541;
w5920 <= not w5918 and not w5919;
w5921 <= not w5917 and w5920;
w5922 <= w3303 and w5074;
w5923 <= w5921 and not w5922;
w5924 <= a(29) and not w5923;
w5925 <= not w5923 and not w5924;
w5926 <= a(29) and not w5924;
w5927 <= not w5925 and not w5926;
w5928 <= not w5793 and not w5796;
w5929 <= w5795 and not w5796;
w5930 <= not w5928 and not w5929;
w5931 <= not w5927 and not w5930;
w5932 <= not w5927 and not w5931;
w5933 <= not w5930 and not w5931;
w5934 <= not w5932 and not w5933;
w5935 <= not w5780 and not w5782;
w5936 <= not w5702 and w5783;
w5937 <= not w5935 and not w5936;
w5938 <= not w1812 and w2955;
w5939 <= not w1848 and w2963;
w5940 <= not w1927 and w2958;
w5941 <= w2807 and not w2809;
w5942 <= not w2810 and not w5941;
w5943 <= w10 and w5942;
w5944 <= not w5940 and not w5943;
w5945 <= not w5939 and w5944;
w5946 <= not w5938 and w5945;
w5947 <= not w5937 and not w5946;
w5948 <= not w5776 and not w5779;
w5949 <= w5778 and not w5779;
w5950 <= not w5948 and not w5949;
w5951 <= not w224 and w1994;
w5952 <= not w555 and w5951;
w5953 <= not w287 and w5952;
w5954 <= not w329 and w5953;
w5955 <= not w538 and w5954;
w5956 <= w1662 and w2640;
w5957 <= w2491 and w5956;
w5958 <= not w265 and w5957;
w5959 <= not w401 and w5958;
w5960 <= w1615 and w5959;
w5961 <= not w205 and w5960;
w5962 <= w4270 and w5087;
w5963 <= w4991 and w5962;
w5964 <= w1019 and w5963;
w5965 <= w2062 and w5964;
w5966 <= w3515 and w5965;
w5967 <= w5961 and w5966;
w5968 <= w2374 and w5967;
w5969 <= w5955 and w5968;
w5970 <= w964 and w5969;
w5971 <= w4721 and w5970;
w5972 <= w553 and w5971;
w5973 <= not w178 and w5972;
w5974 <= not w454 and w5973;
w5975 <= not w62 and w5974;
w5976 <= not w16 and w5975;
w5977 <= a(2) and not w5976;
w5978 <= not a(2) and w5976;
w5979 <= w402 and w1546;
w5980 <= not w355 and w5979;
w5981 <= not w997 and w5980;
w5982 <= not w352 and w5981;
w5983 <= not w335 and w5982;
w5984 <= not w351 and w5983;
w5985 <= not w127 and w5984;
w5986 <= not w498 and w5985;
w5987 <= not w360 and w5986;
w5988 <= not w649 and w5987;
w5989 <= not w178 and w5988;
w5990 <= w625 and w3187;
w5991 <= w553 and w5990;
w5992 <= w4763 and w5991;
w5993 <= w139 and w5992;
w5994 <= w259 and w5993;
w5995 <= w5989 and w5994;
w5996 <= w2558 and w5995;
w5997 <= w2896 and w5996;
w5998 <= w4209 and w5997;
w5999 <= w539 and w5998;
w6000 <= w389 and w5999;
w6001 <= w358 and w6000;
w6002 <= w666 and w6001;
w6003 <= w1314 and w6002;
w6004 <= not w84 and w6003;
w6005 <= not w181 and w6004;
w6006 <= not w726 and w6005;
w6007 <= not w527 and w6006;
w6008 <= not w821 and w6007;
w6009 <= not w384 and w6008;
w6010 <= a(2) and not w6009;
w6011 <= not a(2) and w6009;
w6012 <= w1361 and w1579;
w6013 <= not w125 and w6012;
w6014 <= not w174 and w6013;
w6015 <= not w572 and w6014;
w6016 <= not w240 and w6015;
w6017 <= not w65 and w6016;
w6018 <= not w945 and w6017;
w6019 <= not w230 and not w330;
w6020 <= w2528 and w5085;
w6021 <= w1373 and w6020;
w6022 <= w6019 and w6021;
w6023 <= w5128 and w6022;
w6024 <= w1536 and w6023;
w6025 <= w964 and w6024;
w6026 <= w389 and w6025;
w6027 <= w914 and w6026;
w6028 <= not w687 and w6027;
w6029 <= not w159 and w6028;
w6030 <= not w210 and w6029;
w6031 <= not w161 and w6030;
w6032 <= not w386 and w6031;
w6033 <= w525 and not w1007;
w6034 <= not w141 and w6033;
w6035 <= not w649 and w6034;
w6036 <= not w624 and w6035;
w6037 <= not w409 and w6036;
w6038 <= not w46 and w4302;
w6039 <= not w538 and w6038;
w6040 <= w4204 and w6039;
w6041 <= w2176 and w6040;
w6042 <= w2742 and w6041;
w6043 <= w6037 and w6042;
w6044 <= w2686 and w6043;
w6045 <= w6032 and w6044;
w6046 <= w6018 and w6045;
w6047 <= w268 and w6046;
w6048 <= w1226 and w6047;
w6049 <= w4721 and w6048;
w6050 <= not w136 and w6049;
w6051 <= not w499 and w6050;
w6052 <= not w424 and w6051;
w6053 <= not w821 and w6052;
w6054 <= a(2) and not w6053;
w6055 <= not a(2) and w6053;
w6056 <= w2787 and not w2789;
w6057 <= not w2790 and not w6056;
w6058 <= w10 and w6057;
w6059 <= not w2124 and w2955;
w6060 <= not w2323 and w2958;
w6061 <= not w2226 and w2963;
w6062 <= not w6060 and not w6061;
w6063 <= not w6059 and w6062;
w6064 <= not w6058 and w6063;
w6065 <= not w6054 and not w6064;
w6066 <= not w6055 and w6065;
w6067 <= not w6054 and not w6066;
w6068 <= not w6010 and not w6067;
w6069 <= not w6011 and w6068;
w6070 <= not w6010 and not w6069;
w6071 <= not w5977 and not w6070;
w6072 <= not w5978 and w6071;
w6073 <= not w5977 and not w6072;
w6074 <= a(5) and w5764;
w6075 <= not w5765 and not w6074;
w6076 <= not w6073 and w6075;
w6077 <= w2799 and not w2801;
w6078 <= not w2802 and not w6077;
w6079 <= w10 and w6078;
w6080 <= not w1927 and w2955;
w6081 <= not w2087 and w2958;
w6082 <= not w1992 and w2963;
w6083 <= not w6081 and not w6082;
w6084 <= not w6080 and w6083;
w6085 <= not w6079 and w6084;
w6086 <= w6073 and not w6075;
w6087 <= not w6076 and not w6086;
w6088 <= not w6085 and w6087;
w6089 <= not w6076 and not w6088;
w6090 <= not w5950 and not w6089;
w6091 <= w5950 and w6089;
w6092 <= not w6090 and not w6091;
w6093 <= not w1600 and w3392;
w6094 <= not w1812 and w3477;
w6095 <= not w1714 and w3541;
w6096 <= not w6094 and not w6095;
w6097 <= not w6093 and w6096;
w6098 <= not w3303 and w6097;
w6099 <= not w5263 and w6097;
w6100 <= not w6098 and not w6099;
w6101 <= a(29) and not w6100;
w6102 <= not a(29) and w6100;
w6103 <= not w6101 and not w6102;
w6104 <= w6092 and not w6103;
w6105 <= not w6090 and not w6104;
w6106 <= not w5937 and not w5947;
w6107 <= not w5946 and not w5947;
w6108 <= not w6106 and not w6107;
w6109 <= not w6105 and not w6108;
w6110 <= not w5947 and not w6109;
w6111 <= not w5934 and not w6110;
w6112 <= not w5931 and not w6111;
w6113 <= not w5800 and w5811;
w6114 <= not w5812 and not w6113;
w6115 <= not w6112 and w6114;
w6116 <= w6112 and not w6114;
w6117 <= not w6115 and not w6116;
w6118 <= not w995 and w3819;
w6119 <= not w1170 and w3902;
w6120 <= not w1113 and w3981;
w6121 <= not w6119 and not w6120;
w6122 <= not w6118 and w6121;
w6123 <= w3985 and w4364;
w6124 <= w6122 and not w6123;
w6125 <= a(26) and not w6124;
w6126 <= a(26) and not w6125;
w6127 <= not w6124 and not w6125;
w6128 <= not w6126 and not w6127;
w6129 <= w6117 and not w6128;
w6130 <= not w6115 and not w6129;
w6131 <= not w5916 and not w6130;
w6132 <= w5916 and w6130;
w6133 <= not w6131 and not w6132;
w6134 <= not w522 and w4629;
w6135 <= not w802 and w4468;
w6136 <= not w645 and w4539;
w6137 <= not w6135 and not w6136;
w6138 <= not w6134 and w6137;
w6139 <= w3266 and w4471;
w6140 <= w6138 and not w6139;
w6141 <= a(23) and not w6140;
w6142 <= a(23) and not w6141;
w6143 <= not w6140 and not w6141;
w6144 <= not w6142 and not w6143;
w6145 <= w6133 and not w6144;
w6146 <= not w6131 and not w6145;
w6147 <= not w5913 and not w6146;
w6148 <= not w5910 and not w6147;
w6149 <= not w5896 and not w6148;
w6150 <= w5896 and w6148;
w6151 <= not w6149 and not w6150;
w6152 <= not w3391 and w5431;
w6153 <= not w3474 and w4870;
w6154 <= not w3540 and w5342;
w6155 <= not w6153 and not w6154;
w6156 <= not w6152 and w6155;
w6157 <= w3562 and w4873;
w6158 <= w6156 and not w6157;
w6159 <= a(20) and not w6158;
w6160 <= a(20) and not w6159;
w6161 <= not w6158 and not w6159;
w6162 <= not w6160 and not w6161;
w6163 <= w6151 and not w6162;
w6164 <= not w6149 and not w6163;
w6165 <= not w5893 and not w6164;
w6166 <= w5893 and w6164;
w6167 <= not w6165 and not w6166;
w6168 <= not w5593 and w5596;
w6169 <= not w3812 and w6168;
w6170 <= not w3899 and w5598;
w6171 <= not w3980 and w5874;
w6172 <= not w6170 and not w6171;
w6173 <= not w6169 and w6172;
w6174 <= w4002 and w5601;
w6175 <= w6173 and not w6174;
w6176 <= a(17) and not w6175;
w6177 <= a(17) and not w6176;
w6178 <= not w6175 and not w6176;
w6179 <= not w6177 and not w6178;
w6180 <= w6167 and not w6179;
w6181 <= not w6165 and not w6180;
w6182 <= not w4450 and w6168;
w6183 <= not w3980 and w5598;
w6184 <= not w3812 and w5874;
w6185 <= not w6183 and not w6184;
w6186 <= not w6182 and w6185;
w6187 <= not w5601 and w6186;
w6188 <= not w4650 and w6186;
w6189 <= not w6187 and not w6188;
w6190 <= a(17) and not w6189;
w6191 <= not a(17) and w6189;
w6192 <= not w6190 and not w6191;
w6193 <= not w6181 and not w6192;
w6194 <= w6181 and w6192;
w6195 <= not w6193 and not w6194;
w6196 <= w5865 and not w5867;
w6197 <= not w5868 and not w6196;
w6198 <= w6195 and w6197;
w6199 <= not w6193 and not w6198;
w6200 <= not w5890 and not w6199;
w6201 <= w5890 and w6199;
w6202 <= not w6200 and not w6201;
w6203 <= w6151 and not w6163;
w6204 <= not w6162 and not w6163;
w6205 <= not w6203 and not w6204;
w6206 <= w5913 and w6146;
w6207 <= not w6147 and not w6206;
w6208 <= not w3540 and w5431;
w6209 <= not w2947 and w4870;
w6210 <= not w3474 and w5342;
w6211 <= not w6209 and not w6210;
w6212 <= not w6208 and w6211;
w6213 <= not w4873 and w6212;
w6214 <= not w4019 and w6212;
w6215 <= not w6213 and not w6214;
w6216 <= a(20) and not w6215;
w6217 <= not a(20) and w6215;
w6218 <= not w6216 and not w6217;
w6219 <= w6207 and not w6218;
w6220 <= w6133 and not w6145;
w6221 <= not w6144 and not w6145;
w6222 <= not w6220 and not w6221;
w6223 <= w6117 and not w6129;
w6224 <= not w6128 and not w6129;
w6225 <= not w6223 and not w6224;
w6226 <= w5934 and w6110;
w6227 <= not w6111 and not w6226;
w6228 <= not w1113 and w3819;
w6229 <= not w1299 and w3902;
w6230 <= not w1170 and w3981;
w6231 <= not w6229 and not w6230;
w6232 <= not w6228 and w6231;
w6233 <= not w3985 and w6232;
w6234 <= not w4796 and w6232;
w6235 <= not w6233 and not w6234;
w6236 <= a(26) and not w6235;
w6237 <= not a(26) and w6235;
w6238 <= not w6236 and not w6237;
w6239 <= w6227 and not w6238;
w6240 <= not w6105 and not w6109;
w6241 <= not w6108 and not w6109;
w6242 <= not w6240 and not w6241;
w6243 <= not w1507 and w3392;
w6244 <= not w1714 and w3477;
w6245 <= not w1600 and w3541;
w6246 <= not w6244 and not w6245;
w6247 <= not w6243 and w6246;
w6248 <= not w3303 and w6247;
w6249 <= not w5496 and w6247;
w6250 <= not w6248 and not w6249;
w6251 <= a(29) and not w6250;
w6252 <= not a(29) and w6250;
w6253 <= not w6251 and not w6252;
w6254 <= not w6242 and not w6253;
w6255 <= w6242 and w6253;
w6256 <= not w6254 and not w6255;
w6257 <= not w1170 and w3819;
w6258 <= not w1407 and w3902;
w6259 <= not w1299 and w3981;
w6260 <= not w6258 and not w6259;
w6261 <= not w6257 and w6260;
w6262 <= w3985 and w4783;
w6263 <= w6261 and not w6262;
w6264 <= a(26) and not w6263;
w6265 <= a(26) and not w6264;
w6266 <= not w6263 and not w6264;
w6267 <= not w6265 and not w6266;
w6268 <= w6256 and not w6267;
w6269 <= not w6254 and not w6268;
w6270 <= not w6227 and w6238;
w6271 <= not w6239 and not w6270;
w6272 <= not w6269 and w6271;
w6273 <= not w6239 and not w6272;
w6274 <= not w6225 and not w6273;
w6275 <= w6225 and w6273;
w6276 <= not w6274 and not w6275;
w6277 <= not w645 and w4629;
w6278 <= not w893 and w4468;
w6279 <= not w802 and w4539;
w6280 <= not w6278 and not w6279;
w6281 <= not w6277 and w6280;
w6282 <= w4114 and w4471;
w6283 <= w6281 and not w6282;
w6284 <= a(23) and not w6283;
w6285 <= a(23) and not w6284;
w6286 <= not w6283 and not w6284;
w6287 <= not w6285 and not w6286;
w6288 <= w6276 and not w6287;
w6289 <= not w6274 and not w6288;
w6290 <= not w6222 and not w6289;
w6291 <= w6222 and w6289;
w6292 <= not w6290 and not w6291;
w6293 <= not w3474 and w5431;
w6294 <= not w327 and w4870;
w6295 <= not w2947 and w5342;
w6296 <= not w6294 and not w6295;
w6297 <= not w6293 and w6296;
w6298 <= w3650 and w4873;
w6299 <= w6297 and not w6298;
w6300 <= a(20) and not w6299;
w6301 <= a(20) and not w6300;
w6302 <= not w6299 and not w6300;
w6303 <= not w6301 and not w6302;
w6304 <= w6292 and not w6303;
w6305 <= not w6290 and not w6304;
w6306 <= not w6207 and w6218;
w6307 <= not w6219 and not w6306;
w6308 <= not w6305 and w6307;
w6309 <= not w6219 and not w6308;
w6310 <= not w6205 and not w6309;
w6311 <= w6205 and w6309;
w6312 <= not w6310 and not w6311;
w6313 <= not w3980 and w6168;
w6314 <= not w3740 and w5598;
w6315 <= not w3899 and w5874;
w6316 <= not w6314 and not w6315;
w6317 <= not w6313 and w6316;
w6318 <= w4412 and w5601;
w6319 <= w6317 and not w6318;
w6320 <= a(17) and not w6319;
w6321 <= a(17) and not w6320;
w6322 <= not w6319 and not w6320;
w6323 <= not w6321 and not w6322;
w6324 <= w6312 and not w6323;
w6325 <= not w6310 and not w6324;
w6326 <= a(11) and not a(12);
w6327 <= not a(11) and a(12);
w6328 <= not w6326 and not w6327;
w6329 <= a(13) and not a(14);
w6330 <= not a(13) and a(14);
w6331 <= not w6329 and not w6330;
w6332 <= not w6328 and not w6331;
w6333 <= not a(12) and a(13);
w6334 <= a(12) and not a(13);
w6335 <= not w6333 and not w6334;
w6336 <= w6328 and not w6331;
w6337 <= w6335 and w6336;
w6338 <= not w4450 and w6337;
w6339 <= not w6332 and not w6338;
w6340 <= not w4457 and not w6338;
w6341 <= not w6339 and not w6340;
w6342 <= a(14) and not w6341;
w6343 <= not a(14) and w6341;
w6344 <= not w6342 and not w6343;
w6345 <= not w6325 and not w6344;
w6346 <= w6167 and not w6180;
w6347 <= not w6179 and not w6180;
w6348 <= not w6346 and not w6347;
w6349 <= w6325 and w6344;
w6350 <= not w6345 and not w6349;
w6351 <= not w6348 and w6350;
w6352 <= not w6345 and not w6351;
w6353 <= not w6195 and not w6197;
w6354 <= not w6198 and not w6353;
w6355 <= not w6352 and w6354;
w6356 <= w6352 and not w6354;
w6357 <= not w6355 and not w6356;
w6358 <= not w6348 and not w6351;
w6359 <= w6350 and not w6351;
w6360 <= not w6358 and not w6359;
w6361 <= not w3899 and w6168;
w6362 <= not w3391 and w5598;
w6363 <= not w3740 and w5874;
w6364 <= not w6362 and not w6363;
w6365 <= not w6361 and w6364;
w6366 <= w4493 and w5601;
w6367 <= w6365 and not w6366;
w6368 <= a(17) and not w6367;
w6369 <= not w6367 and not w6368;
w6370 <= a(17) and not w6368;
w6371 <= not w6369 and not w6370;
w6372 <= w6305 and not w6307;
w6373 <= not w6308 and not w6372;
w6374 <= not w6371 and w6373;
w6375 <= not w6371 and not w6374;
w6376 <= w6373 and not w6374;
w6377 <= not w6375 and not w6376;
w6378 <= w6292 and not w6304;
w6379 <= not w6303 and not w6304;
w6380 <= not w6378 and not w6379;
w6381 <= w6276 and not w6288;
w6382 <= not w6287 and not w6288;
w6383 <= not w6381 and not w6382;
w6384 <= not w802 and w4629;
w6385 <= not w995 and w4468;
w6386 <= not w893 and w4539;
w6387 <= not w6385 and not w6386;
w6388 <= not w6384 and w6387;
w6389 <= w4139 and w4471;
w6390 <= w6388 and not w6389;
w6391 <= a(23) and not w6390;
w6392 <= not w6390 and not w6391;
w6393 <= a(23) and not w6391;
w6394 <= not w6392 and not w6393;
w6395 <= w6269 and not w6271;
w6396 <= not w6272 and not w6395;
w6397 <= not w6394 and w6396;
w6398 <= not w6394 and not w6397;
w6399 <= w6396 and not w6397;
w6400 <= not w6398 and not w6399;
w6401 <= w6256 and not w6268;
w6402 <= not w6267 and not w6268;
w6403 <= not w6401 and not w6402;
w6404 <= w6087 and not w6088;
w6405 <= not w6085 and not w6088;
w6406 <= not w6404 and not w6405;
w6407 <= not w6070 and not w6072;
w6408 <= not w5978 and w6073;
w6409 <= not w6407 and not w6408;
w6410 <= not w1992 and w2955;
w6411 <= not w2087 and w2963;
w6412 <= not w2124 and w2958;
w6413 <= w2795 and not w2797;
w6414 <= not w2798 and not w6413;
w6415 <= w10 and w6414;
w6416 <= not w6412 and not w6415;
w6417 <= not w6411 and w6416;
w6418 <= not w6410 and w6417;
w6419 <= not w6409 and not w6418;
w6420 <= not w6067 and not w6069;
w6421 <= not w6011 and w6070;
w6422 <= not w6420 and not w6421;
w6423 <= not w2087 and w2955;
w6424 <= not w2124 and w2963;
w6425 <= not w2226 and w2958;
w6426 <= w2791 and not w2793;
w6427 <= not w2794 and not w6426;
w6428 <= w10 and w6427;
w6429 <= not w6425 and not w6428;
w6430 <= not w6424 and w6429;
w6431 <= not w6423 and w6430;
w6432 <= not w6422 and not w6431;
w6433 <= not w6064 and not w6066;
w6434 <= not w6055 and w6067;
w6435 <= not w6433 and not w6434;
w6436 <= w2543 and w4292;
w6437 <= w4763 and w6436;
w6438 <= w4214 and w6437;
w6439 <= w1729 and w6438;
w6440 <= w1227 and w6439;
w6441 <= w809 and w6440;
w6442 <= w1074 and w6441;
w6443 <= w2928 and w6442;
w6444 <= w51 and w6443;
w6445 <= not w552 and w6444;
w6446 <= not w189 and w6445;
w6447 <= not w744 and w6446;
w6448 <= not w303 and w6447;
w6449 <= not w726 and w6448;
w6450 <= not w110 and w5106;
w6451 <= not w141 and w6450;
w6452 <= not w590 and w6451;
w6453 <= not w58 and not w453;
w6454 <= not w92 and w6453;
w6455 <= not w205 and w6454;
w6456 <= w3459 and w5710;
w6457 <= w626 and w6456;
w6458 <= w6455 and w6457;
w6459 <= w6452 and w6458;
w6460 <= w1644 and w6459;
w6461 <= w4340 and w6460;
w6462 <= w4310 and w6461;
w6463 <= w6449 and w6462;
w6464 <= w389 and w6463;
w6465 <= w666 and w6464;
w6466 <= w1413 and w6465;
w6467 <= not w71 and w6466;
w6468 <= not w183 and w6467;
w6469 <= not w233 and w6468;
w6470 <= not w208 and w6469;
w6471 <= not w371 and w6470;
w6472 <= not w2226 and w2955;
w6473 <= not w2323 and w2963;
w6474 <= not w2399 and w2958;
w6475 <= w2783 and not w2785;
w6476 <= not w2786 and not w6475;
w6477 <= w10 and w6476;
w6478 <= not w6474 and not w6477;
w6479 <= not w6473 and w6478;
w6480 <= not w6472 and w6479;
w6481 <= not w6471 and not w6480;
w6482 <= not w213 and not w331;
w6483 <= not w467 and w6482;
w6484 <= w4956 and w6483;
w6485 <= w1720 and w6484;
w6486 <= w1521 and w6485;
w6487 <= w4062 and w6486;
w6488 <= w2518 and w6487;
w6489 <= w35 and w6488;
w6490 <= not w602 and w6489;
w6491 <= not w576 and w6490;
w6492 <= not w124 and w6491;
w6493 <= not w42 and w6492;
w6494 <= not w712 and w6493;
w6495 <= not w499 and w6494;
w6496 <= not w16 and w6495;
w6497 <= w358 and not w997;
w6498 <= not w819 and w6497;
w6499 <= not w233 and w6498;
w6500 <= not w460 and w6499;
w6501 <= not w219 and w1063;
w6502 <= not w395 and w6501;
w6503 <= w1675 and w3351;
w6504 <= w2155 and w6503;
w6505 <= w6502 and w6504;
w6506 <= w1627 and w6505;
w6507 <= w6500 and w6506;
w6508 <= w812 and w6507;
w6509 <= w1644 and w6508;
w6510 <= w203 and w6509;
w6511 <= w4302 and w6510;
w6512 <= w6496 and w6511;
w6513 <= w4998 and w6512;
w6514 <= w385 and w6513;
w6515 <= w1696 and w6514;
w6516 <= not w129 and w6515;
w6517 <= not w86 and w6516;
w6518 <= not w210 and w6517;
w6519 <= not w108 and w6518;
w6520 <= not w428 and w6519;
w6521 <= not w135 and w6520;
w6522 <= not w2323 and w2955;
w6523 <= not w2399 and w2963;
w6524 <= not w2468 and w2958;
w6525 <= w2779 and not w2781;
w6526 <= not w2782 and not w6525;
w6527 <= w10 and w6526;
w6528 <= not w6524 and not w6527;
w6529 <= not w6523 and w6528;
w6530 <= not w6522 and w6529;
w6531 <= not w6521 and not w6530;
w6532 <= w853 and w2126;
w6533 <= w214 and w6532;
w6534 <= w35 and w6533;
w6535 <= not w224 and w6534;
w6536 <= not w738 and w6535;
w6537 <= not w181 and w6536;
w6538 <= not w401 and w6537;
w6539 <= not w607 and w6538;
w6540 <= not w263 and w450;
w6541 <= not w331 and w6540;
w6542 <= not w403 and w6541;
w6543 <= not w687 and w1759;
w6544 <= not w651 and w6543;
w6545 <= not w424 and w6544;
w6546 <= w1359 and w1523;
w6547 <= w6545 and w6546;
w6548 <= w6542 and w6547;
w6549 <= w5083 and w6548;
w6550 <= w655 and w6549;
w6551 <= w569 and w6550;
w6552 <= not w333 and w6551;
w6553 <= not w87 and w6552;
w6554 <= not w289 and w6553;
w6555 <= not w712 and w6554;
w6556 <= not w351 and w6555;
w6557 <= not w303 and w6556;
w6558 <= not w867 and w6557;
w6559 <= not w207 and w6558;
w6560 <= not w647 and w6559;
w6561 <= not w493 and w2104;
w6562 <= not w274 and w6561;
w6563 <= not w262 and w6562;
w6564 <= w107 and w1432;
w6565 <= w6563 and w6564;
w6566 <= w2305 and w6565;
w6567 <= w3703 and w6566;
w6568 <= w5159 and w6567;
w6569 <= w6560 and w6568;
w6570 <= w6539 and w6569;
w6571 <= not w288 and w6570;
w6572 <= not w302 and w6571;
w6573 <= not w760 and w6572;
w6574 <= not w126 and w6573;
w6575 <= not w160 and w6574;
w6576 <= not w371 and w6575;
w6577 <= not w2399 and w2955;
w6578 <= not w2468 and w2963;
w6579 <= not w2506 and w2958;
w6580 <= w2775 and not w2777;
w6581 <= not w2778 and not w6580;
w6582 <= w10 and w6581;
w6583 <= not w6579 and not w6582;
w6584 <= not w6578 and w6583;
w6585 <= not w6577 and w6584;
w6586 <= not w6576 and not w6585;
w6587 <= w3249 and w3484;
w6588 <= w3344 and w6587;
w6589 <= w1040 and w6588;
w6590 <= w1458 and w6589;
w6591 <= not w58 and w6590;
w6592 <= not w362 and w6591;
w6593 <= not w264 and w6592;
w6594 <= not w263 and w6593;
w6595 <= not w337 and w6594;
w6596 <= not w365 and w6595;
w6597 <= not w275 and w6596;
w6598 <= not w293 and not w453;
w6599 <= not w363 and w6598;
w6600 <= w762 and w6599;
w6601 <= not w241 and w6600;
w6602 <= not w93 and w6601;
w6603 <= not w96 and not w466;
w6604 <= not w239 and w6603;
w6605 <= not w157 and w6604;
w6606 <= not w215 and w539;
w6607 <= not w267 and w6606;
w6608 <= w1513 and w6607;
w6609 <= w4204 and w6608;
w6610 <= w6605 and w6609;
w6611 <= w6602 and w6610;
w6612 <= w2193 and w6611;
w6613 <= w6597 and w6612;
w6614 <= w740 and w6613;
w6615 <= w2508 and w6614;
w6616 <= w1466 and w6615;
w6617 <= w1076 and w6616;
w6618 <= w913 and w6617;
w6619 <= w1096 and w6618;
w6620 <= not w288 and w6619;
w6621 <= not w234 and w6620;
w6622 <= not w425 and w6621;
w6623 <= not w503 and w6622;
w6624 <= not w99 and w6623;
w6625 <= not w558 and w6624;
w6626 <= not w2468 and w2955;
w6627 <= not w2506 and w2963;
w6628 <= not w2609 and w2958;
w6629 <= w2771 and not w2773;
w6630 <= not w2774 and not w6629;
w6631 <= w10 and w6630;
w6632 <= not w6628 and not w6631;
w6633 <= not w6627 and w6632;
w6634 <= not w6626 and w6633;
w6635 <= not w6625 and not w6634;
w6636 <= w235 and not w236;
w6637 <= not w1037 and w6636;
w6638 <= not w138 and w6637;
w6639 <= not w261 and w6638;
w6640 <= not w222 and w6639;
w6641 <= not w80 and not w99;
w6642 <= not w471 and w6641;
w6643 <= w1463 and w1552;
w6644 <= w2568 and w6643;
w6645 <= w3821 and w6644;
w6646 <= not w650 and w6645;
w6647 <= not w307 and w6646;
w6648 <= not w301 and w6647;
w6649 <= not w568 and w6648;
w6650 <= not w67 and w3516;
w6651 <= not w136 and w6650;
w6652 <= not w492 and w2024;
w6653 <= w2358 and w6652;
w6654 <= w6651 and w6653;
w6655 <= w832 and w6654;
w6656 <= w1411 and w6655;
w6657 <= w600 and w6656;
w6658 <= w6649 and w6657;
w6659 <= w1466 and w6658;
w6660 <= w761 and w6659;
w6661 <= w162 and w6660;
w6662 <= not w453 and w6661;
w6663 <= not w1036 and w6662;
w6664 <= not w127 and w6663;
w6665 <= not w867 and w6664;
w6666 <= not w409 and w6665;
w6667 <= not w467 and w6666;
w6668 <= not w168 and w820;
w6669 <= not w79 and w6668;
w6670 <= w1156 and w6669;
w6671 <= w1550 and w6670;
w6672 <= w2567 and w6671;
w6673 <= w1389 and w6672;
w6674 <= w6667 and w6673;
w6675 <= w6642 and w6674;
w6676 <= w1956 and w6675;
w6677 <= w6640 and w6676;
w6678 <= not w266 and w6677;
w6679 <= not w207 and w6678;
w6680 <= not w386 and w6679;
w6681 <= not w1039 and w6680;
w6682 <= not w497 and w6681;
w6683 <= not w590 and w6682;
w6684 <= w235 and w2639;
w6685 <= not w46 and w6684;
w6686 <= not w1241 and w6685;
w6687 <= not w309 and w6686;
w6688 <= not w498 and w6687;
w6689 <= not w266 and w6688;
w6690 <= not w306 and w6689;
w6691 <= w5136 and w5728;
w6692 <= w711 and w6691;
w6693 <= w402 and w6692;
w6694 <= w6605 and w6693;
w6695 <= w2673 and w6694;
w6696 <= w808 and w6695;
w6697 <= w1945 and w6696;
w6698 <= w1759 and w6697;
w6699 <= w2008 and w6698;
w6700 <= not w651 and w6699;
w6701 <= not w357 and w6700;
w6702 <= not w329 and w6701;
w6703 <= not w538 and w6702;
w6704 <= not w818 and w6703;
w6705 <= not w1062 and w3571;
w6706 <= not w568 and w6705;
w6707 <= w670 and w1521;
w6708 <= w6706 and w6707;
w6709 <= w4083 and w6708;
w6710 <= w2039 and w6709;
w6711 <= w6704 and w6710;
w6712 <= w6690 and w6711;
w6713 <= w445 and w6712;
w6714 <= w1603 and w6713;
w6715 <= w223 and w6714;
w6716 <= w804 and w6715;
w6717 <= w2401 and w6716;
w6718 <= w745 and w6717;
w6719 <= not w171 and w6718;
w6720 <= not w224 and w6719;
w6721 <= not w189 and w6720;
w6722 <= not w446 and w6721;
w6723 <= not w138 and w6722;
w6724 <= not w302 and w6723;
w6725 <= not w712 and w6724;
w6726 <= not w181 and w6725;
w6727 <= not w2609 and w2955;
w6728 <= not w2671 and w2963;
w6729 <= not w2764 and w2958;
w6730 <= not w2671 and w2764;
w6731 <= w2609 and not w6730;
w6732 <= w2672 and w2764;
w6733 <= not w6731 and not w6732;
w6734 <= w10 and w6733;
w6735 <= not w6729 and not w6734;
w6736 <= not w6728 and w6735;
w6737 <= not w6727 and w6736;
w6738 <= not w6726 and not w6737;
w6739 <= not w6683 and w6738;
w6740 <= w2767 and not w2769;
w6741 <= not w2770 and not w6740;
w6742 <= w10 and w6741;
w6743 <= not w2506 and w2955;
w6744 <= not w2671 and w2958;
w6745 <= not w2609 and w2963;
w6746 <= not w6744 and not w6745;
w6747 <= not w6743 and w6746;
w6748 <= not w6742 and w6747;
w6749 <= w6683 and not w6738;
w6750 <= not w6739 and not w6749;
w6751 <= not w6748 and w6750;
w6752 <= not w6739 and not w6751;
w6753 <= not w6625 and not w6635;
w6754 <= not w6634 and not w6635;
w6755 <= not w6753 and not w6754;
w6756 <= not w6752 and not w6755;
w6757 <= not w6635 and not w6756;
w6758 <= not w6576 and not w6586;
w6759 <= not w6585 and not w6586;
w6760 <= not w6758 and not w6759;
w6761 <= not w6757 and not w6760;
w6762 <= not w6586 and not w6761;
w6763 <= not w6521 and not w6531;
w6764 <= not w6530 and not w6531;
w6765 <= not w6763 and not w6764;
w6766 <= not w6762 and not w6765;
w6767 <= not w6531 and not w6766;
w6768 <= not w6471 and not w6481;
w6769 <= not w6480 and not w6481;
w6770 <= not w6768 and not w6769;
w6771 <= not w6767 and not w6770;
w6772 <= not w6481 and not w6771;
w6773 <= not w6435 and not w6772;
w6774 <= w6435 and w6772;
w6775 <= not w6773 and not w6774;
w6776 <= not w1927 and w3392;
w6777 <= not w2087 and w3477;
w6778 <= not w1992 and w3541;
w6779 <= not w6777 and not w6778;
w6780 <= not w6776 and w6779;
w6781 <= not w3303 and w6780;
w6782 <= not w6078 and w6780;
w6783 <= not w6781 and not w6782;
w6784 <= a(29) and not w6783;
w6785 <= not a(29) and w6783;
w6786 <= not w6784 and not w6785;
w6787 <= w6775 and not w6786;
w6788 <= not w6773 and not w6787;
w6789 <= not w6422 and not w6432;
w6790 <= not w6431 and not w6432;
w6791 <= not w6789 and not w6790;
w6792 <= not w6788 and not w6791;
w6793 <= not w6432 and not w6792;
w6794 <= not w6409 and not w6419;
w6795 <= not w6418 and not w6419;
w6796 <= not w6794 and not w6795;
w6797 <= not w6793 and not w6796;
w6798 <= not w6419 and not w6797;
w6799 <= not w6406 and not w6798;
w6800 <= w6406 and w6798;
w6801 <= not w6799 and not w6800;
w6802 <= not w1714 and w3392;
w6803 <= not w1848 and w3477;
w6804 <= not w1812 and w3541;
w6805 <= not w6803 and not w6804;
w6806 <= not w6802 and w6805;
w6807 <= w3303 and w5786;
w6808 <= w6806 and not w6807;
w6809 <= a(29) and not w6808;
w6810 <= a(29) and not w6809;
w6811 <= not w6808 and not w6809;
w6812 <= not w6810 and not w6811;
w6813 <= w6801 and not w6812;
w6814 <= not w6799 and not w6813;
w6815 <= not w6092 and w6103;
w6816 <= not w6104 and not w6815;
w6817 <= not w6814 and w6816;
w6818 <= w6814 and not w6816;
w6819 <= not w6817 and not w6818;
w6820 <= not w1299 and w3819;
w6821 <= not w1507 and w3902;
w6822 <= not w1407 and w3981;
w6823 <= not w6821 and not w6822;
w6824 <= not w6820 and w6823;
w6825 <= w3985 and w5049;
w6826 <= w6824 and not w6825;
w6827 <= a(26) and not w6826;
w6828 <= a(26) and not w6827;
w6829 <= not w6826 and not w6827;
w6830 <= not w6828 and not w6829;
w6831 <= w6819 and not w6830;
w6832 <= not w6817 and not w6831;
w6833 <= not w6403 and not w6832;
w6834 <= w6403 and w6832;
w6835 <= not w6833 and not w6834;
w6836 <= not w893 and w4629;
w6837 <= not w1113 and w4468;
w6838 <= not w995 and w4539;
w6839 <= not w6837 and not w6838;
w6840 <= not w6836 and w6839;
w6841 <= w4471 and w4568;
w6842 <= w6840 and not w6841;
w6843 <= a(23) and not w6842;
w6844 <= a(23) and not w6843;
w6845 <= not w6842 and not w6843;
w6846 <= not w6844 and not w6845;
w6847 <= w6835 and not w6846;
w6848 <= not w6833 and not w6847;
w6849 <= not w6400 and not w6848;
w6850 <= not w6397 and not w6849;
w6851 <= not w6383 and not w6850;
w6852 <= w6383 and w6850;
w6853 <= not w6851 and not w6852;
w6854 <= not w2947 and w5431;
w6855 <= not w522 and w4870;
w6856 <= not w327 and w5342;
w6857 <= not w6855 and not w6856;
w6858 <= not w6854 and w6857;
w6859 <= w2953 and w4873;
w6860 <= w6858 and not w6859;
w6861 <= a(20) and not w6860;
w6862 <= a(20) and not w6861;
w6863 <= not w6860 and not w6861;
w6864 <= not w6862 and not w6863;
w6865 <= w6853 and not w6864;
w6866 <= not w6851 and not w6865;
w6867 <= not w6380 and not w6866;
w6868 <= w6380 and w6866;
w6869 <= not w6867 and not w6868;
w6870 <= not w3740 and w6168;
w6871 <= not w3540 and w5598;
w6872 <= not w3391 and w5874;
w6873 <= not w6871 and not w6872;
w6874 <= not w6870 and w6873;
w6875 <= w3753 and w5601;
w6876 <= w6874 and not w6875;
w6877 <= a(17) and not w6876;
w6878 <= a(17) and not w6877;
w6879 <= not w6876 and not w6877;
w6880 <= not w6878 and not w6879;
w6881 <= w6869 and not w6880;
w6882 <= not w6867 and not w6881;
w6883 <= not w6377 and not w6882;
w6884 <= not w6374 and not w6883;
w6885 <= not w3812 and w6337;
w6886 <= w6328 and not w6335;
w6887 <= not w4450 and w6886;
w6888 <= not w6885 and not w6887;
w6889 <= not w6332 and w6888;
w6890 <= not w4544 and w6888;
w6891 <= not w6889 and not w6890;
w6892 <= a(14) and not w6891;
w6893 <= not a(14) and w6891;
w6894 <= not w6892 and not w6893;
w6895 <= not w6884 and not w6894;
w6896 <= w6312 and not w6324;
w6897 <= not w6323 and not w6324;
w6898 <= not w6896 and not w6897;
w6899 <= w6884 and w6894;
w6900 <= not w6895 and not w6899;
w6901 <= not w6898 and w6900;
w6902 <= not w6895 and not w6901;
w6903 <= not w6360 and not w6902;
w6904 <= w6360 and w6902;
w6905 <= not w6903 and not w6904;
w6906 <= w6869 and not w6881;
w6907 <= not w6880 and not w6881;
w6908 <= not w6906 and not w6907;
w6909 <= w6853 and not w6865;
w6910 <= not w6864 and not w6865;
w6911 <= not w6909 and not w6910;
w6912 <= w6400 and w6848;
w6913 <= not w6849 and not w6912;
w6914 <= not w327 and w5431;
w6915 <= not w645 and w4870;
w6916 <= not w522 and w5342;
w6917 <= not w6915 and not w6916;
w6918 <= not w6914 and w6917;
w6919 <= not w4873 and w6918;
w6920 <= not w3282 and w6918;
w6921 <= not w6919 and not w6920;
w6922 <= a(20) and not w6921;
w6923 <= not a(20) and w6921;
w6924 <= not w6922 and not w6923;
w6925 <= w6913 and not w6924;
w6926 <= w6835 and not w6847;
w6927 <= not w6846 and not w6847;
w6928 <= not w6926 and not w6927;
w6929 <= w6819 and not w6831;
w6930 <= not w6830 and not w6831;
w6931 <= not w6929 and not w6930;
w6932 <= w6801 and not w6813;
w6933 <= not w6812 and not w6813;
w6934 <= not w6932 and not w6933;
w6935 <= not w1407 and w3819;
w6936 <= not w1600 and w3902;
w6937 <= not w1507 and w3981;
w6938 <= not w6936 and not w6937;
w6939 <= not w6935 and w6938;
w6940 <= not w3985 and w6939;
w6941 <= not w5074 and w6939;
w6942 <= not w6940 and not w6941;
w6943 <= a(26) and not w6942;
w6944 <= not a(26) and w6942;
w6945 <= not w6943 and not w6944;
w6946 <= not w6934 and not w6945;
w6947 <= not w6793 and not w6797;
w6948 <= not w6796 and not w6797;
w6949 <= not w6947 and not w6948;
w6950 <= not w1812 and w3392;
w6951 <= not w1927 and w3477;
w6952 <= not w1848 and w3541;
w6953 <= not w6951 and not w6952;
w6954 <= not w6950 and w6953;
w6955 <= not w3303 and w6954;
w6956 <= not w5942 and w6954;
w6957 <= not w6955 and not w6956;
w6958 <= a(29) and not w6957;
w6959 <= not a(29) and w6957;
w6960 <= not w6958 and not w6959;
w6961 <= not w6949 and not w6960;
w6962 <= w6949 and w6960;
w6963 <= not w6961 and not w6962;
w6964 <= not w1507 and w3819;
w6965 <= not w1714 and w3902;
w6966 <= not w1600 and w3981;
w6967 <= not w6965 and not w6966;
w6968 <= not w6964 and w6967;
w6969 <= w3985 and w5496;
w6970 <= w6968 and not w6969;
w6971 <= a(26) and not w6970;
w6972 <= a(26) and not w6971;
w6973 <= not w6970 and not w6971;
w6974 <= not w6972 and not w6973;
w6975 <= w6963 and not w6974;
w6976 <= not w6961 and not w6975;
w6977 <= w6934 and w6945;
w6978 <= not w6946 and not w6977;
w6979 <= not w6976 and w6978;
w6980 <= not w6946 and not w6979;
w6981 <= not w6931 and not w6980;
w6982 <= w6931 and w6980;
w6983 <= not w6981 and not w6982;
w6984 <= not w995 and w4629;
w6985 <= not w1170 and w4468;
w6986 <= not w1113 and w4539;
w6987 <= not w6985 and not w6986;
w6988 <= not w6984 and w6987;
w6989 <= w4364 and w4471;
w6990 <= w6988 and not w6989;
w6991 <= a(23) and not w6990;
w6992 <= a(23) and not w6991;
w6993 <= not w6990 and not w6991;
w6994 <= not w6992 and not w6993;
w6995 <= w6983 and not w6994;
w6996 <= not w6981 and not w6995;
w6997 <= not w6928 and not w6996;
w6998 <= w6928 and w6996;
w6999 <= not w6997 and not w6998;
w7000 <= not w522 and w5431;
w7001 <= not w802 and w4870;
w7002 <= not w645 and w5342;
w7003 <= not w7001 and not w7002;
w7004 <= not w7000 and w7003;
w7005 <= w3266 and w4873;
w7006 <= w7004 and not w7005;
w7007 <= a(20) and not w7006;
w7008 <= a(20) and not w7007;
w7009 <= not w7006 and not w7007;
w7010 <= not w7008 and not w7009;
w7011 <= w6999 and not w7010;
w7012 <= not w6997 and not w7011;
w7013 <= not w6913 and w6924;
w7014 <= not w6925 and not w7013;
w7015 <= not w7012 and w7014;
w7016 <= not w6925 and not w7015;
w7017 <= not w6911 and not w7016;
w7018 <= w6911 and w7016;
w7019 <= not w7017 and not w7018;
w7020 <= not w3391 and w6168;
w7021 <= not w3474 and w5598;
w7022 <= not w3540 and w5874;
w7023 <= not w7021 and not w7022;
w7024 <= not w7020 and w7023;
w7025 <= w3562 and w5601;
w7026 <= w7024 and not w7025;
w7027 <= a(17) and not w7026;
w7028 <= a(17) and not w7027;
w7029 <= not w7026 and not w7027;
w7030 <= not w7028 and not w7029;
w7031 <= w7019 and not w7030;
w7032 <= not w7017 and not w7031;
w7033 <= not w6908 and not w7032;
w7034 <= w6908 and w7032;
w7035 <= not w7033 and not w7034;
w7036 <= not w6328 and w6331;
w7037 <= not w3812 and w7036;
w7038 <= not w3899 and w6337;
w7039 <= not w3980 and w6886;
w7040 <= not w7038 and not w7039;
w7041 <= not w7037 and w7040;
w7042 <= w4002 and w6332;
w7043 <= w7041 and not w7042;
w7044 <= a(14) and not w7043;
w7045 <= a(14) and not w7044;
w7046 <= not w7043 and not w7044;
w7047 <= not w7045 and not w7046;
w7048 <= w7035 and not w7047;
w7049 <= not w7033 and not w7048;
w7050 <= not w4450 and w7036;
w7051 <= not w3980 and w6337;
w7052 <= not w3812 and w6886;
w7053 <= not w7051 and not w7052;
w7054 <= not w7050 and w7053;
w7055 <= not w6332 and w7054;
w7056 <= not w4650 and w7054;
w7057 <= not w7055 and not w7056;
w7058 <= a(14) and not w7057;
w7059 <= not a(14) and w7057;
w7060 <= not w7058 and not w7059;
w7061 <= not w7049 and not w7060;
w7062 <= w6377 and w6882;
w7063 <= not w6883 and not w7062;
w7064 <= not w7049 and not w7061;
w7065 <= not w7060 and not w7061;
w7066 <= not w7064 and not w7065;
w7067 <= w7063 and not w7066;
w7068 <= not w7061 and not w7067;
w7069 <= w6898 and not w6900;
w7070 <= not w6901 and not w7069;
w7071 <= not w7068 and w7070;
w7072 <= w7019 and not w7031;
w7073 <= not w7030 and not w7031;
w7074 <= not w7072 and not w7073;
w7075 <= not w3540 and w6168;
w7076 <= not w2947 and w5598;
w7077 <= not w3474 and w5874;
w7078 <= not w7076 and not w7077;
w7079 <= not w7075 and w7078;
w7080 <= w4019 and w5601;
w7081 <= w7079 and not w7080;
w7082 <= a(17) and not w7081;
w7083 <= not w7081 and not w7082;
w7084 <= a(17) and not w7082;
w7085 <= not w7083 and not w7084;
w7086 <= w7012 and not w7014;
w7087 <= not w7015 and not w7086;
w7088 <= not w7085 and w7087;
w7089 <= not w7085 and not w7088;
w7090 <= w7087 and not w7088;
w7091 <= not w7089 and not w7090;
w7092 <= w6999 and not w7011;
w7093 <= not w7010 and not w7011;
w7094 <= not w7092 and not w7093;
w7095 <= w6983 and not w6995;
w7096 <= not w6994 and not w6995;
w7097 <= not w7095 and not w7096;
w7098 <= not w1113 and w4629;
w7099 <= not w1299 and w4468;
w7100 <= not w1170 and w4539;
w7101 <= not w7099 and not w7100;
w7102 <= not w7098 and w7101;
w7103 <= w4471 and w4796;
w7104 <= w7102 and not w7103;
w7105 <= a(23) and not w7104;
w7106 <= not w7104 and not w7105;
w7107 <= a(23) and not w7105;
w7108 <= not w7106 and not w7107;
w7109 <= w6976 and not w6978;
w7110 <= not w6979 and not w7109;
w7111 <= not w7108 and w7110;
w7112 <= not w7108 and not w7111;
w7113 <= w7110 and not w7111;
w7114 <= not w7112 and not w7113;
w7115 <= w6963 and not w6975;
w7116 <= not w6974 and not w6975;
w7117 <= not w7115 and not w7116;
w7118 <= not w6788 and not w6792;
w7119 <= not w6791 and not w6792;
w7120 <= not w7118 and not w7119;
w7121 <= not w1848 and w3392;
w7122 <= not w1992 and w3477;
w7123 <= not w1927 and w3541;
w7124 <= not w7122 and not w7123;
w7125 <= not w7121 and w7124;
w7126 <= not w3303 and w7125;
w7127 <= not w5769 and w7125;
w7128 <= not w7126 and not w7127;
w7129 <= a(29) and not w7128;
w7130 <= not a(29) and w7128;
w7131 <= not w7129 and not w7130;
w7132 <= not w7120 and not w7131;
w7133 <= w7120 and w7131;
w7134 <= not w7132 and not w7133;
w7135 <= not w1600 and w3819;
w7136 <= not w1812 and w3902;
w7137 <= not w1714 and w3981;
w7138 <= not w7136 and not w7137;
w7139 <= not w7135 and w7138;
w7140 <= w3985 and w5263;
w7141 <= w7139 and not w7140;
w7142 <= a(26) and not w7141;
w7143 <= a(26) and not w7142;
w7144 <= not w7141 and not w7142;
w7145 <= not w7143 and not w7144;
w7146 <= w7134 and not w7145;
w7147 <= not w7132 and not w7146;
w7148 <= not w7117 and not w7147;
w7149 <= w7117 and w7147;
w7150 <= not w7148 and not w7149;
w7151 <= not w1170 and w4629;
w7152 <= not w1407 and w4468;
w7153 <= not w1299 and w4539;
w7154 <= not w7152 and not w7153;
w7155 <= not w7151 and w7154;
w7156 <= w4471 and w4783;
w7157 <= w7155 and not w7156;
w7158 <= a(23) and not w7157;
w7159 <= a(23) and not w7158;
w7160 <= not w7157 and not w7158;
w7161 <= not w7159 and not w7160;
w7162 <= w7150 and not w7161;
w7163 <= not w7148 and not w7162;
w7164 <= not w7114 and not w7163;
w7165 <= not w7111 and not w7164;
w7166 <= not w7097 and not w7165;
w7167 <= w7097 and w7165;
w7168 <= not w7166 and not w7167;
w7169 <= not w645 and w5431;
w7170 <= not w893 and w4870;
w7171 <= not w802 and w5342;
w7172 <= not w7170 and not w7171;
w7173 <= not w7169 and w7172;
w7174 <= w4114 and w4873;
w7175 <= w7173 and not w7174;
w7176 <= a(20) and not w7175;
w7177 <= a(20) and not w7176;
w7178 <= not w7175 and not w7176;
w7179 <= not w7177 and not w7178;
w7180 <= w7168 and not w7179;
w7181 <= not w7166 and not w7180;
w7182 <= not w7094 and not w7181;
w7183 <= w7094 and w7181;
w7184 <= not w7182 and not w7183;
w7185 <= not w3474 and w6168;
w7186 <= not w327 and w5598;
w7187 <= not w2947 and w5874;
w7188 <= not w7186 and not w7187;
w7189 <= not w7185 and w7188;
w7190 <= w3650 and w5601;
w7191 <= w7189 and not w7190;
w7192 <= a(17) and not w7191;
w7193 <= a(17) and not w7192;
w7194 <= not w7191 and not w7192;
w7195 <= not w7193 and not w7194;
w7196 <= w7184 and not w7195;
w7197 <= not w7182 and not w7196;
w7198 <= not w7091 and not w7197;
w7199 <= not w7088 and not w7198;
w7200 <= not w7074 and not w7199;
w7201 <= w7074 and w7199;
w7202 <= not w7200 and not w7201;
w7203 <= not w3980 and w7036;
w7204 <= not w3740 and w6337;
w7205 <= not w3899 and w6886;
w7206 <= not w7204 and not w7205;
w7207 <= not w7203 and w7206;
w7208 <= w4412 and w6332;
w7209 <= w7207 and not w7208;
w7210 <= a(14) and not w7209;
w7211 <= a(14) and not w7210;
w7212 <= not w7209 and not w7210;
w7213 <= not w7211 and not w7212;
w7214 <= w7202 and not w7213;
w7215 <= not w7200 and not w7214;
w7216 <= not a(9) and a(10);
w7217 <= a(9) and not a(10);
w7218 <= not w7216 and not w7217;
w7219 <= a(10) and not a(11);
w7220 <= not a(10) and a(11);
w7221 <= not w7219 and not w7220;
w7222 <= a(8) and not a(9);
w7223 <= not a(8) and a(9);
w7224 <= not w7222 and not w7223;
w7225 <= not w7221 and w7224;
w7226 <= w7218 and w7225;
w7227 <= not w4450 and w7226;
w7228 <= not w4457 and not w7227;
w7229 <= not w7221 and not w7224;
w7230 <= not w7227 and not w7229;
w7231 <= not w7228 and not w7230;
w7232 <= a(11) and not w7231;
w7233 <= not a(11) and w7231;
w7234 <= not w7232 and not w7233;
w7235 <= not w7215 and not w7234;
w7236 <= w7035 and not w7048;
w7237 <= not w7047 and not w7048;
w7238 <= not w7236 and not w7237;
w7239 <= w7215 and w7234;
w7240 <= not w7235 and not w7239;
w7241 <= not w7238 and w7240;
w7242 <= not w7235 and not w7241;
w7243 <= not w7063 and not w7065;
w7244 <= not w7064 and w7243;
w7245 <= not w7067 and not w7244;
w7246 <= not w7242 and w7245;
w7247 <= not w7238 and not w7241;
w7248 <= w7240 and not w7241;
w7249 <= not w7247 and not w7248;
w7250 <= w7091 and w7197;
w7251 <= not w7198 and not w7250;
w7252 <= not w3899 and w7036;
w7253 <= not w3391 and w6337;
w7254 <= not w3740 and w6886;
w7255 <= not w7253 and not w7254;
w7256 <= not w7252 and w7255;
w7257 <= not w6332 and w7256;
w7258 <= not w4493 and w7256;
w7259 <= not w7257 and not w7258;
w7260 <= a(14) and not w7259;
w7261 <= not a(14) and w7259;
w7262 <= not w7260 and not w7261;
w7263 <= w7251 and not w7262;
w7264 <= w7184 and not w7196;
w7265 <= not w7195 and not w7196;
w7266 <= not w7264 and not w7265;
w7267 <= w7168 and not w7180;
w7268 <= not w7179 and not w7180;
w7269 <= not w7267 and not w7268;
w7270 <= w7114 and w7163;
w7271 <= not w7164 and not w7270;
w7272 <= not w802 and w5431;
w7273 <= not w995 and w4870;
w7274 <= not w893 and w5342;
w7275 <= not w7273 and not w7274;
w7276 <= not w7272 and w7275;
w7277 <= not w4873 and w7276;
w7278 <= not w4139 and w7276;
w7279 <= not w7277 and not w7278;
w7280 <= a(20) and not w7279;
w7281 <= not a(20) and w7279;
w7282 <= not w7280 and not w7281;
w7283 <= w7271 and not w7282;
w7284 <= w7150 and not w7162;
w7285 <= not w7161 and not w7162;
w7286 <= not w7284 and not w7285;
w7287 <= w7134 and not w7146;
w7288 <= not w7145 and not w7146;
w7289 <= not w7287 and not w7288;
w7290 <= not w6767 and not w6771;
w7291 <= not w6770 and not w6771;
w7292 <= not w7290 and not w7291;
w7293 <= not w1992 and w3392;
w7294 <= not w2124 and w3477;
w7295 <= not w2087 and w3541;
w7296 <= not w7294 and not w7295;
w7297 <= not w7293 and w7296;
w7298 <= not w3303 and w7297;
w7299 <= not w6414 and w7297;
w7300 <= not w7298 and not w7299;
w7301 <= a(29) and not w7300;
w7302 <= not a(29) and w7300;
w7303 <= not w7301 and not w7302;
w7304 <= not w7292 and not w7303;
w7305 <= not w6762 and not w6766;
w7306 <= not w6765 and not w6766;
w7307 <= not w7305 and not w7306;
w7308 <= not w2087 and w3392;
w7309 <= not w2226 and w3477;
w7310 <= not w2124 and w3541;
w7311 <= not w7309 and not w7310;
w7312 <= not w7308 and w7311;
w7313 <= not w3303 and w7312;
w7314 <= not w6427 and w7312;
w7315 <= not w7313 and not w7314;
w7316 <= a(29) and not w7315;
w7317 <= not a(29) and w7315;
w7318 <= not w7316 and not w7317;
w7319 <= not w7307 and not w7318;
w7320 <= not w2124 and w3392;
w7321 <= not w2323 and w3477;
w7322 <= not w2226 and w3541;
w7323 <= not w7321 and not w7322;
w7324 <= not w7320 and w7323;
w7325 <= w3303 and w6057;
w7326 <= w7324 and not w7325;
w7327 <= a(29) and not w7326;
w7328 <= not w7326 and not w7327;
w7329 <= a(29) and not w7327;
w7330 <= not w7328 and not w7329;
w7331 <= not w6757 and not w6761;
w7332 <= not w6760 and not w6761;
w7333 <= not w7331 and not w7332;
w7334 <= not w7330 and not w7333;
w7335 <= not w7330 and not w7334;
w7336 <= not w7333 and not w7334;
w7337 <= not w7335 and not w7336;
w7338 <= not w2226 and w3392;
w7339 <= not w2399 and w3477;
w7340 <= not w2323 and w3541;
w7341 <= not w7339 and not w7340;
w7342 <= not w7338 and w7341;
w7343 <= w3303 and w6476;
w7344 <= w7342 and not w7343;
w7345 <= a(29) and not w7344;
w7346 <= not w7344 and not w7345;
w7347 <= a(29) and not w7345;
w7348 <= not w7346 and not w7347;
w7349 <= not w6752 and not w6756;
w7350 <= not w6755 and not w6756;
w7351 <= not w7349 and not w7350;
w7352 <= not w7348 and not w7351;
w7353 <= not w7348 and not w7352;
w7354 <= not w7351 and not w7352;
w7355 <= not w7353 and not w7354;
w7356 <= not w2323 and w3392;
w7357 <= not w2468 and w3477;
w7358 <= not w2399 and w3541;
w7359 <= not w7357 and not w7358;
w7360 <= not w7356 and w7359;
w7361 <= w3303 and w6526;
w7362 <= w7360 and not w7361;
w7363 <= a(29) and not w7362;
w7364 <= not w7362 and not w7363;
w7365 <= a(29) and not w7363;
w7366 <= not w7364 and not w7365;
w7367 <= not w6748 and not w6751;
w7368 <= w6750 and not w6751;
w7369 <= not w7367 and not w7368;
w7370 <= not w7366 and not w7369;
w7371 <= not w7366 and not w7370;
w7372 <= not w7369 and not w7370;
w7373 <= not w7371 and not w7372;
w7374 <= not w2399 and w3392;
w7375 <= not w2506 and w3477;
w7376 <= not w2468 and w3541;
w7377 <= not w7375 and not w7376;
w7378 <= not w7374 and w7377;
w7379 <= w3303 and w6581;
w7380 <= w7378 and not w7379;
w7381 <= a(29) and not w7380;
w7382 <= not w7380 and not w7381;
w7383 <= a(29) and not w7381;
w7384 <= not w7382 and not w7383;
w7385 <= not w6726 and not w6738;
w7386 <= not w6737 and not w6738;
w7387 <= not w7385 and not w7386;
w7388 <= not w7384 and not w7387;
w7389 <= not w7384 and not w7388;
w7390 <= not w7387 and not w7388;
w7391 <= not w7389 and not w7390;
w7392 <= not w2468 and w3392;
w7393 <= not w2609 and w3477;
w7394 <= not w2506 and w3541;
w7395 <= not w7393 and not w7394;
w7396 <= not w7392 and w7395;
w7397 <= w3303 and w6630;
w7398 <= w7396 and not w7397;
w7399 <= a(29) and not w7398;
w7400 <= not w7398 and not w7399;
w7401 <= a(29) and not w7399;
w7402 <= not w7400 and not w7401;
w7403 <= w2671 and not w2764;
w7404 <= not w6730 and not w7403;
w7405 <= w10 and not w7404;
w7406 <= not w2764 and w2963;
w7407 <= not w2671 and w2955;
w7408 <= not w7406 and not w7407;
w7409 <= not w7405 and w7408;
w7410 <= not w7402 and not w7409;
w7411 <= not w7402 and not w7410;
w7412 <= not w7409 and not w7410;
w7413 <= not w7411 and not w7412;
w7414 <= not w10 and not w2955;
w7415 <= not w2764 and not w7414;
w7416 <= not w2764 and w3541;
w7417 <= not w2671 and w3392;
w7418 <= not w7416 and not w7417;
w7419 <= w3303 and not w7404;
w7420 <= w7418 and not w7419;
w7421 <= a(29) and not w7420;
w7422 <= a(29) and not w7421;
w7423 <= not w7420 and not w7421;
w7424 <= not w7422 and not w7423;
w7425 <= not w2764 and not w3302;
w7426 <= a(29) and not w7425;
w7427 <= not w7424 and w7426;
w7428 <= not w2609 and w3392;
w7429 <= not w2764 and w3477;
w7430 <= not w2671 and w3541;
w7431 <= not w7429 and not w7430;
w7432 <= not w7428 and w7431;
w7433 <= not w3303 and w7432;
w7434 <= not w6733 and w7432;
w7435 <= not w7433 and not w7434;
w7436 <= a(29) and not w7435;
w7437 <= not a(29) and w7435;
w7438 <= not w7436 and not w7437;
w7439 <= w7427 and not w7438;
w7440 <= w7415 and w7439;
w7441 <= not w2506 and w3392;
w7442 <= not w2671 and w3477;
w7443 <= not w2609 and w3541;
w7444 <= not w7442 and not w7443;
w7445 <= not w7441 and w7444;
w7446 <= w3303 and w6741;
w7447 <= w7445 and not w7446;
w7448 <= a(29) and not w7447;
w7449 <= not w7447 and not w7448;
w7450 <= a(29) and not w7448;
w7451 <= not w7449 and not w7450;
w7452 <= not w7415 and w7439;
w7453 <= w7415 and not w7439;
w7454 <= not w7452 and not w7453;
w7455 <= not w7451 and not w7454;
w7456 <= not w7440 and not w7455;
w7457 <= not w7413 and not w7456;
w7458 <= not w7410 and not w7457;
w7459 <= not w7391 and not w7458;
w7460 <= not w7388 and not w7459;
w7461 <= not w7373 and not w7460;
w7462 <= not w7370 and not w7461;
w7463 <= not w7355 and not w7462;
w7464 <= not w7352 and not w7463;
w7465 <= not w7337 and not w7464;
w7466 <= not w7334 and not w7465;
w7467 <= w7307 and w7318;
w7468 <= not w7319 and not w7467;
w7469 <= not w7466 and w7468;
w7470 <= not w7319 and not w7469;
w7471 <= w7292 and w7303;
w7472 <= not w7304 and not w7471;
w7473 <= not w7470 and w7472;
w7474 <= not w7304 and not w7473;
w7475 <= not w6775 and w6786;
w7476 <= not w6787 and not w7475;
w7477 <= not w7474 and w7476;
w7478 <= not w1714 and w3819;
w7479 <= not w1848 and w3902;
w7480 <= not w1812 and w3981;
w7481 <= not w7479 and not w7480;
w7482 <= not w7478 and w7481;
w7483 <= w3985 and w5786;
w7484 <= w7482 and not w7483;
w7485 <= a(26) and not w7484;
w7486 <= not w7484 and not w7485;
w7487 <= a(26) and not w7485;
w7488 <= not w7486 and not w7487;
w7489 <= w7474 and not w7476;
w7490 <= not w7477 and not w7489;
w7491 <= not w7488 and w7490;
w7492 <= not w7477 and not w7491;
w7493 <= not w7289 and not w7492;
w7494 <= w7289 and w7492;
w7495 <= not w7493 and not w7494;
w7496 <= not w1299 and w4629;
w7497 <= not w1507 and w4468;
w7498 <= not w1407 and w4539;
w7499 <= not w7497 and not w7498;
w7500 <= not w7496 and w7499;
w7501 <= w4471 and w5049;
w7502 <= w7500 and not w7501;
w7503 <= a(23) and not w7502;
w7504 <= a(23) and not w7503;
w7505 <= not w7502 and not w7503;
w7506 <= not w7504 and not w7505;
w7507 <= w7495 and not w7506;
w7508 <= not w7493 and not w7507;
w7509 <= not w7286 and not w7508;
w7510 <= w7286 and w7508;
w7511 <= not w7509 and not w7510;
w7512 <= not w893 and w5431;
w7513 <= not w1113 and w4870;
w7514 <= not w995 and w5342;
w7515 <= not w7513 and not w7514;
w7516 <= not w7512 and w7515;
w7517 <= w4568 and w4873;
w7518 <= w7516 and not w7517;
w7519 <= a(20) and not w7518;
w7520 <= a(20) and not w7519;
w7521 <= not w7518 and not w7519;
w7522 <= not w7520 and not w7521;
w7523 <= w7511 and not w7522;
w7524 <= not w7509 and not w7523;
w7525 <= not w7271 and w7282;
w7526 <= not w7283 and not w7525;
w7527 <= not w7524 and w7526;
w7528 <= not w7283 and not w7527;
w7529 <= not w7269 and not w7528;
w7530 <= w7269 and w7528;
w7531 <= not w7529 and not w7530;
w7532 <= not w2947 and w6168;
w7533 <= not w522 and w5598;
w7534 <= not w327 and w5874;
w7535 <= not w7533 and not w7534;
w7536 <= not w7532 and w7535;
w7537 <= w2953 and w5601;
w7538 <= w7536 and not w7537;
w7539 <= a(17) and not w7538;
w7540 <= a(17) and not w7539;
w7541 <= not w7538 and not w7539;
w7542 <= not w7540 and not w7541;
w7543 <= w7531 and not w7542;
w7544 <= not w7529 and not w7543;
w7545 <= not w7266 and not w7544;
w7546 <= w7266 and w7544;
w7547 <= not w7545 and not w7546;
w7548 <= not w3740 and w7036;
w7549 <= not w3540 and w6337;
w7550 <= not w3391 and w6886;
w7551 <= not w7549 and not w7550;
w7552 <= not w7548 and w7551;
w7553 <= w3753 and w6332;
w7554 <= w7552 and not w7553;
w7555 <= a(14) and not w7554;
w7556 <= a(14) and not w7555;
w7557 <= not w7554 and not w7555;
w7558 <= not w7556 and not w7557;
w7559 <= w7547 and not w7558;
w7560 <= not w7545 and not w7559;
w7561 <= w7251 and not w7263;
w7562 <= not w7262 and not w7263;
w7563 <= not w7561 and not w7562;
w7564 <= not w7560 and not w7563;
w7565 <= not w7263 and not w7564;
w7566 <= not w3812 and w7226;
w7567 <= not w7218 and w7224;
w7568 <= not w4450 and w7567;
w7569 <= not w7566 and not w7568;
w7570 <= not w7229 and w7569;
w7571 <= not w4544 and w7569;
w7572 <= not w7570 and not w7571;
w7573 <= a(11) and not w7572;
w7574 <= not a(11) and w7572;
w7575 <= not w7573 and not w7574;
w7576 <= not w7565 and not w7575;
w7577 <= w7202 and not w7214;
w7578 <= not w7213 and not w7214;
w7579 <= not w7577 and not w7578;
w7580 <= w7565 and w7575;
w7581 <= not w7576 and not w7580;
w7582 <= not w7579 and w7581;
w7583 <= not w7576 and not w7582;
w7584 <= not w7249 and not w7583;
w7585 <= w7249 and w7583;
w7586 <= not w7584 and not w7585;
w7587 <= w7547 and not w7559;
w7588 <= not w7558 and not w7559;
w7589 <= not w7587 and not w7588;
w7590 <= w7531 and not w7543;
w7591 <= not w7542 and not w7543;
w7592 <= not w7590 and not w7591;
w7593 <= not w327 and w6168;
w7594 <= not w645 and w5598;
w7595 <= not w522 and w5874;
w7596 <= not w7594 and not w7595;
w7597 <= not w7593 and w7596;
w7598 <= w3282 and w5601;
w7599 <= w7597 and not w7598;
w7600 <= a(17) and not w7599;
w7601 <= not w7599 and not w7600;
w7602 <= a(17) and not w7600;
w7603 <= not w7601 and not w7602;
w7604 <= w7524 and not w7526;
w7605 <= not w7527 and not w7604;
w7606 <= not w7603 and w7605;
w7607 <= not w7603 and not w7606;
w7608 <= w7605 and not w7606;
w7609 <= not w7607 and not w7608;
w7610 <= w7511 and not w7523;
w7611 <= not w7522 and not w7523;
w7612 <= not w7610 and not w7611;
w7613 <= w7495 and not w7507;
w7614 <= not w7506 and not w7507;
w7615 <= not w7613 and not w7614;
w7616 <= w7470 and not w7472;
w7617 <= not w7473 and not w7616;
w7618 <= not w1812 and w3819;
w7619 <= not w1927 and w3902;
w7620 <= not w1848 and w3981;
w7621 <= not w7619 and not w7620;
w7622 <= not w7618 and w7621;
w7623 <= not w3985 and w7622;
w7624 <= not w5942 and w7622;
w7625 <= not w7623 and not w7624;
w7626 <= a(26) and not w7625;
w7627 <= not a(26) and w7625;
w7628 <= not w7626 and not w7627;
w7629 <= w7617 and not w7628;
w7630 <= w7466 and not w7468;
w7631 <= not w7469 and not w7630;
w7632 <= not w1848 and w3819;
w7633 <= not w1992 and w3902;
w7634 <= not w1927 and w3981;
w7635 <= not w7633 and not w7634;
w7636 <= not w7632 and w7635;
w7637 <= not w3985 and w7636;
w7638 <= not w5769 and w7636;
w7639 <= not w7637 and not w7638;
w7640 <= a(26) and not w7639;
w7641 <= not a(26) and w7639;
w7642 <= not w7640 and not w7641;
w7643 <= w7631 and not w7642;
w7644 <= w7337 and w7464;
w7645 <= not w7465 and not w7644;
w7646 <= not w1927 and w3819;
w7647 <= not w2087 and w3902;
w7648 <= not w1992 and w3981;
w7649 <= not w7647 and not w7648;
w7650 <= not w7646 and w7649;
w7651 <= not w3985 and w7650;
w7652 <= not w6078 and w7650;
w7653 <= not w7651 and not w7652;
w7654 <= a(26) and not w7653;
w7655 <= not a(26) and w7653;
w7656 <= not w7654 and not w7655;
w7657 <= w7645 and not w7656;
w7658 <= w7355 and w7462;
w7659 <= not w7463 and not w7658;
w7660 <= not w1992 and w3819;
w7661 <= not w2124 and w3902;
w7662 <= not w2087 and w3981;
w7663 <= not w7661 and not w7662;
w7664 <= not w7660 and w7663;
w7665 <= not w3985 and w7664;
w7666 <= not w6414 and w7664;
w7667 <= not w7665 and not w7666;
w7668 <= a(26) and not w7667;
w7669 <= not a(26) and w7667;
w7670 <= not w7668 and not w7669;
w7671 <= w7659 and not w7670;
w7672 <= w7373 and w7460;
w7673 <= not w7461 and not w7672;
w7674 <= not w2087 and w3819;
w7675 <= not w2226 and w3902;
w7676 <= not w2124 and w3981;
w7677 <= not w7675 and not w7676;
w7678 <= not w7674 and w7677;
w7679 <= not w3985 and w7678;
w7680 <= not w6427 and w7678;
w7681 <= not w7679 and not w7680;
w7682 <= a(26) and not w7681;
w7683 <= not a(26) and w7681;
w7684 <= not w7682 and not w7683;
w7685 <= w7673 and not w7684;
w7686 <= w7391 and w7458;
w7687 <= not w7459 and not w7686;
w7688 <= not w2124 and w3819;
w7689 <= not w2323 and w3902;
w7690 <= not w2226 and w3981;
w7691 <= not w7689 and not w7690;
w7692 <= not w7688 and w7691;
w7693 <= not w3985 and w7692;
w7694 <= not w6057 and w7692;
w7695 <= not w7693 and not w7694;
w7696 <= a(26) and not w7695;
w7697 <= not a(26) and w7695;
w7698 <= not w7696 and not w7697;
w7699 <= w7687 and not w7698;
w7700 <= not w7413 and not w7457;
w7701 <= not w7456 and not w7457;
w7702 <= not w7700 and not w7701;
w7703 <= not w2226 and w3819;
w7704 <= not w2399 and w3902;
w7705 <= not w2323 and w3981;
w7706 <= not w7704 and not w7705;
w7707 <= not w7703 and w7706;
w7708 <= not w3985 and w7707;
w7709 <= not w6476 and w7707;
w7710 <= not w7708 and not w7709;
w7711 <= a(26) and not w7710;
w7712 <= not a(26) and w7710;
w7713 <= not w7711 and not w7712;
w7714 <= not w7702 and not w7713;
w7715 <= not w2323 and w3819;
w7716 <= not w2468 and w3902;
w7717 <= not w2399 and w3981;
w7718 <= not w7716 and not w7717;
w7719 <= not w7715 and w7718;
w7720 <= w3985 and w6526;
w7721 <= w7719 and not w7720;
w7722 <= a(26) and not w7721;
w7723 <= not w7721 and not w7722;
w7724 <= a(26) and not w7722;
w7725 <= not w7723 and not w7724;
w7726 <= w7451 and w7454;
w7727 <= not w7455 and not w7726;
w7728 <= not w7725 and w7727;
w7729 <= not w7725 and not w7728;
w7730 <= w7727 and not w7728;
w7731 <= not w7729 and not w7730;
w7732 <= not w2399 and w3819;
w7733 <= not w2506 and w3902;
w7734 <= not w2468 and w3981;
w7735 <= not w7733 and not w7734;
w7736 <= not w7732 and w7735;
w7737 <= w3985 and w6581;
w7738 <= w7736 and not w7737;
w7739 <= a(26) and not w7738;
w7740 <= not w7738 and not w7739;
w7741 <= a(26) and not w7739;
w7742 <= not w7740 and not w7741;
w7743 <= not w7427 and w7438;
w7744 <= not w7439 and not w7743;
w7745 <= not w7742 and w7744;
w7746 <= not w7742 and not w7745;
w7747 <= w7744 and not w7745;
w7748 <= not w7746 and not w7747;
w7749 <= w7424 and not w7426;
w7750 <= not w7427 and not w7749;
w7751 <= not w2468 and w3819;
w7752 <= not w2609 and w3902;
w7753 <= not w2506 and w3981;
w7754 <= not w7752 and not w7753;
w7755 <= not w7751 and w7754;
w7756 <= not w3985 and w7755;
w7757 <= not w6630 and w7755;
w7758 <= not w7756 and not w7757;
w7759 <= a(26) and not w7758;
w7760 <= not a(26) and w7758;
w7761 <= not w7759 and not w7760;
w7762 <= w7750 and not w7761;
w7763 <= not w2764 and w3981;
w7764 <= not w2671 and w3819;
w7765 <= not w7763 and not w7764;
w7766 <= w3985 and not w7404;
w7767 <= w7765 and not w7766;
w7768 <= a(26) and not w7767;
w7769 <= a(26) and not w7768;
w7770 <= not w7767 and not w7768;
w7771 <= not w7769 and not w7770;
w7772 <= not w2764 and not w3815;
w7773 <= a(26) and not w7772;
w7774 <= not w7771 and w7773;
w7775 <= not w2609 and w3819;
w7776 <= not w2764 and w3902;
w7777 <= not w2671 and w3981;
w7778 <= not w7776 and not w7777;
w7779 <= not w7775 and w7778;
w7780 <= not w3985 and w7779;
w7781 <= not w6733 and w7779;
w7782 <= not w7780 and not w7781;
w7783 <= a(26) and not w7782;
w7784 <= not a(26) and w7782;
w7785 <= not w7783 and not w7784;
w7786 <= w7774 and not w7785;
w7787 <= w7425 and w7786;
w7788 <= w7786 and not w7787;
w7789 <= w7425 and not w7787;
w7790 <= not w7788 and not w7789;
w7791 <= not w2506 and w3819;
w7792 <= not w2671 and w3902;
w7793 <= not w2609 and w3981;
w7794 <= not w7792 and not w7793;
w7795 <= not w7791 and w7794;
w7796 <= w3985 and w6741;
w7797 <= w7795 and not w7796;
w7798 <= a(26) and not w7797;
w7799 <= a(26) and not w7798;
w7800 <= not w7797 and not w7798;
w7801 <= not w7799 and not w7800;
w7802 <= not w7790 and not w7801;
w7803 <= not w7787 and not w7802;
w7804 <= not w7750 and w7761;
w7805 <= not w7762 and not w7804;
w7806 <= not w7803 and w7805;
w7807 <= not w7762 and not w7806;
w7808 <= not w7748 and not w7807;
w7809 <= not w7745 and not w7808;
w7810 <= not w7731 and not w7809;
w7811 <= not w7728 and not w7810;
w7812 <= not w7702 and not w7714;
w7813 <= not w7713 and not w7714;
w7814 <= not w7812 and not w7813;
w7815 <= not w7811 and not w7814;
w7816 <= not w7714 and not w7815;
w7817 <= w7687 and not w7699;
w7818 <= not w7698 and not w7699;
w7819 <= not w7817 and not w7818;
w7820 <= not w7816 and not w7819;
w7821 <= not w7699 and not w7820;
w7822 <= w7673 and not w7685;
w7823 <= not w7684 and not w7685;
w7824 <= not w7822 and not w7823;
w7825 <= not w7821 and not w7824;
w7826 <= not w7685 and not w7825;
w7827 <= w7659 and not w7671;
w7828 <= not w7670 and not w7671;
w7829 <= not w7827 and not w7828;
w7830 <= not w7826 and not w7829;
w7831 <= not w7671 and not w7830;
w7832 <= w7645 and not w7657;
w7833 <= not w7656 and not w7657;
w7834 <= not w7832 and not w7833;
w7835 <= not w7831 and not w7834;
w7836 <= not w7657 and not w7835;
w7837 <= w7631 and not w7643;
w7838 <= not w7642 and not w7643;
w7839 <= not w7837 and not w7838;
w7840 <= not w7836 and not w7839;
w7841 <= not w7643 and not w7840;
w7842 <= w7617 and not w7629;
w7843 <= not w7628 and not w7629;
w7844 <= not w7842 and not w7843;
w7845 <= not w7841 and not w7844;
w7846 <= not w7629 and not w7845;
w7847 <= w7488 and not w7490;
w7848 <= not w7491 and not w7847;
w7849 <= not w7846 and w7848;
w7850 <= not w1407 and w4629;
w7851 <= not w1600 and w4468;
w7852 <= not w1507 and w4539;
w7853 <= not w7851 and not w7852;
w7854 <= not w7850 and w7853;
w7855 <= w4471 and w5074;
w7856 <= w7854 and not w7855;
w7857 <= a(23) and not w7856;
w7858 <= not w7856 and not w7857;
w7859 <= a(23) and not w7857;
w7860 <= not w7858 and not w7859;
w7861 <= w7846 and not w7848;
w7862 <= not w7849 and not w7861;
w7863 <= not w7860 and w7862;
w7864 <= not w7849 and not w7863;
w7865 <= not w7615 and not w7864;
w7866 <= w7615 and w7864;
w7867 <= not w7865 and not w7866;
w7868 <= not w995 and w5431;
w7869 <= not w1170 and w4870;
w7870 <= not w1113 and w5342;
w7871 <= not w7869 and not w7870;
w7872 <= not w7868 and w7871;
w7873 <= w4364 and w4873;
w7874 <= w7872 and not w7873;
w7875 <= a(20) and not w7874;
w7876 <= a(20) and not w7875;
w7877 <= not w7874 and not w7875;
w7878 <= not w7876 and not w7877;
w7879 <= w7867 and not w7878;
w7880 <= not w7865 and not w7879;
w7881 <= not w7612 and not w7880;
w7882 <= w7612 and w7880;
w7883 <= not w7881 and not w7882;
w7884 <= not w522 and w6168;
w7885 <= not w802 and w5598;
w7886 <= not w645 and w5874;
w7887 <= not w7885 and not w7886;
w7888 <= not w7884 and w7887;
w7889 <= w3266 and w5601;
w7890 <= w7888 and not w7889;
w7891 <= a(17) and not w7890;
w7892 <= a(17) and not w7891;
w7893 <= not w7890 and not w7891;
w7894 <= not w7892 and not w7893;
w7895 <= w7883 and not w7894;
w7896 <= not w7881 and not w7895;
w7897 <= not w7609 and not w7896;
w7898 <= not w7606 and not w7897;
w7899 <= not w7592 and not w7898;
w7900 <= w7592 and w7898;
w7901 <= not w7899 and not w7900;
w7902 <= not w3391 and w7036;
w7903 <= not w3474 and w6337;
w7904 <= not w3540 and w6886;
w7905 <= not w7903 and not w7904;
w7906 <= not w7902 and w7905;
w7907 <= w3562 and w6332;
w7908 <= w7906 and not w7907;
w7909 <= a(14) and not w7908;
w7910 <= a(14) and not w7909;
w7911 <= not w7908 and not w7909;
w7912 <= not w7910 and not w7911;
w7913 <= w7901 and not w7912;
w7914 <= not w7899 and not w7913;
w7915 <= not w7589 and not w7914;
w7916 <= w7589 and w7914;
w7917 <= not w7915 and not w7916;
w7918 <= w7221 and not w7224;
w7919 <= not w3812 and w7918;
w7920 <= not w3899 and w7226;
w7921 <= not w3980 and w7567;
w7922 <= not w7920 and not w7921;
w7923 <= not w7919 and w7922;
w7924 <= w4002 and w7229;
w7925 <= w7923 and not w7924;
w7926 <= a(11) and not w7925;
w7927 <= a(11) and not w7926;
w7928 <= not w7925 and not w7926;
w7929 <= not w7927 and not w7928;
w7930 <= w7917 and not w7929;
w7931 <= not w7915 and not w7930;
w7932 <= not w4450 and w7918;
w7933 <= not w3980 and w7226;
w7934 <= not w3812 and w7567;
w7935 <= not w7933 and not w7934;
w7936 <= not w7932 and w7935;
w7937 <= not w7229 and w7936;
w7938 <= not w4650 and w7936;
w7939 <= not w7937 and not w7938;
w7940 <= a(11) and not w7939;
w7941 <= not a(11) and w7939;
w7942 <= not w7940 and not w7941;
w7943 <= not w7931 and not w7942;
w7944 <= w7931 and w7942;
w7945 <= not w7943 and not w7944;
w7946 <= not w7560 and not w7564;
w7947 <= not w7563 and not w7564;
w7948 <= not w7946 and not w7947;
w7949 <= w7945 and not w7948;
w7950 <= not w7943 and not w7949;
w7951 <= w7579 and not w7581;
w7952 <= not w7582 and not w7951;
w7953 <= not w7950 and w7952;
w7954 <= w7945 and not w7949;
w7955 <= not w7948 and not w7949;
w7956 <= not w7954 and not w7955;
w7957 <= w7901 and not w7913;
w7958 <= not w7912 and not w7913;
w7959 <= not w7957 and not w7958;
w7960 <= w7609 and w7896;
w7961 <= not w7897 and not w7960;
w7962 <= not w3540 and w7036;
w7963 <= not w2947 and w6337;
w7964 <= not w3474 and w6886;
w7965 <= not w7963 and not w7964;
w7966 <= not w7962 and w7965;
w7967 <= not w6332 and w7966;
w7968 <= not w4019 and w7966;
w7969 <= not w7967 and not w7968;
w7970 <= a(14) and not w7969;
w7971 <= not a(14) and w7969;
w7972 <= not w7970 and not w7971;
w7973 <= w7961 and not w7972;
w7974 <= w7883 and not w7895;
w7975 <= not w7894 and not w7895;
w7976 <= not w7974 and not w7975;
w7977 <= w7867 and not w7879;
w7978 <= not w7878 and not w7879;
w7979 <= not w7977 and not w7978;
w7980 <= not w1507 and w4629;
w7981 <= not w1714 and w4468;
w7982 <= not w1600 and w4539;
w7983 <= not w7981 and not w7982;
w7984 <= not w7980 and w7983;
w7985 <= w4471 and w5496;
w7986 <= w7984 and not w7985;
w7987 <= a(23) and not w7986;
w7988 <= not w7986 and not w7987;
w7989 <= a(23) and not w7987;
w7990 <= not w7988 and not w7989;
w7991 <= not w7841 and not w7845;
w7992 <= not w7844 and not w7845;
w7993 <= not w7991 and not w7992;
w7994 <= not w7990 and not w7993;
w7995 <= not w7990 and not w7994;
w7996 <= not w7993 and not w7994;
w7997 <= not w7995 and not w7996;
w7998 <= not w1600 and w4629;
w7999 <= not w1812 and w4468;
w8000 <= not w1714 and w4539;
w8001 <= not w7999 and not w8000;
w8002 <= not w7998 and w8001;
w8003 <= w4471 and w5263;
w8004 <= w8002 and not w8003;
w8005 <= a(23) and not w8004;
w8006 <= not w8004 and not w8005;
w8007 <= a(23) and not w8005;
w8008 <= not w8006 and not w8007;
w8009 <= not w7836 and not w7840;
w8010 <= not w7839 and not w7840;
w8011 <= not w8009 and not w8010;
w8012 <= not w8008 and not w8011;
w8013 <= not w8008 and not w8012;
w8014 <= not w8011 and not w8012;
w8015 <= not w8013 and not w8014;
w8016 <= not w1714 and w4629;
w8017 <= not w1848 and w4468;
w8018 <= not w1812 and w4539;
w8019 <= not w8017 and not w8018;
w8020 <= not w8016 and w8019;
w8021 <= w4471 and w5786;
w8022 <= w8020 and not w8021;
w8023 <= a(23) and not w8022;
w8024 <= not w8022 and not w8023;
w8025 <= a(23) and not w8023;
w8026 <= not w8024 and not w8025;
w8027 <= not w7831 and not w7835;
w8028 <= not w7834 and not w7835;
w8029 <= not w8027 and not w8028;
w8030 <= not w8026 and not w8029;
w8031 <= not w8026 and not w8030;
w8032 <= not w8029 and not w8030;
w8033 <= not w8031 and not w8032;
w8034 <= not w1812 and w4629;
w8035 <= not w1927 and w4468;
w8036 <= not w1848 and w4539;
w8037 <= not w8035 and not w8036;
w8038 <= not w8034 and w8037;
w8039 <= w4471 and w5942;
w8040 <= w8038 and not w8039;
w8041 <= a(23) and not w8040;
w8042 <= not w8040 and not w8041;
w8043 <= a(23) and not w8041;
w8044 <= not w8042 and not w8043;
w8045 <= not w7826 and not w7830;
w8046 <= not w7829 and not w7830;
w8047 <= not w8045 and not w8046;
w8048 <= not w8044 and not w8047;
w8049 <= not w8044 and not w8048;
w8050 <= not w8047 and not w8048;
w8051 <= not w8049 and not w8050;
w8052 <= not w1848 and w4629;
w8053 <= not w1992 and w4468;
w8054 <= not w1927 and w4539;
w8055 <= not w8053 and not w8054;
w8056 <= not w8052 and w8055;
w8057 <= w4471 and w5769;
w8058 <= w8056 and not w8057;
w8059 <= a(23) and not w8058;
w8060 <= not w8058 and not w8059;
w8061 <= a(23) and not w8059;
w8062 <= not w8060 and not w8061;
w8063 <= not w7821 and not w7825;
w8064 <= not w7824 and not w7825;
w8065 <= not w8063 and not w8064;
w8066 <= not w8062 and not w8065;
w8067 <= not w8062 and not w8066;
w8068 <= not w8065 and not w8066;
w8069 <= not w8067 and not w8068;
w8070 <= not w1927 and w4629;
w8071 <= not w2087 and w4468;
w8072 <= not w1992 and w4539;
w8073 <= not w8071 and not w8072;
w8074 <= not w8070 and w8073;
w8075 <= w4471 and w6078;
w8076 <= w8074 and not w8075;
w8077 <= a(23) and not w8076;
w8078 <= not w8076 and not w8077;
w8079 <= a(23) and not w8077;
w8080 <= not w8078 and not w8079;
w8081 <= not w7816 and not w7820;
w8082 <= not w7819 and not w7820;
w8083 <= not w8081 and not w8082;
w8084 <= not w8080 and not w8083;
w8085 <= not w8080 and not w8084;
w8086 <= not w8083 and not w8084;
w8087 <= not w8085 and not w8086;
w8088 <= not w1992 and w4629;
w8089 <= not w2124 and w4468;
w8090 <= not w2087 and w4539;
w8091 <= not w8089 and not w8090;
w8092 <= not w8088 and w8091;
w8093 <= w4471 and w6414;
w8094 <= w8092 and not w8093;
w8095 <= a(23) and not w8094;
w8096 <= not w8094 and not w8095;
w8097 <= a(23) and not w8095;
w8098 <= not w8096 and not w8097;
w8099 <= not w7811 and not w7815;
w8100 <= not w7814 and not w7815;
w8101 <= not w8099 and not w8100;
w8102 <= not w8098 and not w8101;
w8103 <= not w8098 and not w8102;
w8104 <= not w8101 and not w8102;
w8105 <= not w8103 and not w8104;
w8106 <= w7731 and w7809;
w8107 <= not w7810 and not w8106;
w8108 <= not w2087 and w4629;
w8109 <= not w2226 and w4468;
w8110 <= not w2124 and w4539;
w8111 <= not w8109 and not w8110;
w8112 <= not w8108 and w8111;
w8113 <= not w4471 and w8112;
w8114 <= not w6427 and w8112;
w8115 <= not w8113 and not w8114;
w8116 <= a(23) and not w8115;
w8117 <= not a(23) and w8115;
w8118 <= not w8116 and not w8117;
w8119 <= w8107 and not w8118;
w8120 <= w7748 and w7807;
w8121 <= not w7808 and not w8120;
w8122 <= not w2124 and w4629;
w8123 <= not w2323 and w4468;
w8124 <= not w2226 and w4539;
w8125 <= not w8123 and not w8124;
w8126 <= not w8122 and w8125;
w8127 <= not w4471 and w8126;
w8128 <= not w6057 and w8126;
w8129 <= not w8127 and not w8128;
w8130 <= a(23) and not w8129;
w8131 <= not a(23) and w8129;
w8132 <= not w8130 and not w8131;
w8133 <= w8121 and not w8132;
w8134 <= not w2226 and w4629;
w8135 <= not w2399 and w4468;
w8136 <= not w2323 and w4539;
w8137 <= not w8135 and not w8136;
w8138 <= not w8134 and w8137;
w8139 <= w4471 and w6476;
w8140 <= w8138 and not w8139;
w8141 <= a(23) and not w8140;
w8142 <= not w8140 and not w8141;
w8143 <= a(23) and not w8141;
w8144 <= not w8142 and not w8143;
w8145 <= w7803 and not w7805;
w8146 <= not w7806 and not w8145;
w8147 <= not w8144 and w8146;
w8148 <= not w8144 and not w8147;
w8149 <= w8146 and not w8147;
w8150 <= not w8148 and not w8149;
w8151 <= not w7790 and not w7802;
w8152 <= not w7801 and not w7802;
w8153 <= not w8151 and not w8152;
w8154 <= not w2323 and w4629;
w8155 <= not w2468 and w4468;
w8156 <= not w2399 and w4539;
w8157 <= not w8155 and not w8156;
w8158 <= not w8154 and w8157;
w8159 <= not w4471 and w8158;
w8160 <= not w6526 and w8158;
w8161 <= not w8159 and not w8160;
w8162 <= a(23) and not w8161;
w8163 <= not a(23) and w8161;
w8164 <= not w8162 and not w8163;
w8165 <= not w8153 and not w8164;
w8166 <= not w2399 and w4629;
w8167 <= not w2506 and w4468;
w8168 <= not w2468 and w4539;
w8169 <= not w8167 and not w8168;
w8170 <= not w8166 and w8169;
w8171 <= w4471 and w6581;
w8172 <= w8170 and not w8171;
w8173 <= a(23) and not w8172;
w8174 <= not w8172 and not w8173;
w8175 <= a(23) and not w8173;
w8176 <= not w8174 and not w8175;
w8177 <= not w7774 and w7785;
w8178 <= not w7786 and not w8177;
w8179 <= not w8176 and w8178;
w8180 <= not w8176 and not w8179;
w8181 <= w8178 and not w8179;
w8182 <= not w8180 and not w8181;
w8183 <= w7771 and not w7773;
w8184 <= not w7774 and not w8183;
w8185 <= not w2468 and w4629;
w8186 <= not w2609 and w4468;
w8187 <= not w2506 and w4539;
w8188 <= not w8186 and not w8187;
w8189 <= not w8185 and w8188;
w8190 <= not w4471 and w8189;
w8191 <= not w6630 and w8189;
w8192 <= not w8190 and not w8191;
w8193 <= a(23) and not w8192;
w8194 <= not a(23) and w8192;
w8195 <= not w8193 and not w8194;
w8196 <= w8184 and not w8195;
w8197 <= not w2764 and w4539;
w8198 <= not w2671 and w4629;
w8199 <= not w8197 and not w8198;
w8200 <= w4471 and not w7404;
w8201 <= w8199 and not w8200;
w8202 <= a(23) and not w8201;
w8203 <= a(23) and not w8202;
w8204 <= not w8201 and not w8202;
w8205 <= not w8203 and not w8204;
w8206 <= not w2764 and not w4463;
w8207 <= a(23) and not w8206;
w8208 <= not w8205 and w8207;
w8209 <= not w2609 and w4629;
w8210 <= not w2764 and w4468;
w8211 <= not w2671 and w4539;
w8212 <= not w8210 and not w8211;
w8213 <= not w8209 and w8212;
w8214 <= not w4471 and w8213;
w8215 <= not w6733 and w8213;
w8216 <= not w8214 and not w8215;
w8217 <= a(23) and not w8216;
w8218 <= not a(23) and w8216;
w8219 <= not w8217 and not w8218;
w8220 <= w8208 and not w8219;
w8221 <= w7772 and w8220;
w8222 <= w8220 and not w8221;
w8223 <= w7772 and not w8221;
w8224 <= not w8222 and not w8223;
w8225 <= not w2506 and w4629;
w8226 <= not w2671 and w4468;
w8227 <= not w2609 and w4539;
w8228 <= not w8226 and not w8227;
w8229 <= not w8225 and w8228;
w8230 <= w4471 and w6741;
w8231 <= w8229 and not w8230;
w8232 <= a(23) and not w8231;
w8233 <= a(23) and not w8232;
w8234 <= not w8231 and not w8232;
w8235 <= not w8233 and not w8234;
w8236 <= not w8224 and not w8235;
w8237 <= not w8221 and not w8236;
w8238 <= not w8184 and w8195;
w8239 <= not w8196 and not w8238;
w8240 <= not w8237 and w8239;
w8241 <= not w8196 and not w8240;
w8242 <= not w8182 and not w8241;
w8243 <= not w8179 and not w8242;
w8244 <= w8153 and w8164;
w8245 <= not w8165 and not w8244;
w8246 <= not w8243 and w8245;
w8247 <= not w8165 and not w8246;
w8248 <= not w8150 and not w8247;
w8249 <= not w8147 and not w8248;
w8250 <= w8121 and not w8133;
w8251 <= not w8132 and not w8133;
w8252 <= not w8250 and not w8251;
w8253 <= not w8249 and not w8252;
w8254 <= not w8133 and not w8253;
w8255 <= not w8107 and w8118;
w8256 <= not w8119 and not w8255;
w8257 <= not w8254 and w8256;
w8258 <= not w8119 and not w8257;
w8259 <= not w8105 and not w8258;
w8260 <= not w8102 and not w8259;
w8261 <= not w8087 and not w8260;
w8262 <= not w8084 and not w8261;
w8263 <= not w8069 and not w8262;
w8264 <= not w8066 and not w8263;
w8265 <= not w8051 and not w8264;
w8266 <= not w8048 and not w8265;
w8267 <= not w8033 and not w8266;
w8268 <= not w8030 and not w8267;
w8269 <= not w8015 and not w8268;
w8270 <= not w8012 and not w8269;
w8271 <= not w7997 and not w8270;
w8272 <= not w7994 and not w8271;
w8273 <= w7860 and not w7862;
w8274 <= not w7863 and not w8273;
w8275 <= not w8272 and w8274;
w8276 <= not w1113 and w5431;
w8277 <= not w1299 and w4870;
w8278 <= not w1170 and w5342;
w8279 <= not w8277 and not w8278;
w8280 <= not w8276 and w8279;
w8281 <= w4796 and w4873;
w8282 <= w8280 and not w8281;
w8283 <= a(20) and not w8282;
w8284 <= not w8282 and not w8283;
w8285 <= a(20) and not w8283;
w8286 <= not w8284 and not w8285;
w8287 <= w8272 and not w8274;
w8288 <= not w8275 and not w8287;
w8289 <= not w8286 and w8288;
w8290 <= not w8275 and not w8289;
w8291 <= not w7979 and not w8290;
w8292 <= w7979 and w8290;
w8293 <= not w8291 and not w8292;
w8294 <= not w645 and w6168;
w8295 <= not w893 and w5598;
w8296 <= not w802 and w5874;
w8297 <= not w8295 and not w8296;
w8298 <= not w8294 and w8297;
w8299 <= w4114 and w5601;
w8300 <= w8298 and not w8299;
w8301 <= a(17) and not w8300;
w8302 <= a(17) and not w8301;
w8303 <= not w8300 and not w8301;
w8304 <= not w8302 and not w8303;
w8305 <= w8293 and not w8304;
w8306 <= not w8291 and not w8305;
w8307 <= not w7976 and not w8306;
w8308 <= w7976 and w8306;
w8309 <= not w8307 and not w8308;
w8310 <= not w3474 and w7036;
w8311 <= not w327 and w6337;
w8312 <= not w2947 and w6886;
w8313 <= not w8311 and not w8312;
w8314 <= not w8310 and w8313;
w8315 <= w3650 and w6332;
w8316 <= w8314 and not w8315;
w8317 <= a(14) and not w8316;
w8318 <= a(14) and not w8317;
w8319 <= not w8316 and not w8317;
w8320 <= not w8318 and not w8319;
w8321 <= w8309 and not w8320;
w8322 <= not w8307 and not w8321;
w8323 <= not w7961 and w7972;
w8324 <= not w7973 and not w8323;
w8325 <= not w8322 and w8324;
w8326 <= not w7973 and not w8325;
w8327 <= not w7959 and not w8326;
w8328 <= w7959 and w8326;
w8329 <= not w8327 and not w8328;
w8330 <= not w3980 and w7918;
w8331 <= not w3740 and w7226;
w8332 <= not w3899 and w7567;
w8333 <= not w8331 and not w8332;
w8334 <= not w8330 and w8333;
w8335 <= w4412 and w7229;
w8336 <= w8334 and not w8335;
w8337 <= a(11) and not w8336;
w8338 <= a(11) and not w8337;
w8339 <= not w8336 and not w8337;
w8340 <= not w8338 and not w8339;
w8341 <= w8329 and not w8340;
w8342 <= not w8327 and not w8341;
w8343 <= not a(6) and a(7);
w8344 <= a(6) and not a(7);
w8345 <= not w8343 and not w8344;
w8346 <= a(7) and not a(8);
w8347 <= not a(7) and a(8);
w8348 <= not w8346 and not w8347;
w8349 <= a(5) and not a(6);
w8350 <= not a(5) and a(6);
w8351 <= not w8349 and not w8350;
w8352 <= not w8348 and w8351;
w8353 <= w8345 and w8352;
w8354 <= not w4450 and w8353;
w8355 <= not w4457 and not w8354;
w8356 <= not w8348 and not w8351;
w8357 <= not w8354 and not w8356;
w8358 <= not w8355 and not w8357;
w8359 <= a(8) and not w8358;
w8360 <= not a(8) and w8358;
w8361 <= not w8359 and not w8360;
w8362 <= not w8342 and not w8361;
w8363 <= w7917 and not w7930;
w8364 <= not w7929 and not w7930;
w8365 <= not w8363 and not w8364;
w8366 <= w8342 and w8361;
w8367 <= not w8362 and not w8366;
w8368 <= not w8365 and w8367;
w8369 <= not w8362 and not w8368;
w8370 <= not w7956 and not w8369;
w8371 <= w7956 and w8369;
w8372 <= not w8370 and not w8371;
w8373 <= not w8365 and not w8368;
w8374 <= w8367 and not w8368;
w8375 <= not w8373 and not w8374;
w8376 <= w8309 and not w8321;
w8377 <= not w8320 and not w8321;
w8378 <= not w8376 and not w8377;
w8379 <= w8293 and not w8305;
w8380 <= not w8304 and not w8305;
w8381 <= not w8379 and not w8380;
w8382 <= w7997 and w8270;
w8383 <= not w8271 and not w8382;
w8384 <= not w1170 and w5431;
w8385 <= not w1407 and w4870;
w8386 <= not w1299 and w5342;
w8387 <= not w8385 and not w8386;
w8388 <= not w8384 and w8387;
w8389 <= not w4873 and w8388;
w8390 <= not w4783 and w8388;
w8391 <= not w8389 and not w8390;
w8392 <= a(20) and not w8391;
w8393 <= not a(20) and w8391;
w8394 <= not w8392 and not w8393;
w8395 <= w8383 and not w8394;
w8396 <= w8015 and w8268;
w8397 <= not w8269 and not w8396;
w8398 <= not w1299 and w5431;
w8399 <= not w1507 and w4870;
w8400 <= not w1407 and w5342;
w8401 <= not w8399 and not w8400;
w8402 <= not w8398 and w8401;
w8403 <= not w4873 and w8402;
w8404 <= not w5049 and w8402;
w8405 <= not w8403 and not w8404;
w8406 <= a(20) and not w8405;
w8407 <= not a(20) and w8405;
w8408 <= not w8406 and not w8407;
w8409 <= w8397 and not w8408;
w8410 <= w8033 and w8266;
w8411 <= not w8267 and not w8410;
w8412 <= not w1407 and w5431;
w8413 <= not w1600 and w4870;
w8414 <= not w1507 and w5342;
w8415 <= not w8413 and not w8414;
w8416 <= not w8412 and w8415;
w8417 <= not w4873 and w8416;
w8418 <= not w5074 and w8416;
w8419 <= not w8417 and not w8418;
w8420 <= a(20) and not w8419;
w8421 <= not a(20) and w8419;
w8422 <= not w8420 and not w8421;
w8423 <= w8411 and not w8422;
w8424 <= w8051 and w8264;
w8425 <= not w8265 and not w8424;
w8426 <= not w1507 and w5431;
w8427 <= not w1714 and w4870;
w8428 <= not w1600 and w5342;
w8429 <= not w8427 and not w8428;
w8430 <= not w8426 and w8429;
w8431 <= not w4873 and w8430;
w8432 <= not w5496 and w8430;
w8433 <= not w8431 and not w8432;
w8434 <= a(20) and not w8433;
w8435 <= not a(20) and w8433;
w8436 <= not w8434 and not w8435;
w8437 <= w8425 and not w8436;
w8438 <= w8069 and w8262;
w8439 <= not w8263 and not w8438;
w8440 <= not w1600 and w5431;
w8441 <= not w1812 and w4870;
w8442 <= not w1714 and w5342;
w8443 <= not w8441 and not w8442;
w8444 <= not w8440 and w8443;
w8445 <= not w4873 and w8444;
w8446 <= not w5263 and w8444;
w8447 <= not w8445 and not w8446;
w8448 <= a(20) and not w8447;
w8449 <= not a(20) and w8447;
w8450 <= not w8448 and not w8449;
w8451 <= w8439 and not w8450;
w8452 <= w8087 and w8260;
w8453 <= not w8261 and not w8452;
w8454 <= not w1714 and w5431;
w8455 <= not w1848 and w4870;
w8456 <= not w1812 and w5342;
w8457 <= not w8455 and not w8456;
w8458 <= not w8454 and w8457;
w8459 <= not w4873 and w8458;
w8460 <= not w5786 and w8458;
w8461 <= not w8459 and not w8460;
w8462 <= a(20) and not w8461;
w8463 <= not a(20) and w8461;
w8464 <= not w8462 and not w8463;
w8465 <= w8453 and not w8464;
w8466 <= w8105 and w8258;
w8467 <= not w8259 and not w8466;
w8468 <= not w1812 and w5431;
w8469 <= not w1927 and w4870;
w8470 <= not w1848 and w5342;
w8471 <= not w8469 and not w8470;
w8472 <= not w8468 and w8471;
w8473 <= not w4873 and w8472;
w8474 <= not w5942 and w8472;
w8475 <= not w8473 and not w8474;
w8476 <= a(20) and not w8475;
w8477 <= not a(20) and w8475;
w8478 <= not w8476 and not w8477;
w8479 <= w8467 and not w8478;
w8480 <= not w1848 and w5431;
w8481 <= not w1992 and w4870;
w8482 <= not w1927 and w5342;
w8483 <= not w8481 and not w8482;
w8484 <= not w8480 and w8483;
w8485 <= w4873 and w5769;
w8486 <= w8484 and not w8485;
w8487 <= a(20) and not w8486;
w8488 <= not w8486 and not w8487;
w8489 <= a(20) and not w8487;
w8490 <= not w8488 and not w8489;
w8491 <= w8254 and not w8256;
w8492 <= not w8257 and not w8491;
w8493 <= not w8490 and w8492;
w8494 <= not w8490 and not w8493;
w8495 <= w8492 and not w8493;
w8496 <= not w8494 and not w8495;
w8497 <= not w1927 and w5431;
w8498 <= not w2087 and w4870;
w8499 <= not w1992 and w5342;
w8500 <= not w8498 and not w8499;
w8501 <= not w8497 and w8500;
w8502 <= w4873 and w6078;
w8503 <= w8501 and not w8502;
w8504 <= a(20) and not w8503;
w8505 <= not w8503 and not w8504;
w8506 <= a(20) and not w8504;
w8507 <= not w8505 and not w8506;
w8508 <= not w8249 and not w8253;
w8509 <= not w8252 and not w8253;
w8510 <= not w8508 and not w8509;
w8511 <= not w8507 and not w8510;
w8512 <= not w8507 and not w8511;
w8513 <= not w8510 and not w8511;
w8514 <= not w8512 and not w8513;
w8515 <= w8150 and w8247;
w8516 <= not w8248 and not w8515;
w8517 <= not w1992 and w5431;
w8518 <= not w2124 and w4870;
w8519 <= not w2087 and w5342;
w8520 <= not w8518 and not w8519;
w8521 <= not w8517 and w8520;
w8522 <= not w4873 and w8521;
w8523 <= not w6414 and w8521;
w8524 <= not w8522 and not w8523;
w8525 <= a(20) and not w8524;
w8526 <= not a(20) and w8524;
w8527 <= not w8525 and not w8526;
w8528 <= w8516 and not w8527;
w8529 <= w8243 and not w8245;
w8530 <= not w8246 and not w8529;
w8531 <= not w2087 and w5431;
w8532 <= not w2226 and w4870;
w8533 <= not w2124 and w5342;
w8534 <= not w8532 and not w8533;
w8535 <= not w8531 and w8534;
w8536 <= not w4873 and w8535;
w8537 <= not w6427 and w8535;
w8538 <= not w8536 and not w8537;
w8539 <= a(20) and not w8538;
w8540 <= not a(20) and w8538;
w8541 <= not w8539 and not w8540;
w8542 <= w8530 and not w8541;
w8543 <= w8182 and w8241;
w8544 <= not w8242 and not w8543;
w8545 <= not w2124 and w5431;
w8546 <= not w2323 and w4870;
w8547 <= not w2226 and w5342;
w8548 <= not w8546 and not w8547;
w8549 <= not w8545 and w8548;
w8550 <= not w4873 and w8549;
w8551 <= not w6057 and w8549;
w8552 <= not w8550 and not w8551;
w8553 <= a(20) and not w8552;
w8554 <= not a(20) and w8552;
w8555 <= not w8553 and not w8554;
w8556 <= w8544 and not w8555;
w8557 <= not w2226 and w5431;
w8558 <= not w2399 and w4870;
w8559 <= not w2323 and w5342;
w8560 <= not w8558 and not w8559;
w8561 <= not w8557 and w8560;
w8562 <= w4873 and w6476;
w8563 <= w8561 and not w8562;
w8564 <= a(20) and not w8563;
w8565 <= not w8563 and not w8564;
w8566 <= a(20) and not w8564;
w8567 <= not w8565 and not w8566;
w8568 <= w8237 and not w8239;
w8569 <= not w8240 and not w8568;
w8570 <= not w8567 and w8569;
w8571 <= not w8567 and not w8570;
w8572 <= w8569 and not w8570;
w8573 <= not w8571 and not w8572;
w8574 <= not w8224 and not w8236;
w8575 <= not w8235 and not w8236;
w8576 <= not w8574 and not w8575;
w8577 <= not w2323 and w5431;
w8578 <= not w2468 and w4870;
w8579 <= not w2399 and w5342;
w8580 <= not w8578 and not w8579;
w8581 <= not w8577 and w8580;
w8582 <= not w4873 and w8581;
w8583 <= not w6526 and w8581;
w8584 <= not w8582 and not w8583;
w8585 <= a(20) and not w8584;
w8586 <= not a(20) and w8584;
w8587 <= not w8585 and not w8586;
w8588 <= not w8576 and not w8587;
w8589 <= not w2399 and w5431;
w8590 <= not w2506 and w4870;
w8591 <= not w2468 and w5342;
w8592 <= not w8590 and not w8591;
w8593 <= not w8589 and w8592;
w8594 <= w4873 and w6581;
w8595 <= w8593 and not w8594;
w8596 <= a(20) and not w8595;
w8597 <= not w8595 and not w8596;
w8598 <= a(20) and not w8596;
w8599 <= not w8597 and not w8598;
w8600 <= not w8208 and w8219;
w8601 <= not w8220 and not w8600;
w8602 <= not w8599 and w8601;
w8603 <= not w8599 and not w8602;
w8604 <= w8601 and not w8602;
w8605 <= not w8603 and not w8604;
w8606 <= w8205 and not w8207;
w8607 <= not w8208 and not w8606;
w8608 <= not w2468 and w5431;
w8609 <= not w2609 and w4870;
w8610 <= not w2506 and w5342;
w8611 <= not w8609 and not w8610;
w8612 <= not w8608 and w8611;
w8613 <= not w4873 and w8612;
w8614 <= not w6630 and w8612;
w8615 <= not w8613 and not w8614;
w8616 <= a(20) and not w8615;
w8617 <= not a(20) and w8615;
w8618 <= not w8616 and not w8617;
w8619 <= w8607 and not w8618;
w8620 <= not w2764 and w5342;
w8621 <= not w2671 and w5431;
w8622 <= not w8620 and not w8621;
w8623 <= w4873 and not w7404;
w8624 <= w8622 and not w8623;
w8625 <= a(20) and not w8624;
w8626 <= a(20) and not w8625;
w8627 <= not w8624 and not w8625;
w8628 <= not w8626 and not w8627;
w8629 <= not w2764 and not w4868;
w8630 <= a(20) and not w8629;
w8631 <= not w8628 and w8630;
w8632 <= not w2609 and w5431;
w8633 <= not w2764 and w4870;
w8634 <= not w2671 and w5342;
w8635 <= not w8633 and not w8634;
w8636 <= not w8632 and w8635;
w8637 <= not w4873 and w8636;
w8638 <= not w6733 and w8636;
w8639 <= not w8637 and not w8638;
w8640 <= a(20) and not w8639;
w8641 <= not a(20) and w8639;
w8642 <= not w8640 and not w8641;
w8643 <= w8631 and not w8642;
w8644 <= w8206 and w8643;
w8645 <= w8643 and not w8644;
w8646 <= w8206 and not w8644;
w8647 <= not w8645 and not w8646;
w8648 <= not w2506 and w5431;
w8649 <= not w2671 and w4870;
w8650 <= not w2609 and w5342;
w8651 <= not w8649 and not w8650;
w8652 <= not w8648 and w8651;
w8653 <= w4873 and w6741;
w8654 <= w8652 and not w8653;
w8655 <= a(20) and not w8654;
w8656 <= a(20) and not w8655;
w8657 <= not w8654 and not w8655;
w8658 <= not w8656 and not w8657;
w8659 <= not w8647 and not w8658;
w8660 <= not w8644 and not w8659;
w8661 <= not w8607 and w8618;
w8662 <= not w8619 and not w8661;
w8663 <= not w8660 and w8662;
w8664 <= not w8619 and not w8663;
w8665 <= not w8605 and not w8664;
w8666 <= not w8602 and not w8665;
w8667 <= w8576 and w8587;
w8668 <= not w8588 and not w8667;
w8669 <= not w8666 and w8668;
w8670 <= not w8588 and not w8669;
w8671 <= not w8573 and not w8670;
w8672 <= not w8570 and not w8671;
w8673 <= w8544 and not w8556;
w8674 <= not w8555 and not w8556;
w8675 <= not w8673 and not w8674;
w8676 <= not w8672 and not w8675;
w8677 <= not w8556 and not w8676;
w8678 <= w8530 and not w8542;
w8679 <= not w8541 and not w8542;
w8680 <= not w8678 and not w8679;
w8681 <= not w8677 and not w8680;
w8682 <= not w8542 and not w8681;
w8683 <= not w8516 and w8527;
w8684 <= not w8528 and not w8683;
w8685 <= not w8682 and w8684;
w8686 <= not w8528 and not w8685;
w8687 <= not w8514 and not w8686;
w8688 <= not w8511 and not w8687;
w8689 <= not w8496 and not w8688;
w8690 <= not w8493 and not w8689;
w8691 <= w8467 and not w8479;
w8692 <= not w8478 and not w8479;
w8693 <= not w8691 and not w8692;
w8694 <= not w8690 and not w8693;
w8695 <= not w8479 and not w8694;
w8696 <= w8453 and not w8465;
w8697 <= not w8464 and not w8465;
w8698 <= not w8696 and not w8697;
w8699 <= not w8695 and not w8698;
w8700 <= not w8465 and not w8699;
w8701 <= w8439 and not w8451;
w8702 <= not w8450 and not w8451;
w8703 <= not w8701 and not w8702;
w8704 <= not w8700 and not w8703;
w8705 <= not w8451 and not w8704;
w8706 <= w8425 and not w8437;
w8707 <= not w8436 and not w8437;
w8708 <= not w8706 and not w8707;
w8709 <= not w8705 and not w8708;
w8710 <= not w8437 and not w8709;
w8711 <= w8411 and not w8423;
w8712 <= not w8422 and not w8423;
w8713 <= not w8711 and not w8712;
w8714 <= not w8710 and not w8713;
w8715 <= not w8423 and not w8714;
w8716 <= w8397 and not w8409;
w8717 <= not w8408 and not w8409;
w8718 <= not w8716 and not w8717;
w8719 <= not w8715 and not w8718;
w8720 <= not w8409 and not w8719;
w8721 <= w8383 and not w8395;
w8722 <= not w8394 and not w8395;
w8723 <= not w8721 and not w8722;
w8724 <= not w8720 and not w8723;
w8725 <= not w8395 and not w8724;
w8726 <= w8286 and not w8288;
w8727 <= not w8289 and not w8726;
w8728 <= not w8725 and w8727;
w8729 <= not w802 and w6168;
w8730 <= not w995 and w5598;
w8731 <= not w893 and w5874;
w8732 <= not w8730 and not w8731;
w8733 <= not w8729 and w8732;
w8734 <= w4139 and w5601;
w8735 <= w8733 and not w8734;
w8736 <= a(17) and not w8735;
w8737 <= not w8735 and not w8736;
w8738 <= a(17) and not w8736;
w8739 <= not w8737 and not w8738;
w8740 <= w8725 and not w8727;
w8741 <= not w8728 and not w8740;
w8742 <= not w8739 and w8741;
w8743 <= not w8728 and not w8742;
w8744 <= not w8381 and not w8743;
w8745 <= w8381 and w8743;
w8746 <= not w8744 and not w8745;
w8747 <= not w2947 and w7036;
w8748 <= not w522 and w6337;
w8749 <= not w327 and w6886;
w8750 <= not w8748 and not w8749;
w8751 <= not w8747 and w8750;
w8752 <= w2953 and w6332;
w8753 <= w8751 and not w8752;
w8754 <= a(14) and not w8753;
w8755 <= a(14) and not w8754;
w8756 <= not w8753 and not w8754;
w8757 <= not w8755 and not w8756;
w8758 <= w8746 and not w8757;
w8759 <= not w8744 and not w8758;
w8760 <= not w8378 and not w8759;
w8761 <= w8378 and w8759;
w8762 <= not w8760 and not w8761;
w8763 <= not w3740 and w7918;
w8764 <= not w3540 and w7226;
w8765 <= not w3391 and w7567;
w8766 <= not w8764 and not w8765;
w8767 <= not w8763 and w8766;
w8768 <= w3753 and w7229;
w8769 <= w8767 and not w8768;
w8770 <= a(11) and not w8769;
w8771 <= a(11) and not w8770;
w8772 <= not w8769 and not w8770;
w8773 <= not w8771 and not w8772;
w8774 <= w8762 and not w8773;
w8775 <= not w8760 and not w8774;
w8776 <= not w3899 and w7918;
w8777 <= not w3391 and w7226;
w8778 <= not w3740 and w7567;
w8779 <= not w8777 and not w8778;
w8780 <= not w8776 and w8779;
w8781 <= not w7229 and w8780;
w8782 <= not w4493 and w8780;
w8783 <= not w8781 and not w8782;
w8784 <= a(11) and not w8783;
w8785 <= not a(11) and w8783;
w8786 <= not w8784 and not w8785;
w8787 <= not w8775 and not w8786;
w8788 <= w8775 and w8786;
w8789 <= not w8787 and not w8788;
w8790 <= w8322 and not w8324;
w8791 <= not w8325 and not w8790;
w8792 <= w8789 and w8791;
w8793 <= not w8787 and not w8792;
w8794 <= not w3812 and w8353;
w8795 <= not w8345 and w8351;
w8796 <= not w4450 and w8795;
w8797 <= not w8794 and not w8796;
w8798 <= not w8356 and w8797;
w8799 <= not w4544 and w8797;
w8800 <= not w8798 and not w8799;
w8801 <= a(8) and not w8800;
w8802 <= not a(8) and w8800;
w8803 <= not w8801 and not w8802;
w8804 <= not w8793 and not w8803;
w8805 <= w8329 and not w8341;
w8806 <= not w8340 and not w8341;
w8807 <= not w8805 and not w8806;
w8808 <= w8793 and w8803;
w8809 <= not w8804 and not w8808;
w8810 <= not w8807 and w8809;
w8811 <= not w8804 and not w8810;
w8812 <= not w8375 and not w8811;
w8813 <= w8375 and w8811;
w8814 <= not w8812 and not w8813;
w8815 <= w8762 and not w8774;
w8816 <= not w8773 and not w8774;
w8817 <= not w8815 and not w8816;
w8818 <= w8746 and not w8758;
w8819 <= not w8757 and not w8758;
w8820 <= not w8818 and not w8819;
w8821 <= not w893 and w6168;
w8822 <= not w1113 and w5598;
w8823 <= not w995 and w5874;
w8824 <= not w8822 and not w8823;
w8825 <= not w8821 and w8824;
w8826 <= w4568 and w5601;
w8827 <= w8825 and not w8826;
w8828 <= a(17) and not w8827;
w8829 <= not w8827 and not w8828;
w8830 <= a(17) and not w8828;
w8831 <= not w8829 and not w8830;
w8832 <= not w8720 and not w8724;
w8833 <= not w8723 and not w8724;
w8834 <= not w8832 and not w8833;
w8835 <= not w8831 and not w8834;
w8836 <= not w8831 and not w8835;
w8837 <= not w8834 and not w8835;
w8838 <= not w8836 and not w8837;
w8839 <= not w995 and w6168;
w8840 <= not w1170 and w5598;
w8841 <= not w1113 and w5874;
w8842 <= not w8840 and not w8841;
w8843 <= not w8839 and w8842;
w8844 <= w4364 and w5601;
w8845 <= w8843 and not w8844;
w8846 <= a(17) and not w8845;
w8847 <= not w8845 and not w8846;
w8848 <= a(17) and not w8846;
w8849 <= not w8847 and not w8848;
w8850 <= not w8715 and not w8719;
w8851 <= not w8718 and not w8719;
w8852 <= not w8850 and not w8851;
w8853 <= not w8849 and not w8852;
w8854 <= not w8849 and not w8853;
w8855 <= not w8852 and not w8853;
w8856 <= not w8854 and not w8855;
w8857 <= not w1113 and w6168;
w8858 <= not w1299 and w5598;
w8859 <= not w1170 and w5874;
w8860 <= not w8858 and not w8859;
w8861 <= not w8857 and w8860;
w8862 <= w4796 and w5601;
w8863 <= w8861 and not w8862;
w8864 <= a(17) and not w8863;
w8865 <= not w8863 and not w8864;
w8866 <= a(17) and not w8864;
w8867 <= not w8865 and not w8866;
w8868 <= not w8710 and not w8714;
w8869 <= not w8713 and not w8714;
w8870 <= not w8868 and not w8869;
w8871 <= not w8867 and not w8870;
w8872 <= not w8867 and not w8871;
w8873 <= not w8870 and not w8871;
w8874 <= not w8872 and not w8873;
w8875 <= not w1170 and w6168;
w8876 <= not w1407 and w5598;
w8877 <= not w1299 and w5874;
w8878 <= not w8876 and not w8877;
w8879 <= not w8875 and w8878;
w8880 <= w4783 and w5601;
w8881 <= w8879 and not w8880;
w8882 <= a(17) and not w8881;
w8883 <= not w8881 and not w8882;
w8884 <= a(17) and not w8882;
w8885 <= not w8883 and not w8884;
w8886 <= not w8705 and not w8709;
w8887 <= not w8708 and not w8709;
w8888 <= not w8886 and not w8887;
w8889 <= not w8885 and not w8888;
w8890 <= not w8885 and not w8889;
w8891 <= not w8888 and not w8889;
w8892 <= not w8890 and not w8891;
w8893 <= not w1299 and w6168;
w8894 <= not w1507 and w5598;
w8895 <= not w1407 and w5874;
w8896 <= not w8894 and not w8895;
w8897 <= not w8893 and w8896;
w8898 <= w5049 and w5601;
w8899 <= w8897 and not w8898;
w8900 <= a(17) and not w8899;
w8901 <= not w8899 and not w8900;
w8902 <= a(17) and not w8900;
w8903 <= not w8901 and not w8902;
w8904 <= not w8700 and not w8704;
w8905 <= not w8703 and not w8704;
w8906 <= not w8904 and not w8905;
w8907 <= not w8903 and not w8906;
w8908 <= not w8903 and not w8907;
w8909 <= not w8906 and not w8907;
w8910 <= not w8908 and not w8909;
w8911 <= not w1407 and w6168;
w8912 <= not w1600 and w5598;
w8913 <= not w1507 and w5874;
w8914 <= not w8912 and not w8913;
w8915 <= not w8911 and w8914;
w8916 <= w5074 and w5601;
w8917 <= w8915 and not w8916;
w8918 <= a(17) and not w8917;
w8919 <= not w8917 and not w8918;
w8920 <= a(17) and not w8918;
w8921 <= not w8919 and not w8920;
w8922 <= not w8695 and not w8699;
w8923 <= not w8698 and not w8699;
w8924 <= not w8922 and not w8923;
w8925 <= not w8921 and not w8924;
w8926 <= not w8921 and not w8925;
w8927 <= not w8924 and not w8925;
w8928 <= not w8926 and not w8927;
w8929 <= not w1507 and w6168;
w8930 <= not w1714 and w5598;
w8931 <= not w1600 and w5874;
w8932 <= not w8930 and not w8931;
w8933 <= not w8929 and w8932;
w8934 <= w5496 and w5601;
w8935 <= w8933 and not w8934;
w8936 <= a(17) and not w8935;
w8937 <= not w8935 and not w8936;
w8938 <= a(17) and not w8936;
w8939 <= not w8937 and not w8938;
w8940 <= not w8690 and not w8694;
w8941 <= not w8693 and not w8694;
w8942 <= not w8940 and not w8941;
w8943 <= not w8939 and not w8942;
w8944 <= not w8939 and not w8943;
w8945 <= not w8942 and not w8943;
w8946 <= not w8944 and not w8945;
w8947 <= w8496 and w8688;
w8948 <= not w8689 and not w8947;
w8949 <= not w1600 and w6168;
w8950 <= not w1812 and w5598;
w8951 <= not w1714 and w5874;
w8952 <= not w8950 and not w8951;
w8953 <= not w8949 and w8952;
w8954 <= not w5601 and w8953;
w8955 <= not w5263 and w8953;
w8956 <= not w8954 and not w8955;
w8957 <= a(17) and not w8956;
w8958 <= not a(17) and w8956;
w8959 <= not w8957 and not w8958;
w8960 <= w8948 and not w8959;
w8961 <= w8514 and w8686;
w8962 <= not w8687 and not w8961;
w8963 <= not w1714 and w6168;
w8964 <= not w1848 and w5598;
w8965 <= not w1812 and w5874;
w8966 <= not w8964 and not w8965;
w8967 <= not w8963 and w8966;
w8968 <= not w5601 and w8967;
w8969 <= not w5786 and w8967;
w8970 <= not w8968 and not w8969;
w8971 <= a(17) and not w8970;
w8972 <= not a(17) and w8970;
w8973 <= not w8971 and not w8972;
w8974 <= w8962 and not w8973;
w8975 <= not w1812 and w6168;
w8976 <= not w1927 and w5598;
w8977 <= not w1848 and w5874;
w8978 <= not w8976 and not w8977;
w8979 <= not w8975 and w8978;
w8980 <= w5601 and w5942;
w8981 <= w8979 and not w8980;
w8982 <= a(17) and not w8981;
w8983 <= not w8981 and not w8982;
w8984 <= a(17) and not w8982;
w8985 <= not w8983 and not w8984;
w8986 <= w8682 and not w8684;
w8987 <= not w8685 and not w8986;
w8988 <= not w8985 and w8987;
w8989 <= not w8985 and not w8988;
w8990 <= w8987 and not w8988;
w8991 <= not w8989 and not w8990;
w8992 <= not w1848 and w6168;
w8993 <= not w1992 and w5598;
w8994 <= not w1927 and w5874;
w8995 <= not w8993 and not w8994;
w8996 <= not w8992 and w8995;
w8997 <= w5601 and w5769;
w8998 <= w8996 and not w8997;
w8999 <= a(17) and not w8998;
w9000 <= not w8998 and not w8999;
w9001 <= a(17) and not w8999;
w9002 <= not w9000 and not w9001;
w9003 <= not w8677 and not w8681;
w9004 <= not w8680 and not w8681;
w9005 <= not w9003 and not w9004;
w9006 <= not w9002 and not w9005;
w9007 <= not w9002 and not w9006;
w9008 <= not w9005 and not w9006;
w9009 <= not w9007 and not w9008;
w9010 <= not w1927 and w6168;
w9011 <= not w2087 and w5598;
w9012 <= not w1992 and w5874;
w9013 <= not w9011 and not w9012;
w9014 <= not w9010 and w9013;
w9015 <= w5601 and w6078;
w9016 <= w9014 and not w9015;
w9017 <= a(17) and not w9016;
w9018 <= not w9016 and not w9017;
w9019 <= a(17) and not w9017;
w9020 <= not w9018 and not w9019;
w9021 <= not w8672 and not w8676;
w9022 <= not w8675 and not w8676;
w9023 <= not w9021 and not w9022;
w9024 <= not w9020 and not w9023;
w9025 <= not w9020 and not w9024;
w9026 <= not w9023 and not w9024;
w9027 <= not w9025 and not w9026;
w9028 <= w8573 and w8670;
w9029 <= not w8671 and not w9028;
w9030 <= not w1992 and w6168;
w9031 <= not w2124 and w5598;
w9032 <= not w2087 and w5874;
w9033 <= not w9031 and not w9032;
w9034 <= not w9030 and w9033;
w9035 <= not w5601 and w9034;
w9036 <= not w6414 and w9034;
w9037 <= not w9035 and not w9036;
w9038 <= a(17) and not w9037;
w9039 <= not a(17) and w9037;
w9040 <= not w9038 and not w9039;
w9041 <= w9029 and not w9040;
w9042 <= w8666 and not w8668;
w9043 <= not w8669 and not w9042;
w9044 <= not w2087 and w6168;
w9045 <= not w2226 and w5598;
w9046 <= not w2124 and w5874;
w9047 <= not w9045 and not w9046;
w9048 <= not w9044 and w9047;
w9049 <= not w5601 and w9048;
w9050 <= not w6427 and w9048;
w9051 <= not w9049 and not w9050;
w9052 <= a(17) and not w9051;
w9053 <= not a(17) and w9051;
w9054 <= not w9052 and not w9053;
w9055 <= w9043 and not w9054;
w9056 <= w8605 and w8664;
w9057 <= not w8665 and not w9056;
w9058 <= not w2124 and w6168;
w9059 <= not w2323 and w5598;
w9060 <= not w2226 and w5874;
w9061 <= not w9059 and not w9060;
w9062 <= not w9058 and w9061;
w9063 <= not w5601 and w9062;
w9064 <= not w6057 and w9062;
w9065 <= not w9063 and not w9064;
w9066 <= a(17) and not w9065;
w9067 <= not a(17) and w9065;
w9068 <= not w9066 and not w9067;
w9069 <= w9057 and not w9068;
w9070 <= not w2226 and w6168;
w9071 <= not w2399 and w5598;
w9072 <= not w2323 and w5874;
w9073 <= not w9071 and not w9072;
w9074 <= not w9070 and w9073;
w9075 <= w5601 and w6476;
w9076 <= w9074 and not w9075;
w9077 <= a(17) and not w9076;
w9078 <= not w9076 and not w9077;
w9079 <= a(17) and not w9077;
w9080 <= not w9078 and not w9079;
w9081 <= w8660 and not w8662;
w9082 <= not w8663 and not w9081;
w9083 <= not w9080 and w9082;
w9084 <= not w9080 and not w9083;
w9085 <= w9082 and not w9083;
w9086 <= not w9084 and not w9085;
w9087 <= not w8647 and not w8659;
w9088 <= not w8658 and not w8659;
w9089 <= not w9087 and not w9088;
w9090 <= not w2323 and w6168;
w9091 <= not w2468 and w5598;
w9092 <= not w2399 and w5874;
w9093 <= not w9091 and not w9092;
w9094 <= not w9090 and w9093;
w9095 <= not w5601 and w9094;
w9096 <= not w6526 and w9094;
w9097 <= not w9095 and not w9096;
w9098 <= a(17) and not w9097;
w9099 <= not a(17) and w9097;
w9100 <= not w9098 and not w9099;
w9101 <= not w9089 and not w9100;
w9102 <= not w2399 and w6168;
w9103 <= not w2506 and w5598;
w9104 <= not w2468 and w5874;
w9105 <= not w9103 and not w9104;
w9106 <= not w9102 and w9105;
w9107 <= w5601 and w6581;
w9108 <= w9106 and not w9107;
w9109 <= a(17) and not w9108;
w9110 <= not w9108 and not w9109;
w9111 <= a(17) and not w9109;
w9112 <= not w9110 and not w9111;
w9113 <= not w8631 and w8642;
w9114 <= not w8643 and not w9113;
w9115 <= not w9112 and w9114;
w9116 <= not w9112 and not w9115;
w9117 <= w9114 and not w9115;
w9118 <= not w9116 and not w9117;
w9119 <= w8628 and not w8630;
w9120 <= not w8631 and not w9119;
w9121 <= not w2468 and w6168;
w9122 <= not w2609 and w5598;
w9123 <= not w2506 and w5874;
w9124 <= not w9122 and not w9123;
w9125 <= not w9121 and w9124;
w9126 <= not w5601 and w9125;
w9127 <= not w6630 and w9125;
w9128 <= not w9126 and not w9127;
w9129 <= a(17) and not w9128;
w9130 <= not a(17) and w9128;
w9131 <= not w9129 and not w9130;
w9132 <= w9120 and not w9131;
w9133 <= not w2764 and w5874;
w9134 <= not w2671 and w6168;
w9135 <= not w9133 and not w9134;
w9136 <= w5601 and not w7404;
w9137 <= w9135 and not w9136;
w9138 <= a(17) and not w9137;
w9139 <= a(17) and not w9138;
w9140 <= not w9137 and not w9138;
w9141 <= not w9139 and not w9140;
w9142 <= not w2764 and not w5593;
w9143 <= a(17) and not w9142;
w9144 <= not w9141 and w9143;
w9145 <= not w2609 and w6168;
w9146 <= not w2764 and w5598;
w9147 <= not w2671 and w5874;
w9148 <= not w9146 and not w9147;
w9149 <= not w9145 and w9148;
w9150 <= not w5601 and w9149;
w9151 <= not w6733 and w9149;
w9152 <= not w9150 and not w9151;
w9153 <= a(17) and not w9152;
w9154 <= not a(17) and w9152;
w9155 <= not w9153 and not w9154;
w9156 <= w9144 and not w9155;
w9157 <= w8629 and w9156;
w9158 <= w9156 and not w9157;
w9159 <= w8629 and not w9157;
w9160 <= not w9158 and not w9159;
w9161 <= not w2506 and w6168;
w9162 <= not w2671 and w5598;
w9163 <= not w2609 and w5874;
w9164 <= not w9162 and not w9163;
w9165 <= not w9161 and w9164;
w9166 <= w5601 and w6741;
w9167 <= w9165 and not w9166;
w9168 <= a(17) and not w9167;
w9169 <= a(17) and not w9168;
w9170 <= not w9167 and not w9168;
w9171 <= not w9169 and not w9170;
w9172 <= not w9160 and not w9171;
w9173 <= not w9157 and not w9172;
w9174 <= not w9120 and w9131;
w9175 <= not w9132 and not w9174;
w9176 <= not w9173 and w9175;
w9177 <= not w9132 and not w9176;
w9178 <= not w9118 and not w9177;
w9179 <= not w9115 and not w9178;
w9180 <= w9089 and w9100;
w9181 <= not w9101 and not w9180;
w9182 <= not w9179 and w9181;
w9183 <= not w9101 and not w9182;
w9184 <= not w9086 and not w9183;
w9185 <= not w9083 and not w9184;
w9186 <= w9057 and not w9069;
w9187 <= not w9068 and not w9069;
w9188 <= not w9186 and not w9187;
w9189 <= not w9185 and not w9188;
w9190 <= not w9069 and not w9189;
w9191 <= w9043 and not w9055;
w9192 <= not w9054 and not w9055;
w9193 <= not w9191 and not w9192;
w9194 <= not w9190 and not w9193;
w9195 <= not w9055 and not w9194;
w9196 <= not w9029 and w9040;
w9197 <= not w9041 and not w9196;
w9198 <= not w9195 and w9197;
w9199 <= not w9041 and not w9198;
w9200 <= not w9027 and not w9199;
w9201 <= not w9024 and not w9200;
w9202 <= not w9009 and not w9201;
w9203 <= not w9006 and not w9202;
w9204 <= not w8991 and not w9203;
w9205 <= not w8988 and not w9204;
w9206 <= w8962 and not w8974;
w9207 <= not w8973 and not w8974;
w9208 <= not w9206 and not w9207;
w9209 <= not w9205 and not w9208;
w9210 <= not w8974 and not w9209;
w9211 <= not w8948 and w8959;
w9212 <= not w8960 and not w9211;
w9213 <= not w9210 and w9212;
w9214 <= not w8960 and not w9213;
w9215 <= not w8946 and not w9214;
w9216 <= not w8943 and not w9215;
w9217 <= not w8928 and not w9216;
w9218 <= not w8925 and not w9217;
w9219 <= not w8910 and not w9218;
w9220 <= not w8907 and not w9219;
w9221 <= not w8892 and not w9220;
w9222 <= not w8889 and not w9221;
w9223 <= not w8874 and not w9222;
w9224 <= not w8871 and not w9223;
w9225 <= not w8856 and not w9224;
w9226 <= not w8853 and not w9225;
w9227 <= not w8838 and not w9226;
w9228 <= not w8835 and not w9227;
w9229 <= w8739 and not w8741;
w9230 <= not w8742 and not w9229;
w9231 <= not w9228 and w9230;
w9232 <= not w327 and w7036;
w9233 <= not w645 and w6337;
w9234 <= not w522 and w6886;
w9235 <= not w9233 and not w9234;
w9236 <= not w9232 and w9235;
w9237 <= w3282 and w6332;
w9238 <= w9236 and not w9237;
w9239 <= a(14) and not w9238;
w9240 <= not w9238 and not w9239;
w9241 <= a(14) and not w9239;
w9242 <= not w9240 and not w9241;
w9243 <= w9228 and not w9230;
w9244 <= not w9231 and not w9243;
w9245 <= not w9242 and w9244;
w9246 <= not w9231 and not w9245;
w9247 <= not w8820 and not w9246;
w9248 <= w8820 and w9246;
w9249 <= not w9247 and not w9248;
w9250 <= not w3391 and w7918;
w9251 <= not w3474 and w7226;
w9252 <= not w3540 and w7567;
w9253 <= not w9251 and not w9252;
w9254 <= not w9250 and w9253;
w9255 <= w3562 and w7229;
w9256 <= w9254 and not w9255;
w9257 <= a(11) and not w9256;
w9258 <= a(11) and not w9257;
w9259 <= not w9256 and not w9257;
w9260 <= not w9258 and not w9259;
w9261 <= w9249 and not w9260;
w9262 <= not w9247 and not w9261;
w9263 <= not w8817 and not w9262;
w9264 <= w8817 and w9262;
w9265 <= not w9263 and not w9264;
w9266 <= w8348 and not w8351;
w9267 <= not w3812 and w9266;
w9268 <= not w3899 and w8353;
w9269 <= not w3980 and w8795;
w9270 <= not w9268 and not w9269;
w9271 <= not w9267 and w9270;
w9272 <= w4002 and w8356;
w9273 <= w9271 and not w9272;
w9274 <= a(8) and not w9273;
w9275 <= a(8) and not w9274;
w9276 <= not w9273 and not w9274;
w9277 <= not w9275 and not w9276;
w9278 <= w9265 and not w9277;
w9279 <= not w9263 and not w9278;
w9280 <= not w4450 and w9266;
w9281 <= not w3980 and w8353;
w9282 <= not w3812 and w8795;
w9283 <= not w9281 and not w9282;
w9284 <= not w9280 and w9283;
w9285 <= not w8356 and w9284;
w9286 <= not w4650 and w9284;
w9287 <= not w9285 and not w9286;
w9288 <= a(8) and not w9287;
w9289 <= not a(8) and w9287;
w9290 <= not w9288 and not w9289;
w9291 <= not w9279 and not w9290;
w9292 <= not w9279 and not w9291;
w9293 <= not w9290 and not w9291;
w9294 <= not w9292 and not w9293;
w9295 <= not w8789 and not w8791;
w9296 <= not w8792 and not w9295;
w9297 <= not w9294 and w9296;
w9298 <= not w9291 and not w9297;
w9299 <= w8807 and not w8809;
w9300 <= not w8810 and not w9299;
w9301 <= not w9298 and w9300;
w9302 <= w9249 and not w9261;
w9303 <= not w9260 and not w9261;
w9304 <= not w9302 and not w9303;
w9305 <= w8838 and w9226;
w9306 <= not w9227 and not w9305;
w9307 <= not w522 and w7036;
w9308 <= not w802 and w6337;
w9309 <= not w645 and w6886;
w9310 <= not w9308 and not w9309;
w9311 <= not w9307 and w9310;
w9312 <= not w6332 and w9311;
w9313 <= not w3266 and w9311;
w9314 <= not w9312 and not w9313;
w9315 <= a(14) and not w9314;
w9316 <= not a(14) and w9314;
w9317 <= not w9315 and not w9316;
w9318 <= w9306 and not w9317;
w9319 <= w8856 and w9224;
w9320 <= not w9225 and not w9319;
w9321 <= not w645 and w7036;
w9322 <= not w893 and w6337;
w9323 <= not w802 and w6886;
w9324 <= not w9322 and not w9323;
w9325 <= not w9321 and w9324;
w9326 <= not w6332 and w9325;
w9327 <= not w4114 and w9325;
w9328 <= not w9326 and not w9327;
w9329 <= a(14) and not w9328;
w9330 <= not a(14) and w9328;
w9331 <= not w9329 and not w9330;
w9332 <= w9320 and not w9331;
w9333 <= w8874 and w9222;
w9334 <= not w9223 and not w9333;
w9335 <= not w802 and w7036;
w9336 <= not w995 and w6337;
w9337 <= not w893 and w6886;
w9338 <= not w9336 and not w9337;
w9339 <= not w9335 and w9338;
w9340 <= not w6332 and w9339;
w9341 <= not w4139 and w9339;
w9342 <= not w9340 and not w9341;
w9343 <= a(14) and not w9342;
w9344 <= not a(14) and w9342;
w9345 <= not w9343 and not w9344;
w9346 <= w9334 and not w9345;
w9347 <= w8892 and w9220;
w9348 <= not w9221 and not w9347;
w9349 <= not w893 and w7036;
w9350 <= not w1113 and w6337;
w9351 <= not w995 and w6886;
w9352 <= not w9350 and not w9351;
w9353 <= not w9349 and w9352;
w9354 <= not w6332 and w9353;
w9355 <= not w4568 and w9353;
w9356 <= not w9354 and not w9355;
w9357 <= a(14) and not w9356;
w9358 <= not a(14) and w9356;
w9359 <= not w9357 and not w9358;
w9360 <= w9348 and not w9359;
w9361 <= w8910 and w9218;
w9362 <= not w9219 and not w9361;
w9363 <= not w995 and w7036;
w9364 <= not w1170 and w6337;
w9365 <= not w1113 and w6886;
w9366 <= not w9364 and not w9365;
w9367 <= not w9363 and w9366;
w9368 <= not w6332 and w9367;
w9369 <= not w4364 and w9367;
w9370 <= not w9368 and not w9369;
w9371 <= a(14) and not w9370;
w9372 <= not a(14) and w9370;
w9373 <= not w9371 and not w9372;
w9374 <= w9362 and not w9373;
w9375 <= w8928 and w9216;
w9376 <= not w9217 and not w9375;
w9377 <= not w1113 and w7036;
w9378 <= not w1299 and w6337;
w9379 <= not w1170 and w6886;
w9380 <= not w9378 and not w9379;
w9381 <= not w9377 and w9380;
w9382 <= not w6332 and w9381;
w9383 <= not w4796 and w9381;
w9384 <= not w9382 and not w9383;
w9385 <= a(14) and not w9384;
w9386 <= not a(14) and w9384;
w9387 <= not w9385 and not w9386;
w9388 <= w9376 and not w9387;
w9389 <= w8946 and w9214;
w9390 <= not w9215 and not w9389;
w9391 <= not w1170 and w7036;
w9392 <= not w1407 and w6337;
w9393 <= not w1299 and w6886;
w9394 <= not w9392 and not w9393;
w9395 <= not w9391 and w9394;
w9396 <= not w6332 and w9395;
w9397 <= not w4783 and w9395;
w9398 <= not w9396 and not w9397;
w9399 <= a(14) and not w9398;
w9400 <= not a(14) and w9398;
w9401 <= not w9399 and not w9400;
w9402 <= w9390 and not w9401;
w9403 <= not w1299 and w7036;
w9404 <= not w1507 and w6337;
w9405 <= not w1407 and w6886;
w9406 <= not w9404 and not w9405;
w9407 <= not w9403 and w9406;
w9408 <= w5049 and w6332;
w9409 <= w9407 and not w9408;
w9410 <= a(14) and not w9409;
w9411 <= not w9409 and not w9410;
w9412 <= a(14) and not w9410;
w9413 <= not w9411 and not w9412;
w9414 <= w9210 and not w9212;
w9415 <= not w9213 and not w9414;
w9416 <= not w9413 and w9415;
w9417 <= not w9413 and not w9416;
w9418 <= w9415 and not w9416;
w9419 <= not w9417 and not w9418;
w9420 <= not w1407 and w7036;
w9421 <= not w1600 and w6337;
w9422 <= not w1507 and w6886;
w9423 <= not w9421 and not w9422;
w9424 <= not w9420 and w9423;
w9425 <= w5074 and w6332;
w9426 <= w9424 and not w9425;
w9427 <= a(14) and not w9426;
w9428 <= not w9426 and not w9427;
w9429 <= a(14) and not w9427;
w9430 <= not w9428 and not w9429;
w9431 <= not w9205 and not w9209;
w9432 <= not w9208 and not w9209;
w9433 <= not w9431 and not w9432;
w9434 <= not w9430 and not w9433;
w9435 <= not w9430 and not w9434;
w9436 <= not w9433 and not w9434;
w9437 <= not w9435 and not w9436;
w9438 <= w8991 and w9203;
w9439 <= not w9204 and not w9438;
w9440 <= not w1507 and w7036;
w9441 <= not w1714 and w6337;
w9442 <= not w1600 and w6886;
w9443 <= not w9441 and not w9442;
w9444 <= not w9440 and w9443;
w9445 <= not w6332 and w9444;
w9446 <= not w5496 and w9444;
w9447 <= not w9445 and not w9446;
w9448 <= a(14) and not w9447;
w9449 <= not a(14) and w9447;
w9450 <= not w9448 and not w9449;
w9451 <= w9439 and not w9450;
w9452 <= w9009 and w9201;
w9453 <= not w9202 and not w9452;
w9454 <= not w1600 and w7036;
w9455 <= not w1812 and w6337;
w9456 <= not w1714 and w6886;
w9457 <= not w9455 and not w9456;
w9458 <= not w9454 and w9457;
w9459 <= not w6332 and w9458;
w9460 <= not w5263 and w9458;
w9461 <= not w9459 and not w9460;
w9462 <= a(14) and not w9461;
w9463 <= not a(14) and w9461;
w9464 <= not w9462 and not w9463;
w9465 <= w9453 and not w9464;
w9466 <= w9027 and w9199;
w9467 <= not w9200 and not w9466;
w9468 <= not w1714 and w7036;
w9469 <= not w1848 and w6337;
w9470 <= not w1812 and w6886;
w9471 <= not w9469 and not w9470;
w9472 <= not w9468 and w9471;
w9473 <= not w6332 and w9472;
w9474 <= not w5786 and w9472;
w9475 <= not w9473 and not w9474;
w9476 <= a(14) and not w9475;
w9477 <= not a(14) and w9475;
w9478 <= not w9476 and not w9477;
w9479 <= w9467 and not w9478;
w9480 <= not w1812 and w7036;
w9481 <= not w1927 and w6337;
w9482 <= not w1848 and w6886;
w9483 <= not w9481 and not w9482;
w9484 <= not w9480 and w9483;
w9485 <= w5942 and w6332;
w9486 <= w9484 and not w9485;
w9487 <= a(14) and not w9486;
w9488 <= not w9486 and not w9487;
w9489 <= a(14) and not w9487;
w9490 <= not w9488 and not w9489;
w9491 <= w9195 and not w9197;
w9492 <= not w9198 and not w9491;
w9493 <= not w9490 and w9492;
w9494 <= not w9490 and not w9493;
w9495 <= w9492 and not w9493;
w9496 <= not w9494 and not w9495;
w9497 <= not w1848 and w7036;
w9498 <= not w1992 and w6337;
w9499 <= not w1927 and w6886;
w9500 <= not w9498 and not w9499;
w9501 <= not w9497 and w9500;
w9502 <= w5769 and w6332;
w9503 <= w9501 and not w9502;
w9504 <= a(14) and not w9503;
w9505 <= not w9503 and not w9504;
w9506 <= a(14) and not w9504;
w9507 <= not w9505 and not w9506;
w9508 <= not w9190 and not w9194;
w9509 <= not w9193 and not w9194;
w9510 <= not w9508 and not w9509;
w9511 <= not w9507 and not w9510;
w9512 <= not w9507 and not w9511;
w9513 <= not w9510 and not w9511;
w9514 <= not w9512 and not w9513;
w9515 <= not w1927 and w7036;
w9516 <= not w2087 and w6337;
w9517 <= not w1992 and w6886;
w9518 <= not w9516 and not w9517;
w9519 <= not w9515 and w9518;
w9520 <= w6078 and w6332;
w9521 <= w9519 and not w9520;
w9522 <= a(14) and not w9521;
w9523 <= not w9521 and not w9522;
w9524 <= a(14) and not w9522;
w9525 <= not w9523 and not w9524;
w9526 <= not w9185 and not w9189;
w9527 <= not w9188 and not w9189;
w9528 <= not w9526 and not w9527;
w9529 <= not w9525 and not w9528;
w9530 <= not w9525 and not w9529;
w9531 <= not w9528 and not w9529;
w9532 <= not w9530 and not w9531;
w9533 <= w9086 and w9183;
w9534 <= not w9184 and not w9533;
w9535 <= not w1992 and w7036;
w9536 <= not w2124 and w6337;
w9537 <= not w2087 and w6886;
w9538 <= not w9536 and not w9537;
w9539 <= not w9535 and w9538;
w9540 <= not w6332 and w9539;
w9541 <= not w6414 and w9539;
w9542 <= not w9540 and not w9541;
w9543 <= a(14) and not w9542;
w9544 <= not a(14) and w9542;
w9545 <= not w9543 and not w9544;
w9546 <= w9534 and not w9545;
w9547 <= w9179 and not w9181;
w9548 <= not w9182 and not w9547;
w9549 <= not w2087 and w7036;
w9550 <= not w2226 and w6337;
w9551 <= not w2124 and w6886;
w9552 <= not w9550 and not w9551;
w9553 <= not w9549 and w9552;
w9554 <= not w6332 and w9553;
w9555 <= not w6427 and w9553;
w9556 <= not w9554 and not w9555;
w9557 <= a(14) and not w9556;
w9558 <= not a(14) and w9556;
w9559 <= not w9557 and not w9558;
w9560 <= w9548 and not w9559;
w9561 <= w9118 and w9177;
w9562 <= not w9178 and not w9561;
w9563 <= not w2124 and w7036;
w9564 <= not w2323 and w6337;
w9565 <= not w2226 and w6886;
w9566 <= not w9564 and not w9565;
w9567 <= not w9563 and w9566;
w9568 <= not w6332 and w9567;
w9569 <= not w6057 and w9567;
w9570 <= not w9568 and not w9569;
w9571 <= a(14) and not w9570;
w9572 <= not a(14) and w9570;
w9573 <= not w9571 and not w9572;
w9574 <= w9562 and not w9573;
w9575 <= not w2226 and w7036;
w9576 <= not w2399 and w6337;
w9577 <= not w2323 and w6886;
w9578 <= not w9576 and not w9577;
w9579 <= not w9575 and w9578;
w9580 <= w6332 and w6476;
w9581 <= w9579 and not w9580;
w9582 <= a(14) and not w9581;
w9583 <= not w9581 and not w9582;
w9584 <= a(14) and not w9582;
w9585 <= not w9583 and not w9584;
w9586 <= w9173 and not w9175;
w9587 <= not w9176 and not w9586;
w9588 <= not w9585 and w9587;
w9589 <= not w9585 and not w9588;
w9590 <= w9587 and not w9588;
w9591 <= not w9589 and not w9590;
w9592 <= not w9160 and not w9172;
w9593 <= not w9171 and not w9172;
w9594 <= not w9592 and not w9593;
w9595 <= not w2323 and w7036;
w9596 <= not w2468 and w6337;
w9597 <= not w2399 and w6886;
w9598 <= not w9596 and not w9597;
w9599 <= not w9595 and w9598;
w9600 <= not w6332 and w9599;
w9601 <= not w6526 and w9599;
w9602 <= not w9600 and not w9601;
w9603 <= a(14) and not w9602;
w9604 <= not a(14) and w9602;
w9605 <= not w9603 and not w9604;
w9606 <= not w9594 and not w9605;
w9607 <= not w2399 and w7036;
w9608 <= not w2506 and w6337;
w9609 <= not w2468 and w6886;
w9610 <= not w9608 and not w9609;
w9611 <= not w9607 and w9610;
w9612 <= w6332 and w6581;
w9613 <= w9611 and not w9612;
w9614 <= a(14) and not w9613;
w9615 <= not w9613 and not w9614;
w9616 <= a(14) and not w9614;
w9617 <= not w9615 and not w9616;
w9618 <= not w9144 and w9155;
w9619 <= not w9156 and not w9618;
w9620 <= not w9617 and w9619;
w9621 <= not w9617 and not w9620;
w9622 <= w9619 and not w9620;
w9623 <= not w9621 and not w9622;
w9624 <= w9141 and not w9143;
w9625 <= not w9144 and not w9624;
w9626 <= not w2468 and w7036;
w9627 <= not w2609 and w6337;
w9628 <= not w2506 and w6886;
w9629 <= not w9627 and not w9628;
w9630 <= not w9626 and w9629;
w9631 <= not w6332 and w9630;
w9632 <= not w6630 and w9630;
w9633 <= not w9631 and not w9632;
w9634 <= a(14) and not w9633;
w9635 <= not a(14) and w9633;
w9636 <= not w9634 and not w9635;
w9637 <= w9625 and not w9636;
w9638 <= not w2764 and w6886;
w9639 <= not w2671 and w7036;
w9640 <= not w9638 and not w9639;
w9641 <= w6332 and not w7404;
w9642 <= w9640 and not w9641;
w9643 <= a(14) and not w9642;
w9644 <= a(14) and not w9643;
w9645 <= not w9642 and not w9643;
w9646 <= not w9644 and not w9645;
w9647 <= not w2764 and not w6328;
w9648 <= a(14) and not w9647;
w9649 <= not w9646 and w9648;
w9650 <= not w2609 and w7036;
w9651 <= not w2764 and w6337;
w9652 <= not w2671 and w6886;
w9653 <= not w9651 and not w9652;
w9654 <= not w9650 and w9653;
w9655 <= not w6332 and w9654;
w9656 <= not w6733 and w9654;
w9657 <= not w9655 and not w9656;
w9658 <= a(14) and not w9657;
w9659 <= not a(14) and w9657;
w9660 <= not w9658 and not w9659;
w9661 <= w9649 and not w9660;
w9662 <= w9142 and w9661;
w9663 <= w9661 and not w9662;
w9664 <= w9142 and not w9662;
w9665 <= not w9663 and not w9664;
w9666 <= not w2506 and w7036;
w9667 <= not w2671 and w6337;
w9668 <= not w2609 and w6886;
w9669 <= not w9667 and not w9668;
w9670 <= not w9666 and w9669;
w9671 <= w6332 and w6741;
w9672 <= w9670 and not w9671;
w9673 <= a(14) and not w9672;
w9674 <= a(14) and not w9673;
w9675 <= not w9672 and not w9673;
w9676 <= not w9674 and not w9675;
w9677 <= not w9665 and not w9676;
w9678 <= not w9662 and not w9677;
w9679 <= not w9625 and w9636;
w9680 <= not w9637 and not w9679;
w9681 <= not w9678 and w9680;
w9682 <= not w9637 and not w9681;
w9683 <= not w9623 and not w9682;
w9684 <= not w9620 and not w9683;
w9685 <= w9594 and w9605;
w9686 <= not w9606 and not w9685;
w9687 <= not w9684 and w9686;
w9688 <= not w9606 and not w9687;
w9689 <= not w9591 and not w9688;
w9690 <= not w9588 and not w9689;
w9691 <= w9562 and not w9574;
w9692 <= not w9573 and not w9574;
w9693 <= not w9691 and not w9692;
w9694 <= not w9690 and not w9693;
w9695 <= not w9574 and not w9694;
w9696 <= w9548 and not w9560;
w9697 <= not w9559 and not w9560;
w9698 <= not w9696 and not w9697;
w9699 <= not w9695 and not w9698;
w9700 <= not w9560 and not w9699;
w9701 <= not w9534 and w9545;
w9702 <= not w9546 and not w9701;
w9703 <= not w9700 and w9702;
w9704 <= not w9546 and not w9703;
w9705 <= not w9532 and not w9704;
w9706 <= not w9529 and not w9705;
w9707 <= not w9514 and not w9706;
w9708 <= not w9511 and not w9707;
w9709 <= not w9496 and not w9708;
w9710 <= not w9493 and not w9709;
w9711 <= w9467 and not w9479;
w9712 <= not w9478 and not w9479;
w9713 <= not w9711 and not w9712;
w9714 <= not w9710 and not w9713;
w9715 <= not w9479 and not w9714;
w9716 <= w9453 and not w9465;
w9717 <= not w9464 and not w9465;
w9718 <= not w9716 and not w9717;
w9719 <= not w9715 and not w9718;
w9720 <= not w9465 and not w9719;
w9721 <= not w9439 and w9450;
w9722 <= not w9451 and not w9721;
w9723 <= not w9720 and w9722;
w9724 <= not w9451 and not w9723;
w9725 <= not w9437 and not w9724;
w9726 <= not w9434 and not w9725;
w9727 <= not w9419 and not w9726;
w9728 <= not w9416 and not w9727;
w9729 <= w9390 and not w9402;
w9730 <= not w9401 and not w9402;
w9731 <= not w9729 and not w9730;
w9732 <= not w9728 and not w9731;
w9733 <= not w9402 and not w9732;
w9734 <= w9376 and not w9388;
w9735 <= not w9387 and not w9388;
w9736 <= not w9734 and not w9735;
w9737 <= not w9733 and not w9736;
w9738 <= not w9388 and not w9737;
w9739 <= w9362 and not w9374;
w9740 <= not w9373 and not w9374;
w9741 <= not w9739 and not w9740;
w9742 <= not w9738 and not w9741;
w9743 <= not w9374 and not w9742;
w9744 <= w9348 and not w9360;
w9745 <= not w9359 and not w9360;
w9746 <= not w9744 and not w9745;
w9747 <= not w9743 and not w9746;
w9748 <= not w9360 and not w9747;
w9749 <= w9334 and not w9346;
w9750 <= not w9345 and not w9346;
w9751 <= not w9749 and not w9750;
w9752 <= not w9748 and not w9751;
w9753 <= not w9346 and not w9752;
w9754 <= w9320 and not w9332;
w9755 <= not w9331 and not w9332;
w9756 <= not w9754 and not w9755;
w9757 <= not w9753 and not w9756;
w9758 <= not w9332 and not w9757;
w9759 <= w9306 and not w9318;
w9760 <= not w9317 and not w9318;
w9761 <= not w9759 and not w9760;
w9762 <= not w9758 and not w9761;
w9763 <= not w9318 and not w9762;
w9764 <= w9242 and not w9244;
w9765 <= not w9245 and not w9764;
w9766 <= not w9763 and w9765;
w9767 <= not w3540 and w7918;
w9768 <= not w2947 and w7226;
w9769 <= not w3474 and w7567;
w9770 <= not w9768 and not w9769;
w9771 <= not w9767 and w9770;
w9772 <= w4019 and w7229;
w9773 <= w9771 and not w9772;
w9774 <= a(11) and not w9773;
w9775 <= not w9773 and not w9774;
w9776 <= a(11) and not w9774;
w9777 <= not w9775 and not w9776;
w9778 <= w9763 and not w9765;
w9779 <= not w9766 and not w9778;
w9780 <= not w9777 and w9779;
w9781 <= not w9766 and not w9780;
w9782 <= not w9304 and not w9781;
w9783 <= w9304 and w9781;
w9784 <= not w9782 and not w9783;
w9785 <= not w3980 and w9266;
w9786 <= not w3740 and w8353;
w9787 <= not w3899 and w8795;
w9788 <= not w9786 and not w9787;
w9789 <= not w9785 and w9788;
w9790 <= w4412 and w8356;
w9791 <= w9789 and not w9790;
w9792 <= a(8) and not w9791;
w9793 <= a(8) and not w9792;
w9794 <= not w9791 and not w9792;
w9795 <= not w9793 and not w9794;
w9796 <= w9784 and not w9795;
w9797 <= not w9782 and not w9796;
w9798 <= not a(3) and a(4);
w9799 <= a(3) and not a(4);
w9800 <= not w9798 and not w9799;
w9801 <= not w2 and w5;
w9802 <= w9800 and w9801;
w9803 <= not w4450 and w9802;
w9804 <= not w4457 and not w9803;
w9805 <= not w2 and not w5;
w9806 <= not w9803 and not w9805;
w9807 <= not w9804 and not w9806;
w9808 <= a(5) and not w9807;
w9809 <= not a(5) and w9807;
w9810 <= not w9808 and not w9809;
w9811 <= not w9797 and not w9810;
w9812 <= w9265 and not w9278;
w9813 <= not w9277 and not w9278;
w9814 <= not w9812 and not w9813;
w9815 <= w9797 and w9810;
w9816 <= not w9811 and not w9815;
w9817 <= not w9814 and w9816;
w9818 <= not w9811 and not w9817;
w9819 <= not w9293 and not w9296;
w9820 <= not w9292 and w9819;
w9821 <= not w9297 and not w9820;
w9822 <= not w9818 and w9821;
w9823 <= not w9814 and not w9817;
w9824 <= w9816 and not w9817;
w9825 <= not w9823 and not w9824;
w9826 <= not w3474 and w7918;
w9827 <= not w327 and w7226;
w9828 <= not w2947 and w7567;
w9829 <= not w9827 and not w9828;
w9830 <= not w9826 and w9829;
w9831 <= w3650 and w7229;
w9832 <= w9830 and not w9831;
w9833 <= a(11) and not w9832;
w9834 <= not w9832 and not w9833;
w9835 <= a(11) and not w9833;
w9836 <= not w9834 and not w9835;
w9837 <= not w9758 and not w9762;
w9838 <= not w9761 and not w9762;
w9839 <= not w9837 and not w9838;
w9840 <= not w9836 and not w9839;
w9841 <= not w9836 and not w9840;
w9842 <= not w9839 and not w9840;
w9843 <= not w9841 and not w9842;
w9844 <= not w2947 and w7918;
w9845 <= not w522 and w7226;
w9846 <= not w327 and w7567;
w9847 <= not w9845 and not w9846;
w9848 <= not w9844 and w9847;
w9849 <= w2953 and w7229;
w9850 <= w9848 and not w9849;
w9851 <= a(11) and not w9850;
w9852 <= not w9850 and not w9851;
w9853 <= a(11) and not w9851;
w9854 <= not w9852 and not w9853;
w9855 <= not w9753 and not w9757;
w9856 <= not w9756 and not w9757;
w9857 <= not w9855 and not w9856;
w9858 <= not w9854 and not w9857;
w9859 <= not w9854 and not w9858;
w9860 <= not w9857 and not w9858;
w9861 <= not w9859 and not w9860;
w9862 <= not w327 and w7918;
w9863 <= not w645 and w7226;
w9864 <= not w522 and w7567;
w9865 <= not w9863 and not w9864;
w9866 <= not w9862 and w9865;
w9867 <= w3282 and w7229;
w9868 <= w9866 and not w9867;
w9869 <= a(11) and not w9868;
w9870 <= not w9868 and not w9869;
w9871 <= a(11) and not w9869;
w9872 <= not w9870 and not w9871;
w9873 <= not w9748 and not w9752;
w9874 <= not w9751 and not w9752;
w9875 <= not w9873 and not w9874;
w9876 <= not w9872 and not w9875;
w9877 <= not w9872 and not w9876;
w9878 <= not w9875 and not w9876;
w9879 <= not w9877 and not w9878;
w9880 <= not w522 and w7918;
w9881 <= not w802 and w7226;
w9882 <= not w645 and w7567;
w9883 <= not w9881 and not w9882;
w9884 <= not w9880 and w9883;
w9885 <= w3266 and w7229;
w9886 <= w9884 and not w9885;
w9887 <= a(11) and not w9886;
w9888 <= not w9886 and not w9887;
w9889 <= a(11) and not w9887;
w9890 <= not w9888 and not w9889;
w9891 <= not w9743 and not w9747;
w9892 <= not w9746 and not w9747;
w9893 <= not w9891 and not w9892;
w9894 <= not w9890 and not w9893;
w9895 <= not w9890 and not w9894;
w9896 <= not w9893 and not w9894;
w9897 <= not w9895 and not w9896;
w9898 <= not w645 and w7918;
w9899 <= not w893 and w7226;
w9900 <= not w802 and w7567;
w9901 <= not w9899 and not w9900;
w9902 <= not w9898 and w9901;
w9903 <= w4114 and w7229;
w9904 <= w9902 and not w9903;
w9905 <= a(11) and not w9904;
w9906 <= not w9904 and not w9905;
w9907 <= a(11) and not w9905;
w9908 <= not w9906 and not w9907;
w9909 <= not w9738 and not w9742;
w9910 <= not w9741 and not w9742;
w9911 <= not w9909 and not w9910;
w9912 <= not w9908 and not w9911;
w9913 <= not w9908 and not w9912;
w9914 <= not w9911 and not w9912;
w9915 <= not w9913 and not w9914;
w9916 <= not w802 and w7918;
w9917 <= not w995 and w7226;
w9918 <= not w893 and w7567;
w9919 <= not w9917 and not w9918;
w9920 <= not w9916 and w9919;
w9921 <= w4139 and w7229;
w9922 <= w9920 and not w9921;
w9923 <= a(11) and not w9922;
w9924 <= not w9922 and not w9923;
w9925 <= a(11) and not w9923;
w9926 <= not w9924 and not w9925;
w9927 <= not w9733 and not w9737;
w9928 <= not w9736 and not w9737;
w9929 <= not w9927 and not w9928;
w9930 <= not w9926 and not w9929;
w9931 <= not w9926 and not w9930;
w9932 <= not w9929 and not w9930;
w9933 <= not w9931 and not w9932;
w9934 <= not w893 and w7918;
w9935 <= not w1113 and w7226;
w9936 <= not w995 and w7567;
w9937 <= not w9935 and not w9936;
w9938 <= not w9934 and w9937;
w9939 <= w4568 and w7229;
w9940 <= w9938 and not w9939;
w9941 <= a(11) and not w9940;
w9942 <= not w9940 and not w9941;
w9943 <= a(11) and not w9941;
w9944 <= not w9942 and not w9943;
w9945 <= not w9728 and not w9732;
w9946 <= not w9731 and not w9732;
w9947 <= not w9945 and not w9946;
w9948 <= not w9944 and not w9947;
w9949 <= not w9944 and not w9948;
w9950 <= not w9947 and not w9948;
w9951 <= not w9949 and not w9950;
w9952 <= w9419 and w9726;
w9953 <= not w9727 and not w9952;
w9954 <= not w995 and w7918;
w9955 <= not w1170 and w7226;
w9956 <= not w1113 and w7567;
w9957 <= not w9955 and not w9956;
w9958 <= not w9954 and w9957;
w9959 <= not w7229 and w9958;
w9960 <= not w4364 and w9958;
w9961 <= not w9959 and not w9960;
w9962 <= a(11) and not w9961;
w9963 <= not a(11) and w9961;
w9964 <= not w9962 and not w9963;
w9965 <= w9953 and not w9964;
w9966 <= w9437 and w9724;
w9967 <= not w9725 and not w9966;
w9968 <= not w1113 and w7918;
w9969 <= not w1299 and w7226;
w9970 <= not w1170 and w7567;
w9971 <= not w9969 and not w9970;
w9972 <= not w9968 and w9971;
w9973 <= not w7229 and w9972;
w9974 <= not w4796 and w9972;
w9975 <= not w9973 and not w9974;
w9976 <= a(11) and not w9975;
w9977 <= not a(11) and w9975;
w9978 <= not w9976 and not w9977;
w9979 <= w9967 and not w9978;
w9980 <= not w1170 and w7918;
w9981 <= not w1407 and w7226;
w9982 <= not w1299 and w7567;
w9983 <= not w9981 and not w9982;
w9984 <= not w9980 and w9983;
w9985 <= w4783 and w7229;
w9986 <= w9984 and not w9985;
w9987 <= a(11) and not w9986;
w9988 <= not w9986 and not w9987;
w9989 <= a(11) and not w9987;
w9990 <= not w9988 and not w9989;
w9991 <= w9720 and not w9722;
w9992 <= not w9723 and not w9991;
w9993 <= not w9990 and w9992;
w9994 <= not w9990 and not w9993;
w9995 <= w9992 and not w9993;
w9996 <= not w9994 and not w9995;
w9997 <= not w1299 and w7918;
w9998 <= not w1507 and w7226;
w9999 <= not w1407 and w7567;
w10000 <= not w9998 and not w9999;
w10001 <= not w9997 and w10000;
w10002 <= w5049 and w7229;
w10003 <= w10001 and not w10002;
w10004 <= a(11) and not w10003;
w10005 <= not w10003 and not w10004;
w10006 <= a(11) and not w10004;
w10007 <= not w10005 and not w10006;
w10008 <= not w9715 and not w9719;
w10009 <= not w9718 and not w9719;
w10010 <= not w10008 and not w10009;
w10011 <= not w10007 and not w10010;
w10012 <= not w10007 and not w10011;
w10013 <= not w10010 and not w10011;
w10014 <= not w10012 and not w10013;
w10015 <= not w1407 and w7918;
w10016 <= not w1600 and w7226;
w10017 <= not w1507 and w7567;
w10018 <= not w10016 and not w10017;
w10019 <= not w10015 and w10018;
w10020 <= w5074 and w7229;
w10021 <= w10019 and not w10020;
w10022 <= a(11) and not w10021;
w10023 <= not w10021 and not w10022;
w10024 <= a(11) and not w10022;
w10025 <= not w10023 and not w10024;
w10026 <= not w9710 and not w9714;
w10027 <= not w9713 and not w9714;
w10028 <= not w10026 and not w10027;
w10029 <= not w10025 and not w10028;
w10030 <= not w10025 and not w10029;
w10031 <= not w10028 and not w10029;
w10032 <= not w10030 and not w10031;
w10033 <= w9496 and w9708;
w10034 <= not w9709 and not w10033;
w10035 <= not w1507 and w7918;
w10036 <= not w1714 and w7226;
w10037 <= not w1600 and w7567;
w10038 <= not w10036 and not w10037;
w10039 <= not w10035 and w10038;
w10040 <= not w7229 and w10039;
w10041 <= not w5496 and w10039;
w10042 <= not w10040 and not w10041;
w10043 <= a(11) and not w10042;
w10044 <= not a(11) and w10042;
w10045 <= not w10043 and not w10044;
w10046 <= w10034 and not w10045;
w10047 <= w9514 and w9706;
w10048 <= not w9707 and not w10047;
w10049 <= not w1600 and w7918;
w10050 <= not w1812 and w7226;
w10051 <= not w1714 and w7567;
w10052 <= not w10050 and not w10051;
w10053 <= not w10049 and w10052;
w10054 <= not w7229 and w10053;
w10055 <= not w5263 and w10053;
w10056 <= not w10054 and not w10055;
w10057 <= a(11) and not w10056;
w10058 <= not a(11) and w10056;
w10059 <= not w10057 and not w10058;
w10060 <= w10048 and not w10059;
w10061 <= w9532 and w9704;
w10062 <= not w9705 and not w10061;
w10063 <= not w1714 and w7918;
w10064 <= not w1848 and w7226;
w10065 <= not w1812 and w7567;
w10066 <= not w10064 and not w10065;
w10067 <= not w10063 and w10066;
w10068 <= not w7229 and w10067;
w10069 <= not w5786 and w10067;
w10070 <= not w10068 and not w10069;
w10071 <= a(11) and not w10070;
w10072 <= not a(11) and w10070;
w10073 <= not w10071 and not w10072;
w10074 <= w10062 and not w10073;
w10075 <= not w1812 and w7918;
w10076 <= not w1927 and w7226;
w10077 <= not w1848 and w7567;
w10078 <= not w10076 and not w10077;
w10079 <= not w10075 and w10078;
w10080 <= w5942 and w7229;
w10081 <= w10079 and not w10080;
w10082 <= a(11) and not w10081;
w10083 <= not w10081 and not w10082;
w10084 <= a(11) and not w10082;
w10085 <= not w10083 and not w10084;
w10086 <= w9700 and not w9702;
w10087 <= not w9703 and not w10086;
w10088 <= not w10085 and w10087;
w10089 <= not w10085 and not w10088;
w10090 <= w10087 and not w10088;
w10091 <= not w10089 and not w10090;
w10092 <= not w1848 and w7918;
w10093 <= not w1992 and w7226;
w10094 <= not w1927 and w7567;
w10095 <= not w10093 and not w10094;
w10096 <= not w10092 and w10095;
w10097 <= w5769 and w7229;
w10098 <= w10096 and not w10097;
w10099 <= a(11) and not w10098;
w10100 <= not w10098 and not w10099;
w10101 <= a(11) and not w10099;
w10102 <= not w10100 and not w10101;
w10103 <= not w9695 and not w9699;
w10104 <= not w9698 and not w9699;
w10105 <= not w10103 and not w10104;
w10106 <= not w10102 and not w10105;
w10107 <= not w10102 and not w10106;
w10108 <= not w10105 and not w10106;
w10109 <= not w10107 and not w10108;
w10110 <= not w1927 and w7918;
w10111 <= not w2087 and w7226;
w10112 <= not w1992 and w7567;
w10113 <= not w10111 and not w10112;
w10114 <= not w10110 and w10113;
w10115 <= w6078 and w7229;
w10116 <= w10114 and not w10115;
w10117 <= a(11) and not w10116;
w10118 <= not w10116 and not w10117;
w10119 <= a(11) and not w10117;
w10120 <= not w10118 and not w10119;
w10121 <= not w9690 and not w9694;
w10122 <= not w9693 and not w9694;
w10123 <= not w10121 and not w10122;
w10124 <= not w10120 and not w10123;
w10125 <= not w10120 and not w10124;
w10126 <= not w10123 and not w10124;
w10127 <= not w10125 and not w10126;
w10128 <= w9591 and w9688;
w10129 <= not w9689 and not w10128;
w10130 <= not w1992 and w7918;
w10131 <= not w2124 and w7226;
w10132 <= not w2087 and w7567;
w10133 <= not w10131 and not w10132;
w10134 <= not w10130 and w10133;
w10135 <= not w7229 and w10134;
w10136 <= not w6414 and w10134;
w10137 <= not w10135 and not w10136;
w10138 <= a(11) and not w10137;
w10139 <= not a(11) and w10137;
w10140 <= not w10138 and not w10139;
w10141 <= w10129 and not w10140;
w10142 <= w9684 and not w9686;
w10143 <= not w9687 and not w10142;
w10144 <= not w2087 and w7918;
w10145 <= not w2226 and w7226;
w10146 <= not w2124 and w7567;
w10147 <= not w10145 and not w10146;
w10148 <= not w10144 and w10147;
w10149 <= not w7229 and w10148;
w10150 <= not w6427 and w10148;
w10151 <= not w10149 and not w10150;
w10152 <= a(11) and not w10151;
w10153 <= not a(11) and w10151;
w10154 <= not w10152 and not w10153;
w10155 <= w10143 and not w10154;
w10156 <= w9623 and w9682;
w10157 <= not w9683 and not w10156;
w10158 <= not w2124 and w7918;
w10159 <= not w2323 and w7226;
w10160 <= not w2226 and w7567;
w10161 <= not w10159 and not w10160;
w10162 <= not w10158 and w10161;
w10163 <= not w7229 and w10162;
w10164 <= not w6057 and w10162;
w10165 <= not w10163 and not w10164;
w10166 <= a(11) and not w10165;
w10167 <= not a(11) and w10165;
w10168 <= not w10166 and not w10167;
w10169 <= w10157 and not w10168;
w10170 <= not w2226 and w7918;
w10171 <= not w2399 and w7226;
w10172 <= not w2323 and w7567;
w10173 <= not w10171 and not w10172;
w10174 <= not w10170 and w10173;
w10175 <= w6476 and w7229;
w10176 <= w10174 and not w10175;
w10177 <= a(11) and not w10176;
w10178 <= not w10176 and not w10177;
w10179 <= a(11) and not w10177;
w10180 <= not w10178 and not w10179;
w10181 <= w9678 and not w9680;
w10182 <= not w9681 and not w10181;
w10183 <= not w10180 and w10182;
w10184 <= not w10180 and not w10183;
w10185 <= w10182 and not w10183;
w10186 <= not w10184 and not w10185;
w10187 <= not w9665 and not w9677;
w10188 <= not w9676 and not w9677;
w10189 <= not w10187 and not w10188;
w10190 <= not w2323 and w7918;
w10191 <= not w2468 and w7226;
w10192 <= not w2399 and w7567;
w10193 <= not w10191 and not w10192;
w10194 <= not w10190 and w10193;
w10195 <= not w7229 and w10194;
w10196 <= not w6526 and w10194;
w10197 <= not w10195 and not w10196;
w10198 <= a(11) and not w10197;
w10199 <= not a(11) and w10197;
w10200 <= not w10198 and not w10199;
w10201 <= not w10189 and not w10200;
w10202 <= not w2399 and w7918;
w10203 <= not w2506 and w7226;
w10204 <= not w2468 and w7567;
w10205 <= not w10203 and not w10204;
w10206 <= not w10202 and w10205;
w10207 <= w6581 and w7229;
w10208 <= w10206 and not w10207;
w10209 <= a(11) and not w10208;
w10210 <= not w10208 and not w10209;
w10211 <= a(11) and not w10209;
w10212 <= not w10210 and not w10211;
w10213 <= not w9649 and w9660;
w10214 <= not w9661 and not w10213;
w10215 <= not w10212 and w10214;
w10216 <= not w10212 and not w10215;
w10217 <= w10214 and not w10215;
w10218 <= not w10216 and not w10217;
w10219 <= w9646 and not w9648;
w10220 <= not w9649 and not w10219;
w10221 <= not w2468 and w7918;
w10222 <= not w2609 and w7226;
w10223 <= not w2506 and w7567;
w10224 <= not w10222 and not w10223;
w10225 <= not w10221 and w10224;
w10226 <= not w7229 and w10225;
w10227 <= not w6630 and w10225;
w10228 <= not w10226 and not w10227;
w10229 <= a(11) and not w10228;
w10230 <= not a(11) and w10228;
w10231 <= not w10229 and not w10230;
w10232 <= w10220 and not w10231;
w10233 <= not w2764 and w7567;
w10234 <= not w2671 and w7918;
w10235 <= not w10233 and not w10234;
w10236 <= w7229 and not w7404;
w10237 <= w10235 and not w10236;
w10238 <= a(11) and not w10237;
w10239 <= a(11) and not w10238;
w10240 <= not w10237 and not w10238;
w10241 <= not w10239 and not w10240;
w10242 <= not w2764 and not w7224;
w10243 <= a(11) and not w10242;
w10244 <= not w10241 and w10243;
w10245 <= not w2609 and w7918;
w10246 <= not w2764 and w7226;
w10247 <= not w2671 and w7567;
w10248 <= not w10246 and not w10247;
w10249 <= not w10245 and w10248;
w10250 <= not w7229 and w10249;
w10251 <= not w6733 and w10249;
w10252 <= not w10250 and not w10251;
w10253 <= a(11) and not w10252;
w10254 <= not a(11) and w10252;
w10255 <= not w10253 and not w10254;
w10256 <= w10244 and not w10255;
w10257 <= w9647 and w10256;
w10258 <= w10256 and not w10257;
w10259 <= w9647 and not w10257;
w10260 <= not w10258 and not w10259;
w10261 <= not w2506 and w7918;
w10262 <= not w2671 and w7226;
w10263 <= not w2609 and w7567;
w10264 <= not w10262 and not w10263;
w10265 <= not w10261 and w10264;
w10266 <= w6741 and w7229;
w10267 <= w10265 and not w10266;
w10268 <= a(11) and not w10267;
w10269 <= a(11) and not w10268;
w10270 <= not w10267 and not w10268;
w10271 <= not w10269 and not w10270;
w10272 <= not w10260 and not w10271;
w10273 <= not w10257 and not w10272;
w10274 <= not w10220 and w10231;
w10275 <= not w10232 and not w10274;
w10276 <= not w10273 and w10275;
w10277 <= not w10232 and not w10276;
w10278 <= not w10218 and not w10277;
w10279 <= not w10215 and not w10278;
w10280 <= w10189 and w10200;
w10281 <= not w10201 and not w10280;
w10282 <= not w10279 and w10281;
w10283 <= not w10201 and not w10282;
w10284 <= not w10186 and not w10283;
w10285 <= not w10183 and not w10284;
w10286 <= w10157 and not w10169;
w10287 <= not w10168 and not w10169;
w10288 <= not w10286 and not w10287;
w10289 <= not w10285 and not w10288;
w10290 <= not w10169 and not w10289;
w10291 <= w10143 and not w10155;
w10292 <= not w10154 and not w10155;
w10293 <= not w10291 and not w10292;
w10294 <= not w10290 and not w10293;
w10295 <= not w10155 and not w10294;
w10296 <= not w10129 and w10140;
w10297 <= not w10141 and not w10296;
w10298 <= not w10295 and w10297;
w10299 <= not w10141 and not w10298;
w10300 <= not w10127 and not w10299;
w10301 <= not w10124 and not w10300;
w10302 <= not w10109 and not w10301;
w10303 <= not w10106 and not w10302;
w10304 <= not w10091 and not w10303;
w10305 <= not w10088 and not w10304;
w10306 <= w10062 and not w10074;
w10307 <= not w10073 and not w10074;
w10308 <= not w10306 and not w10307;
w10309 <= not w10305 and not w10308;
w10310 <= not w10074 and not w10309;
w10311 <= w10048 and not w10060;
w10312 <= not w10059 and not w10060;
w10313 <= not w10311 and not w10312;
w10314 <= not w10310 and not w10313;
w10315 <= not w10060 and not w10314;
w10316 <= not w10034 and w10045;
w10317 <= not w10046 and not w10316;
w10318 <= not w10315 and w10317;
w10319 <= not w10046 and not w10318;
w10320 <= not w10032 and not w10319;
w10321 <= not w10029 and not w10320;
w10322 <= not w10014 and not w10321;
w10323 <= not w10011 and not w10322;
w10324 <= not w9996 and not w10323;
w10325 <= not w9993 and not w10324;
w10326 <= w9967 and not w9979;
w10327 <= not w9978 and not w9979;
w10328 <= not w10326 and not w10327;
w10329 <= not w10325 and not w10328;
w10330 <= not w9979 and not w10329;
w10331 <= not w9953 and w9964;
w10332 <= not w9965 and not w10331;
w10333 <= not w10330 and w10332;
w10334 <= not w9965 and not w10333;
w10335 <= not w9951 and not w10334;
w10336 <= not w9948 and not w10335;
w10337 <= not w9933 and not w10336;
w10338 <= not w9930 and not w10337;
w10339 <= not w9915 and not w10338;
w10340 <= not w9912 and not w10339;
w10341 <= not w9897 and not w10340;
w10342 <= not w9894 and not w10341;
w10343 <= not w9879 and not w10342;
w10344 <= not w9876 and not w10343;
w10345 <= not w9861 and not w10344;
w10346 <= not w9858 and not w10345;
w10347 <= not w9843 and not w10346;
w10348 <= not w9840 and not w10347;
w10349 <= w9777 and not w9779;
w10350 <= not w9780 and not w10349;
w10351 <= not w10348 and w10350;
w10352 <= not w3899 and w9266;
w10353 <= not w3391 and w8353;
w10354 <= not w3740 and w8795;
w10355 <= not w10353 and not w10354;
w10356 <= not w10352 and w10355;
w10357 <= w4493 and w8356;
w10358 <= w10356 and not w10357;
w10359 <= a(8) and not w10358;
w10360 <= not w10358 and not w10359;
w10361 <= a(8) and not w10359;
w10362 <= not w10360 and not w10361;
w10363 <= not w10348 and not w10351;
w10364 <= w10350 and not w10351;
w10365 <= not w10363 and not w10364;
w10366 <= not w10362 and not w10365;
w10367 <= not w10351 and not w10366;
w10368 <= not w3812 and w9802;
w10369 <= w5 and not w9800;
w10370 <= not w4450 and w10369;
w10371 <= not w10368 and not w10370;
w10372 <= not w9805 and w10371;
w10373 <= not w4544 and w10371;
w10374 <= not w10372 and not w10373;
w10375 <= a(5) and not w10374;
w10376 <= not a(5) and w10374;
w10377 <= not w10375 and not w10376;
w10378 <= not w10367 and not w10377;
w10379 <= w9784 and not w9796;
w10380 <= not w9795 and not w9796;
w10381 <= not w10379 and not w10380;
w10382 <= w10367 and w10377;
w10383 <= not w10378 and not w10382;
w10384 <= not w10381 and w10383;
w10385 <= not w10378 and not w10384;
w10386 <= not w9825 and not w10385;
w10387 <= w9825 and w10385;
w10388 <= not w10386 and not w10387;
w10389 <= w9843 and w10346;
w10390 <= not w10347 and not w10389;
w10391 <= not w3740 and w9266;
w10392 <= not w3540 and w8353;
w10393 <= not w3391 and w8795;
w10394 <= not w10392 and not w10393;
w10395 <= not w10391 and w10394;
w10396 <= not w8356 and w10395;
w10397 <= not w3753 and w10395;
w10398 <= not w10396 and not w10397;
w10399 <= a(8) and not w10398;
w10400 <= not a(8) and w10398;
w10401 <= not w10399 and not w10400;
w10402 <= w10390 and not w10401;
w10403 <= w9861 and w10344;
w10404 <= not w10345 and not w10403;
w10405 <= not w3391 and w9266;
w10406 <= not w3474 and w8353;
w10407 <= not w3540 and w8795;
w10408 <= not w10406 and not w10407;
w10409 <= not w10405 and w10408;
w10410 <= not w8356 and w10409;
w10411 <= not w3562 and w10409;
w10412 <= not w10410 and not w10411;
w10413 <= a(8) and not w10412;
w10414 <= not a(8) and w10412;
w10415 <= not w10413 and not w10414;
w10416 <= w10404 and not w10415;
w10417 <= w9879 and w10342;
w10418 <= not w10343 and not w10417;
w10419 <= not w3540 and w9266;
w10420 <= not w2947 and w8353;
w10421 <= not w3474 and w8795;
w10422 <= not w10420 and not w10421;
w10423 <= not w10419 and w10422;
w10424 <= not w8356 and w10423;
w10425 <= not w4019 and w10423;
w10426 <= not w10424 and not w10425;
w10427 <= a(8) and not w10426;
w10428 <= not a(8) and w10426;
w10429 <= not w10427 and not w10428;
w10430 <= w10418 and not w10429;
w10431 <= w9897 and w10340;
w10432 <= not w10341 and not w10431;
w10433 <= not w3474 and w9266;
w10434 <= not w327 and w8353;
w10435 <= not w2947 and w8795;
w10436 <= not w10434 and not w10435;
w10437 <= not w10433 and w10436;
w10438 <= not w8356 and w10437;
w10439 <= not w3650 and w10437;
w10440 <= not w10438 and not w10439;
w10441 <= a(8) and not w10440;
w10442 <= not a(8) and w10440;
w10443 <= not w10441 and not w10442;
w10444 <= w10432 and not w10443;
w10445 <= w9915 and w10338;
w10446 <= not w10339 and not w10445;
w10447 <= not w2947 and w9266;
w10448 <= not w522 and w8353;
w10449 <= not w327 and w8795;
w10450 <= not w10448 and not w10449;
w10451 <= not w10447 and w10450;
w10452 <= not w8356 and w10451;
w10453 <= not w2953 and w10451;
w10454 <= not w10452 and not w10453;
w10455 <= a(8) and not w10454;
w10456 <= not a(8) and w10454;
w10457 <= not w10455 and not w10456;
w10458 <= w10446 and not w10457;
w10459 <= w9933 and w10336;
w10460 <= not w10337 and not w10459;
w10461 <= not w327 and w9266;
w10462 <= not w645 and w8353;
w10463 <= not w522 and w8795;
w10464 <= not w10462 and not w10463;
w10465 <= not w10461 and w10464;
w10466 <= not w8356 and w10465;
w10467 <= not w3282 and w10465;
w10468 <= not w10466 and not w10467;
w10469 <= a(8) and not w10468;
w10470 <= not a(8) and w10468;
w10471 <= not w10469 and not w10470;
w10472 <= w10460 and not w10471;
w10473 <= w9951 and w10334;
w10474 <= not w10335 and not w10473;
w10475 <= not w522 and w9266;
w10476 <= not w802 and w8353;
w10477 <= not w645 and w8795;
w10478 <= not w10476 and not w10477;
w10479 <= not w10475 and w10478;
w10480 <= not w8356 and w10479;
w10481 <= not w3266 and w10479;
w10482 <= not w10480 and not w10481;
w10483 <= a(8) and not w10482;
w10484 <= not a(8) and w10482;
w10485 <= not w10483 and not w10484;
w10486 <= w10474 and not w10485;
w10487 <= not w645 and w9266;
w10488 <= not w893 and w8353;
w10489 <= not w802 and w8795;
w10490 <= not w10488 and not w10489;
w10491 <= not w10487 and w10490;
w10492 <= w4114 and w8356;
w10493 <= w10491 and not w10492;
w10494 <= a(8) and not w10493;
w10495 <= not w10493 and not w10494;
w10496 <= a(8) and not w10494;
w10497 <= not w10495 and not w10496;
w10498 <= w10330 and not w10332;
w10499 <= not w10333 and not w10498;
w10500 <= not w10497 and w10499;
w10501 <= not w10497 and not w10500;
w10502 <= w10499 and not w10500;
w10503 <= not w10501 and not w10502;
w10504 <= not w802 and w9266;
w10505 <= not w995 and w8353;
w10506 <= not w893 and w8795;
w10507 <= not w10505 and not w10506;
w10508 <= not w10504 and w10507;
w10509 <= w4139 and w8356;
w10510 <= w10508 and not w10509;
w10511 <= a(8) and not w10510;
w10512 <= not w10510 and not w10511;
w10513 <= a(8) and not w10511;
w10514 <= not w10512 and not w10513;
w10515 <= not w10325 and not w10329;
w10516 <= not w10328 and not w10329;
w10517 <= not w10515 and not w10516;
w10518 <= not w10514 and not w10517;
w10519 <= not w10514 and not w10518;
w10520 <= not w10517 and not w10518;
w10521 <= not w10519 and not w10520;
w10522 <= w9996 and w10323;
w10523 <= not w10324 and not w10522;
w10524 <= not w893 and w9266;
w10525 <= not w1113 and w8353;
w10526 <= not w995 and w8795;
w10527 <= not w10525 and not w10526;
w10528 <= not w10524 and w10527;
w10529 <= not w8356 and w10528;
w10530 <= not w4568 and w10528;
w10531 <= not w10529 and not w10530;
w10532 <= a(8) and not w10531;
w10533 <= not a(8) and w10531;
w10534 <= not w10532 and not w10533;
w10535 <= w10523 and not w10534;
w10536 <= w10014 and w10321;
w10537 <= not w10322 and not w10536;
w10538 <= not w995 and w9266;
w10539 <= not w1170 and w8353;
w10540 <= not w1113 and w8795;
w10541 <= not w10539 and not w10540;
w10542 <= not w10538 and w10541;
w10543 <= not w8356 and w10542;
w10544 <= not w4364 and w10542;
w10545 <= not w10543 and not w10544;
w10546 <= a(8) and not w10545;
w10547 <= not a(8) and w10545;
w10548 <= not w10546 and not w10547;
w10549 <= w10537 and not w10548;
w10550 <= w10032 and w10319;
w10551 <= not w10320 and not w10550;
w10552 <= not w1113 and w9266;
w10553 <= not w1299 and w8353;
w10554 <= not w1170 and w8795;
w10555 <= not w10553 and not w10554;
w10556 <= not w10552 and w10555;
w10557 <= not w8356 and w10556;
w10558 <= not w4796 and w10556;
w10559 <= not w10557 and not w10558;
w10560 <= a(8) and not w10559;
w10561 <= not a(8) and w10559;
w10562 <= not w10560 and not w10561;
w10563 <= w10551 and not w10562;
w10564 <= not w1170 and w9266;
w10565 <= not w1407 and w8353;
w10566 <= not w1299 and w8795;
w10567 <= not w10565 and not w10566;
w10568 <= not w10564 and w10567;
w10569 <= w4783 and w8356;
w10570 <= w10568 and not w10569;
w10571 <= a(8) and not w10570;
w10572 <= not w10570 and not w10571;
w10573 <= a(8) and not w10571;
w10574 <= not w10572 and not w10573;
w10575 <= w10315 and not w10317;
w10576 <= not w10318 and not w10575;
w10577 <= not w10574 and w10576;
w10578 <= not w10574 and not w10577;
w10579 <= w10576 and not w10577;
w10580 <= not w10578 and not w10579;
w10581 <= not w1299 and w9266;
w10582 <= not w1507 and w8353;
w10583 <= not w1407 and w8795;
w10584 <= not w10582 and not w10583;
w10585 <= not w10581 and w10584;
w10586 <= w5049 and w8356;
w10587 <= w10585 and not w10586;
w10588 <= a(8) and not w10587;
w10589 <= not w10587 and not w10588;
w10590 <= a(8) and not w10588;
w10591 <= not w10589 and not w10590;
w10592 <= not w10310 and not w10314;
w10593 <= not w10313 and not w10314;
w10594 <= not w10592 and not w10593;
w10595 <= not w10591 and not w10594;
w10596 <= not w10591 and not w10595;
w10597 <= not w10594 and not w10595;
w10598 <= not w10596 and not w10597;
w10599 <= not w1407 and w9266;
w10600 <= not w1600 and w8353;
w10601 <= not w1507 and w8795;
w10602 <= not w10600 and not w10601;
w10603 <= not w10599 and w10602;
w10604 <= w5074 and w8356;
w10605 <= w10603 and not w10604;
w10606 <= a(8) and not w10605;
w10607 <= not w10605 and not w10606;
w10608 <= a(8) and not w10606;
w10609 <= not w10607 and not w10608;
w10610 <= not w10305 and not w10309;
w10611 <= not w10308 and not w10309;
w10612 <= not w10610 and not w10611;
w10613 <= not w10609 and not w10612;
w10614 <= not w10609 and not w10613;
w10615 <= not w10612 and not w10613;
w10616 <= not w10614 and not w10615;
w10617 <= w10091 and w10303;
w10618 <= not w10304 and not w10617;
w10619 <= not w1507 and w9266;
w10620 <= not w1714 and w8353;
w10621 <= not w1600 and w8795;
w10622 <= not w10620 and not w10621;
w10623 <= not w10619 and w10622;
w10624 <= not w8356 and w10623;
w10625 <= not w5496 and w10623;
w10626 <= not w10624 and not w10625;
w10627 <= a(8) and not w10626;
w10628 <= not a(8) and w10626;
w10629 <= not w10627 and not w10628;
w10630 <= w10618 and not w10629;
w10631 <= w10109 and w10301;
w10632 <= not w10302 and not w10631;
w10633 <= not w1600 and w9266;
w10634 <= not w1812 and w8353;
w10635 <= not w1714 and w8795;
w10636 <= not w10634 and not w10635;
w10637 <= not w10633 and w10636;
w10638 <= not w8356 and w10637;
w10639 <= not w5263 and w10637;
w10640 <= not w10638 and not w10639;
w10641 <= a(8) and not w10640;
w10642 <= not a(8) and w10640;
w10643 <= not w10641 and not w10642;
w10644 <= w10632 and not w10643;
w10645 <= w10127 and w10299;
w10646 <= not w10300 and not w10645;
w10647 <= not w1714 and w9266;
w10648 <= not w1848 and w8353;
w10649 <= not w1812 and w8795;
w10650 <= not w10648 and not w10649;
w10651 <= not w10647 and w10650;
w10652 <= not w8356 and w10651;
w10653 <= not w5786 and w10651;
w10654 <= not w10652 and not w10653;
w10655 <= a(8) and not w10654;
w10656 <= not a(8) and w10654;
w10657 <= not w10655 and not w10656;
w10658 <= w10646 and not w10657;
w10659 <= not w1812 and w9266;
w10660 <= not w1927 and w8353;
w10661 <= not w1848 and w8795;
w10662 <= not w10660 and not w10661;
w10663 <= not w10659 and w10662;
w10664 <= w5942 and w8356;
w10665 <= w10663 and not w10664;
w10666 <= a(8) and not w10665;
w10667 <= not w10665 and not w10666;
w10668 <= a(8) and not w10666;
w10669 <= not w10667 and not w10668;
w10670 <= w10295 and not w10297;
w10671 <= not w10298 and not w10670;
w10672 <= not w10669 and w10671;
w10673 <= not w10669 and not w10672;
w10674 <= w10671 and not w10672;
w10675 <= not w10673 and not w10674;
w10676 <= not w1848 and w9266;
w10677 <= not w1992 and w8353;
w10678 <= not w1927 and w8795;
w10679 <= not w10677 and not w10678;
w10680 <= not w10676 and w10679;
w10681 <= w5769 and w8356;
w10682 <= w10680 and not w10681;
w10683 <= a(8) and not w10682;
w10684 <= not w10682 and not w10683;
w10685 <= a(8) and not w10683;
w10686 <= not w10684 and not w10685;
w10687 <= not w10290 and not w10294;
w10688 <= not w10293 and not w10294;
w10689 <= not w10687 and not w10688;
w10690 <= not w10686 and not w10689;
w10691 <= not w10686 and not w10690;
w10692 <= not w10689 and not w10690;
w10693 <= not w10691 and not w10692;
w10694 <= not w1927 and w9266;
w10695 <= not w2087 and w8353;
w10696 <= not w1992 and w8795;
w10697 <= not w10695 and not w10696;
w10698 <= not w10694 and w10697;
w10699 <= w6078 and w8356;
w10700 <= w10698 and not w10699;
w10701 <= a(8) and not w10700;
w10702 <= not w10700 and not w10701;
w10703 <= a(8) and not w10701;
w10704 <= not w10702 and not w10703;
w10705 <= not w10285 and not w10289;
w10706 <= not w10288 and not w10289;
w10707 <= not w10705 and not w10706;
w10708 <= not w10704 and not w10707;
w10709 <= not w10704 and not w10708;
w10710 <= not w10707 and not w10708;
w10711 <= not w10709 and not w10710;
w10712 <= w10186 and w10283;
w10713 <= not w10284 and not w10712;
w10714 <= not w1992 and w9266;
w10715 <= not w2124 and w8353;
w10716 <= not w2087 and w8795;
w10717 <= not w10715 and not w10716;
w10718 <= not w10714 and w10717;
w10719 <= not w8356 and w10718;
w10720 <= not w6414 and w10718;
w10721 <= not w10719 and not w10720;
w10722 <= a(8) and not w10721;
w10723 <= not a(8) and w10721;
w10724 <= not w10722 and not w10723;
w10725 <= w10713 and not w10724;
w10726 <= w10279 and not w10281;
w10727 <= not w10282 and not w10726;
w10728 <= not w2087 and w9266;
w10729 <= not w2226 and w8353;
w10730 <= not w2124 and w8795;
w10731 <= not w10729 and not w10730;
w10732 <= not w10728 and w10731;
w10733 <= not w8356 and w10732;
w10734 <= not w6427 and w10732;
w10735 <= not w10733 and not w10734;
w10736 <= a(8) and not w10735;
w10737 <= not a(8) and w10735;
w10738 <= not w10736 and not w10737;
w10739 <= w10727 and not w10738;
w10740 <= w10218 and w10277;
w10741 <= not w10278 and not w10740;
w10742 <= not w2124 and w9266;
w10743 <= not w2323 and w8353;
w10744 <= not w2226 and w8795;
w10745 <= not w10743 and not w10744;
w10746 <= not w10742 and w10745;
w10747 <= not w8356 and w10746;
w10748 <= not w6057 and w10746;
w10749 <= not w10747 and not w10748;
w10750 <= a(8) and not w10749;
w10751 <= not a(8) and w10749;
w10752 <= not w10750 and not w10751;
w10753 <= w10741 and not w10752;
w10754 <= not w2226 and w9266;
w10755 <= not w2399 and w8353;
w10756 <= not w2323 and w8795;
w10757 <= not w10755 and not w10756;
w10758 <= not w10754 and w10757;
w10759 <= w6476 and w8356;
w10760 <= w10758 and not w10759;
w10761 <= a(8) and not w10760;
w10762 <= not w10760 and not w10761;
w10763 <= a(8) and not w10761;
w10764 <= not w10762 and not w10763;
w10765 <= w10273 and not w10275;
w10766 <= not w10276 and not w10765;
w10767 <= not w10764 and w10766;
w10768 <= not w10764 and not w10767;
w10769 <= w10766 and not w10767;
w10770 <= not w10768 and not w10769;
w10771 <= not w10260 and not w10272;
w10772 <= not w10271 and not w10272;
w10773 <= not w10771 and not w10772;
w10774 <= not w2323 and w9266;
w10775 <= not w2468 and w8353;
w10776 <= not w2399 and w8795;
w10777 <= not w10775 and not w10776;
w10778 <= not w10774 and w10777;
w10779 <= not w8356 and w10778;
w10780 <= not w6526 and w10778;
w10781 <= not w10779 and not w10780;
w10782 <= a(8) and not w10781;
w10783 <= not a(8) and w10781;
w10784 <= not w10782 and not w10783;
w10785 <= not w10773 and not w10784;
w10786 <= not w2399 and w9266;
w10787 <= not w2506 and w8353;
w10788 <= not w2468 and w8795;
w10789 <= not w10787 and not w10788;
w10790 <= not w10786 and w10789;
w10791 <= w6581 and w8356;
w10792 <= w10790 and not w10791;
w10793 <= a(8) and not w10792;
w10794 <= not w10792 and not w10793;
w10795 <= a(8) and not w10793;
w10796 <= not w10794 and not w10795;
w10797 <= not w10244 and w10255;
w10798 <= not w10256 and not w10797;
w10799 <= not w10796 and w10798;
w10800 <= not w10796 and not w10799;
w10801 <= w10798 and not w10799;
w10802 <= not w10800 and not w10801;
w10803 <= w10241 and not w10243;
w10804 <= not w10244 and not w10803;
w10805 <= not w2468 and w9266;
w10806 <= not w2609 and w8353;
w10807 <= not w2506 and w8795;
w10808 <= not w10806 and not w10807;
w10809 <= not w10805 and w10808;
w10810 <= not w8356 and w10809;
w10811 <= not w6630 and w10809;
w10812 <= not w10810 and not w10811;
w10813 <= a(8) and not w10812;
w10814 <= not a(8) and w10812;
w10815 <= not w10813 and not w10814;
w10816 <= w10804 and not w10815;
w10817 <= not w2764 and w8795;
w10818 <= not w2671 and w9266;
w10819 <= not w10817 and not w10818;
w10820 <= not w7404 and w8356;
w10821 <= w10819 and not w10820;
w10822 <= a(8) and not w10821;
w10823 <= a(8) and not w10822;
w10824 <= not w10821 and not w10822;
w10825 <= not w10823 and not w10824;
w10826 <= not w2764 and not w8351;
w10827 <= a(8) and not w10826;
w10828 <= not w10825 and w10827;
w10829 <= not w2609 and w9266;
w10830 <= not w2764 and w8353;
w10831 <= not w2671 and w8795;
w10832 <= not w10830 and not w10831;
w10833 <= not w10829 and w10832;
w10834 <= not w8356 and w10833;
w10835 <= not w6733 and w10833;
w10836 <= not w10834 and not w10835;
w10837 <= a(8) and not w10836;
w10838 <= not a(8) and w10836;
w10839 <= not w10837 and not w10838;
w10840 <= w10828 and not w10839;
w10841 <= w10242 and w10840;
w10842 <= w10840 and not w10841;
w10843 <= w10242 and not w10841;
w10844 <= not w10842 and not w10843;
w10845 <= not w2506 and w9266;
w10846 <= not w2671 and w8353;
w10847 <= not w2609 and w8795;
w10848 <= not w10846 and not w10847;
w10849 <= not w10845 and w10848;
w10850 <= w6741 and w8356;
w10851 <= w10849 and not w10850;
w10852 <= a(8) and not w10851;
w10853 <= a(8) and not w10852;
w10854 <= not w10851 and not w10852;
w10855 <= not w10853 and not w10854;
w10856 <= not w10844 and not w10855;
w10857 <= not w10841 and not w10856;
w10858 <= not w10804 and w10815;
w10859 <= not w10816 and not w10858;
w10860 <= not w10857 and w10859;
w10861 <= not w10816 and not w10860;
w10862 <= not w10802 and not w10861;
w10863 <= not w10799 and not w10862;
w10864 <= w10773 and w10784;
w10865 <= not w10785 and not w10864;
w10866 <= not w10863 and w10865;
w10867 <= not w10785 and not w10866;
w10868 <= not w10770 and not w10867;
w10869 <= not w10767 and not w10868;
w10870 <= w10741 and not w10753;
w10871 <= not w10752 and not w10753;
w10872 <= not w10870 and not w10871;
w10873 <= not w10869 and not w10872;
w10874 <= not w10753 and not w10873;
w10875 <= w10727 and not w10739;
w10876 <= not w10738 and not w10739;
w10877 <= not w10875 and not w10876;
w10878 <= not w10874 and not w10877;
w10879 <= not w10739 and not w10878;
w10880 <= not w10713 and w10724;
w10881 <= not w10725 and not w10880;
w10882 <= not w10879 and w10881;
w10883 <= not w10725 and not w10882;
w10884 <= not w10711 and not w10883;
w10885 <= not w10708 and not w10884;
w10886 <= not w10693 and not w10885;
w10887 <= not w10690 and not w10886;
w10888 <= not w10675 and not w10887;
w10889 <= not w10672 and not w10888;
w10890 <= w10646 and not w10658;
w10891 <= not w10657 and not w10658;
w10892 <= not w10890 and not w10891;
w10893 <= not w10889 and not w10892;
w10894 <= not w10658 and not w10893;
w10895 <= w10632 and not w10644;
w10896 <= not w10643 and not w10644;
w10897 <= not w10895 and not w10896;
w10898 <= not w10894 and not w10897;
w10899 <= not w10644 and not w10898;
w10900 <= not w10618 and w10629;
w10901 <= not w10630 and not w10900;
w10902 <= not w10899 and w10901;
w10903 <= not w10630 and not w10902;
w10904 <= not w10616 and not w10903;
w10905 <= not w10613 and not w10904;
w10906 <= not w10598 and not w10905;
w10907 <= not w10595 and not w10906;
w10908 <= not w10580 and not w10907;
w10909 <= not w10577 and not w10908;
w10910 <= w10551 and not w10563;
w10911 <= not w10562 and not w10563;
w10912 <= not w10910 and not w10911;
w10913 <= not w10909 and not w10912;
w10914 <= not w10563 and not w10913;
w10915 <= w10537 and not w10549;
w10916 <= not w10548 and not w10549;
w10917 <= not w10915 and not w10916;
w10918 <= not w10914 and not w10917;
w10919 <= not w10549 and not w10918;
w10920 <= not w10523 and w10534;
w10921 <= not w10535 and not w10920;
w10922 <= not w10919 and w10921;
w10923 <= not w10535 and not w10922;
w10924 <= not w10521 and not w10923;
w10925 <= not w10518 and not w10924;
w10926 <= not w10503 and not w10925;
w10927 <= not w10500 and not w10926;
w10928 <= w10474 and not w10486;
w10929 <= not w10485 and not w10486;
w10930 <= not w10928 and not w10929;
w10931 <= not w10927 and not w10930;
w10932 <= not w10486 and not w10931;
w10933 <= w10460 and not w10472;
w10934 <= not w10471 and not w10472;
w10935 <= not w10933 and not w10934;
w10936 <= not w10932 and not w10935;
w10937 <= not w10472 and not w10936;
w10938 <= w10446 and not w10458;
w10939 <= not w10457 and not w10458;
w10940 <= not w10938 and not w10939;
w10941 <= not w10937 and not w10940;
w10942 <= not w10458 and not w10941;
w10943 <= w10432 and not w10444;
w10944 <= not w10443 and not w10444;
w10945 <= not w10943 and not w10944;
w10946 <= not w10942 and not w10945;
w10947 <= not w10444 and not w10946;
w10948 <= w10418 and not w10430;
w10949 <= not w10429 and not w10430;
w10950 <= not w10948 and not w10949;
w10951 <= not w10947 and not w10950;
w10952 <= not w10430 and not w10951;
w10953 <= w10404 and not w10416;
w10954 <= not w10415 and not w10416;
w10955 <= not w10953 and not w10954;
w10956 <= not w10952 and not w10955;
w10957 <= not w10416 and not w10956;
w10958 <= w10390 and not w10402;
w10959 <= not w10401 and not w10402;
w10960 <= not w10958 and not w10959;
w10961 <= not w10957 and not w10960;
w10962 <= not w10402 and not w10961;
w10963 <= w10362 and not w10364;
w10964 <= not w10363 and w10963;
w10965 <= not w10366 and not w10964;
w10966 <= not w10962 and w10965;
w10967 <= w6 and not w4450;
w10968 <= not w3980 and w9802;
w10969 <= not w3812 and w10369;
w10970 <= not w10968 and not w10969;
w10971 <= not w10967 and w10970;
w10972 <= w4650 and w9805;
w10973 <= w10971 and not w10972;
w10974 <= a(5) and not w10973;
w10975 <= not w10973 and not w10974;
w10976 <= a(5) and not w10974;
w10977 <= not w10975 and not w10976;
w10978 <= not w10962 and not w10966;
w10979 <= w10965 and not w10966;
w10980 <= not w10978 and not w10979;
w10981 <= not w10977 and not w10980;
w10982 <= not w10966 and not w10981;
w10983 <= w10381 and not w10383;
w10984 <= not w10384 and not w10983;
w10985 <= not w10982 and w10984;
w10986 <= a(1) and not a(2);
w10987 <= not a(1) and a(2);
w10988 <= not w10986 and not w10987;
w10989 <= not a(0) and not a(1);
w10990 <= not w10988 and w10989;
w10991 <= not w4450 and w10990;
w10992 <= a(0) and not w10988;
w10993 <= w4457 and w10992;
w10994 <= not w10991 and not w10993;
w10995 <= a(2) and not w10994;
w10996 <= not w10994 and not w10995;
w10997 <= a(2) and not w10995;
w10998 <= not w10996 and not w10997;
w10999 <= w6 and not w3812;
w11000 <= not w3899 and w9802;
w11001 <= not w3980 and w10369;
w11002 <= not w11000 and not w11001;
w11003 <= not w10999 and w11002;
w11004 <= w4002 and w9805;
w11005 <= w11003 and not w11004;
w11006 <= a(5) and not w11005;
w11007 <= a(5) and not w11006;
w11008 <= not w11005 and not w11006;
w11009 <= not w11007 and not w11008;
w11010 <= not w10998 and not w11009;
w11011 <= not w10998 and not w11010;
w11012 <= not w11009 and not w11010;
w11013 <= not w11011 and not w11012;
w11014 <= not w10957 and not w10961;
w11015 <= not w10960 and not w10961;
w11016 <= not w11014 and not w11015;
w11017 <= not w11013 and not w11016;
w11018 <= not w11010 and not w11017;
w11019 <= w10977 and not w10979;
w11020 <= not w10978 and w11019;
w11021 <= not w10981 and not w11020;
w11022 <= not w11018 and w11021;
w11023 <= not w11013 and not w11017;
w11024 <= not w11016 and not w11017;
w11025 <= not w11023 and not w11024;
w11026 <= w6 and not w3980;
w11027 <= not w3740 and w9802;
w11028 <= not w3899 and w10369;
w11029 <= not w11027 and not w11028;
w11030 <= not w11026 and w11029;
w11031 <= w4412 and w9805;
w11032 <= w11030 and not w11031;
w11033 <= a(5) and not w11032;
w11034 <= not w11032 and not w11033;
w11035 <= a(5) and not w11033;
w11036 <= not w11034 and not w11035;
w11037 <= not w10952 and not w10956;
w11038 <= not w10955 and not w10956;
w11039 <= not w11037 and not w11038;
w11040 <= not w11036 and not w11039;
w11041 <= not w11036 and not w11040;
w11042 <= not w11039 and not w11040;
w11043 <= not w11041 and not w11042;
w11044 <= w6 and not w3899;
w11045 <= not w3391 and w9802;
w11046 <= not w3740 and w10369;
w11047 <= not w11045 and not w11046;
w11048 <= not w11044 and w11047;
w11049 <= w4493 and w9805;
w11050 <= w11048 and not w11049;
w11051 <= a(5) and not w11050;
w11052 <= not w11050 and not w11051;
w11053 <= a(5) and not w11051;
w11054 <= not w11052 and not w11053;
w11055 <= not w10947 and not w10951;
w11056 <= not w10950 and not w10951;
w11057 <= not w11055 and not w11056;
w11058 <= not w11054 and not w11057;
w11059 <= not w11054 and not w11058;
w11060 <= not w11057 and not w11058;
w11061 <= not w11059 and not w11060;
w11062 <= w6 and not w3740;
w11063 <= not w3540 and w9802;
w11064 <= not w3391 and w10369;
w11065 <= not w11063 and not w11064;
w11066 <= not w11062 and w11065;
w11067 <= w3753 and w9805;
w11068 <= w11066 and not w11067;
w11069 <= a(5) and not w11068;
w11070 <= not w11068 and not w11069;
w11071 <= a(5) and not w11069;
w11072 <= not w11070 and not w11071;
w11073 <= not w10942 and not w10946;
w11074 <= not w10945 and not w10946;
w11075 <= not w11073 and not w11074;
w11076 <= not w11072 and not w11075;
w11077 <= not w11072 and not w11076;
w11078 <= not w11075 and not w11076;
w11079 <= not w11077 and not w11078;
w11080 <= w6 and not w3391;
w11081 <= not w3474 and w9802;
w11082 <= not w3540 and w10369;
w11083 <= not w11081 and not w11082;
w11084 <= not w11080 and w11083;
w11085 <= w3562 and w9805;
w11086 <= w11084 and not w11085;
w11087 <= a(5) and not w11086;
w11088 <= not w11086 and not w11087;
w11089 <= a(5) and not w11087;
w11090 <= not w11088 and not w11089;
w11091 <= not w10937 and not w10941;
w11092 <= not w10940 and not w10941;
w11093 <= not w11091 and not w11092;
w11094 <= not w11090 and not w11093;
w11095 <= not w11090 and not w11094;
w11096 <= not w11093 and not w11094;
w11097 <= not w11095 and not w11096;
w11098 <= w6 and not w3540;
w11099 <= not w2947 and w9802;
w11100 <= not w3474 and w10369;
w11101 <= not w11099 and not w11100;
w11102 <= not w11098 and w11101;
w11103 <= w4019 and w9805;
w11104 <= w11102 and not w11103;
w11105 <= a(5) and not w11104;
w11106 <= not w11104 and not w11105;
w11107 <= a(5) and not w11105;
w11108 <= not w11106 and not w11107;
w11109 <= not w10932 and not w10936;
w11110 <= not w10935 and not w10936;
w11111 <= not w11109 and not w11110;
w11112 <= not w11108 and not w11111;
w11113 <= not w11108 and not w11112;
w11114 <= not w11111 and not w11112;
w11115 <= not w11113 and not w11114;
w11116 <= w6 and not w3474;
w11117 <= not w327 and w9802;
w11118 <= not w2947 and w10369;
w11119 <= not w11117 and not w11118;
w11120 <= not w11116 and w11119;
w11121 <= w3650 and w9805;
w11122 <= w11120 and not w11121;
w11123 <= a(5) and not w11122;
w11124 <= not w11122 and not w11123;
w11125 <= a(5) and not w11123;
w11126 <= not w11124 and not w11125;
w11127 <= not w10927 and not w10931;
w11128 <= not w10930 and not w10931;
w11129 <= not w11127 and not w11128;
w11130 <= not w11126 and not w11129;
w11131 <= not w11126 and not w11130;
w11132 <= not w11129 and not w11130;
w11133 <= not w11131 and not w11132;
w11134 <= w10503 and w10925;
w11135 <= not w10926 and not w11134;
w11136 <= w6 and not w2947;
w11137 <= not w522 and w9802;
w11138 <= not w327 and w10369;
w11139 <= not w11137 and not w11138;
w11140 <= not w11136 and w11139;
w11141 <= not w9805 and w11140;
w11142 <= not w2953 and w11140;
w11143 <= not w11141 and not w11142;
w11144 <= a(5) and not w11143;
w11145 <= not a(5) and w11143;
w11146 <= not w11144 and not w11145;
w11147 <= w11135 and not w11146;
w11148 <= w10521 and w10923;
w11149 <= not w10924 and not w11148;
w11150 <= w6 and not w327;
w11151 <= not w645 and w9802;
w11152 <= not w522 and w10369;
w11153 <= not w11151 and not w11152;
w11154 <= not w11150 and w11153;
w11155 <= not w9805 and w11154;
w11156 <= not w3282 and w11154;
w11157 <= not w11155 and not w11156;
w11158 <= a(5) and not w11157;
w11159 <= not a(5) and w11157;
w11160 <= not w11158 and not w11159;
w11161 <= w11149 and not w11160;
w11162 <= w6 and not w522;
w11163 <= not w802 and w9802;
w11164 <= not w645 and w10369;
w11165 <= not w11163 and not w11164;
w11166 <= not w11162 and w11165;
w11167 <= w3266 and w9805;
w11168 <= w11166 and not w11167;
w11169 <= a(5) and not w11168;
w11170 <= not w11168 and not w11169;
w11171 <= a(5) and not w11169;
w11172 <= not w11170 and not w11171;
w11173 <= w10919 and not w10921;
w11174 <= not w10922 and not w11173;
w11175 <= not w11172 and w11174;
w11176 <= not w11172 and not w11175;
w11177 <= w11174 and not w11175;
w11178 <= not w11176 and not w11177;
w11179 <= w6 and not w645;
w11180 <= not w893 and w9802;
w11181 <= not w802 and w10369;
w11182 <= not w11180 and not w11181;
w11183 <= not w11179 and w11182;
w11184 <= w4114 and w9805;
w11185 <= w11183 and not w11184;
w11186 <= a(5) and not w11185;
w11187 <= not w11185 and not w11186;
w11188 <= a(5) and not w11186;
w11189 <= not w11187 and not w11188;
w11190 <= not w10914 and not w10918;
w11191 <= not w10917 and not w10918;
w11192 <= not w11190 and not w11191;
w11193 <= not w11189 and not w11192;
w11194 <= not w11189 and not w11193;
w11195 <= not w11192 and not w11193;
w11196 <= not w11194 and not w11195;
w11197 <= w6 and not w802;
w11198 <= not w995 and w9802;
w11199 <= not w893 and w10369;
w11200 <= not w11198 and not w11199;
w11201 <= not w11197 and w11200;
w11202 <= w4139 and w9805;
w11203 <= w11201 and not w11202;
w11204 <= a(5) and not w11203;
w11205 <= not w11203 and not w11204;
w11206 <= a(5) and not w11204;
w11207 <= not w11205 and not w11206;
w11208 <= not w10909 and not w10913;
w11209 <= not w10912 and not w10913;
w11210 <= not w11208 and not w11209;
w11211 <= not w11207 and not w11210;
w11212 <= not w11207 and not w11211;
w11213 <= not w11210 and not w11211;
w11214 <= not w11212 and not w11213;
w11215 <= w10580 and w10907;
w11216 <= not w10908 and not w11215;
w11217 <= w6 and not w893;
w11218 <= not w1113 and w9802;
w11219 <= not w995 and w10369;
w11220 <= not w11218 and not w11219;
w11221 <= not w11217 and w11220;
w11222 <= not w9805 and w11221;
w11223 <= not w4568 and w11221;
w11224 <= not w11222 and not w11223;
w11225 <= a(5) and not w11224;
w11226 <= not a(5) and w11224;
w11227 <= not w11225 and not w11226;
w11228 <= w11216 and not w11227;
w11229 <= w10598 and w10905;
w11230 <= not w10906 and not w11229;
w11231 <= w6 and not w995;
w11232 <= not w1170 and w9802;
w11233 <= not w1113 and w10369;
w11234 <= not w11232 and not w11233;
w11235 <= not w11231 and w11234;
w11236 <= not w9805 and w11235;
w11237 <= not w4364 and w11235;
w11238 <= not w11236 and not w11237;
w11239 <= a(5) and not w11238;
w11240 <= not a(5) and w11238;
w11241 <= not w11239 and not w11240;
w11242 <= w11230 and not w11241;
w11243 <= w10616 and w10903;
w11244 <= not w10904 and not w11243;
w11245 <= w6 and not w1113;
w11246 <= not w1299 and w9802;
w11247 <= not w1170 and w10369;
w11248 <= not w11246 and not w11247;
w11249 <= not w11245 and w11248;
w11250 <= not w9805 and w11249;
w11251 <= not w4796 and w11249;
w11252 <= not w11250 and not w11251;
w11253 <= a(5) and not w11252;
w11254 <= not a(5) and w11252;
w11255 <= not w11253 and not w11254;
w11256 <= w11244 and not w11255;
w11257 <= w6 and not w1170;
w11258 <= not w1407 and w9802;
w11259 <= not w1299 and w10369;
w11260 <= not w11258 and not w11259;
w11261 <= not w11257 and w11260;
w11262 <= w4783 and w9805;
w11263 <= w11261 and not w11262;
w11264 <= a(5) and not w11263;
w11265 <= not w11263 and not w11264;
w11266 <= a(5) and not w11264;
w11267 <= not w11265 and not w11266;
w11268 <= w10899 and not w10901;
w11269 <= not w10902 and not w11268;
w11270 <= not w11267 and w11269;
w11271 <= not w11267 and not w11270;
w11272 <= w11269 and not w11270;
w11273 <= not w11271 and not w11272;
w11274 <= w6 and not w1299;
w11275 <= not w1507 and w9802;
w11276 <= not w1407 and w10369;
w11277 <= not w11275 and not w11276;
w11278 <= not w11274 and w11277;
w11279 <= w5049 and w9805;
w11280 <= w11278 and not w11279;
w11281 <= a(5) and not w11280;
w11282 <= not w11280 and not w11281;
w11283 <= a(5) and not w11281;
w11284 <= not w11282 and not w11283;
w11285 <= not w10894 and not w10898;
w11286 <= not w10897 and not w10898;
w11287 <= not w11285 and not w11286;
w11288 <= not w11284 and not w11287;
w11289 <= not w11284 and not w11288;
w11290 <= not w11287 and not w11288;
w11291 <= not w11289 and not w11290;
w11292 <= w6 and not w1407;
w11293 <= not w1600 and w9802;
w11294 <= not w1507 and w10369;
w11295 <= not w11293 and not w11294;
w11296 <= not w11292 and w11295;
w11297 <= w5074 and w9805;
w11298 <= w11296 and not w11297;
w11299 <= a(5) and not w11298;
w11300 <= not w11298 and not w11299;
w11301 <= a(5) and not w11299;
w11302 <= not w11300 and not w11301;
w11303 <= not w10889 and not w10893;
w11304 <= not w10892 and not w10893;
w11305 <= not w11303 and not w11304;
w11306 <= not w11302 and not w11305;
w11307 <= not w11302 and not w11306;
w11308 <= not w11305 and not w11306;
w11309 <= not w11307 and not w11308;
w11310 <= w10675 and w10887;
w11311 <= not w10888 and not w11310;
w11312 <= w6 and not w1507;
w11313 <= not w1714 and w9802;
w11314 <= not w1600 and w10369;
w11315 <= not w11313 and not w11314;
w11316 <= not w11312 and w11315;
w11317 <= not w9805 and w11316;
w11318 <= not w5496 and w11316;
w11319 <= not w11317 and not w11318;
w11320 <= a(5) and not w11319;
w11321 <= not a(5) and w11319;
w11322 <= not w11320 and not w11321;
w11323 <= w11311 and not w11322;
w11324 <= w10693 and w10885;
w11325 <= not w10886 and not w11324;
w11326 <= w6 and not w1600;
w11327 <= not w1812 and w9802;
w11328 <= not w1714 and w10369;
w11329 <= not w11327 and not w11328;
w11330 <= not w11326 and w11329;
w11331 <= not w9805 and w11330;
w11332 <= not w5263 and w11330;
w11333 <= not w11331 and not w11332;
w11334 <= a(5) and not w11333;
w11335 <= not a(5) and w11333;
w11336 <= not w11334 and not w11335;
w11337 <= w11325 and not w11336;
w11338 <= w10711 and w10883;
w11339 <= not w10884 and not w11338;
w11340 <= w6 and not w1714;
w11341 <= not w1848 and w9802;
w11342 <= not w1812 and w10369;
w11343 <= not w11341 and not w11342;
w11344 <= not w11340 and w11343;
w11345 <= not w9805 and w11344;
w11346 <= not w5786 and w11344;
w11347 <= not w11345 and not w11346;
w11348 <= a(5) and not w11347;
w11349 <= not a(5) and w11347;
w11350 <= not w11348 and not w11349;
w11351 <= w11339 and not w11350;
w11352 <= w6 and not w1812;
w11353 <= not w1927 and w9802;
w11354 <= not w1848 and w10369;
w11355 <= not w11353 and not w11354;
w11356 <= not w11352 and w11355;
w11357 <= w5942 and w9805;
w11358 <= w11356 and not w11357;
w11359 <= a(5) and not w11358;
w11360 <= not w11358 and not w11359;
w11361 <= a(5) and not w11359;
w11362 <= not w11360 and not w11361;
w11363 <= w10879 and not w10881;
w11364 <= not w10882 and not w11363;
w11365 <= not w11362 and w11364;
w11366 <= not w11362 and not w11365;
w11367 <= w11364 and not w11365;
w11368 <= not w11366 and not w11367;
w11369 <= w6 and not w1848;
w11370 <= not w1992 and w9802;
w11371 <= not w1927 and w10369;
w11372 <= not w11370 and not w11371;
w11373 <= not w11369 and w11372;
w11374 <= w5769 and w9805;
w11375 <= w11373 and not w11374;
w11376 <= a(5) and not w11375;
w11377 <= not w11375 and not w11376;
w11378 <= a(5) and not w11376;
w11379 <= not w11377 and not w11378;
w11380 <= not w10874 and not w10878;
w11381 <= not w10877 and not w10878;
w11382 <= not w11380 and not w11381;
w11383 <= not w11379 and not w11382;
w11384 <= not w11379 and not w11383;
w11385 <= not w11382 and not w11383;
w11386 <= not w11384 and not w11385;
w11387 <= w6 and not w1927;
w11388 <= not w2087 and w9802;
w11389 <= not w1992 and w10369;
w11390 <= not w11388 and not w11389;
w11391 <= not w11387 and w11390;
w11392 <= w6078 and w9805;
w11393 <= w11391 and not w11392;
w11394 <= a(5) and not w11393;
w11395 <= not w11393 and not w11394;
w11396 <= a(5) and not w11394;
w11397 <= not w11395 and not w11396;
w11398 <= not w10869 and not w10873;
w11399 <= not w10872 and not w10873;
w11400 <= not w11398 and not w11399;
w11401 <= not w11397 and not w11400;
w11402 <= not w11397 and not w11401;
w11403 <= not w11400 and not w11401;
w11404 <= not w11402 and not w11403;
w11405 <= w10770 and w10867;
w11406 <= not w10868 and not w11405;
w11407 <= w6 and not w1992;
w11408 <= not w2124 and w9802;
w11409 <= not w2087 and w10369;
w11410 <= not w11408 and not w11409;
w11411 <= not w11407 and w11410;
w11412 <= not w9805 and w11411;
w11413 <= not w6414 and w11411;
w11414 <= not w11412 and not w11413;
w11415 <= a(5) and not w11414;
w11416 <= not a(5) and w11414;
w11417 <= not w11415 and not w11416;
w11418 <= w11406 and not w11417;
w11419 <= w10863 and not w10865;
w11420 <= not w10866 and not w11419;
w11421 <= w6 and not w2087;
w11422 <= not w2226 and w9802;
w11423 <= not w2124 and w10369;
w11424 <= not w11422 and not w11423;
w11425 <= not w11421 and w11424;
w11426 <= not w9805 and w11425;
w11427 <= not w6427 and w11425;
w11428 <= not w11426 and not w11427;
w11429 <= a(5) and not w11428;
w11430 <= not a(5) and w11428;
w11431 <= not w11429 and not w11430;
w11432 <= w11420 and not w11431;
w11433 <= w10802 and w10861;
w11434 <= not w10862 and not w11433;
w11435 <= w6 and not w2124;
w11436 <= not w2323 and w9802;
w11437 <= not w2226 and w10369;
w11438 <= not w11436 and not w11437;
w11439 <= not w11435 and w11438;
w11440 <= not w9805 and w11439;
w11441 <= not w6057 and w11439;
w11442 <= not w11440 and not w11441;
w11443 <= a(5) and not w11442;
w11444 <= not a(5) and w11442;
w11445 <= not w11443 and not w11444;
w11446 <= w11434 and not w11445;
w11447 <= w6 and not w2226;
w11448 <= not w2399 and w9802;
w11449 <= not w2323 and w10369;
w11450 <= not w11448 and not w11449;
w11451 <= not w11447 and w11450;
w11452 <= w6476 and w9805;
w11453 <= w11451 and not w11452;
w11454 <= a(5) and not w11453;
w11455 <= not w11453 and not w11454;
w11456 <= a(5) and not w11454;
w11457 <= not w11455 and not w11456;
w11458 <= w10857 and not w10859;
w11459 <= not w10860 and not w11458;
w11460 <= not w11457 and w11459;
w11461 <= not w11457 and not w11460;
w11462 <= w11459 and not w11460;
w11463 <= not w11461 and not w11462;
w11464 <= not w10844 and not w10856;
w11465 <= not w10855 and not w10856;
w11466 <= not w11464 and not w11465;
w11467 <= w6 and not w2323;
w11468 <= not w2468 and w9802;
w11469 <= not w2399 and w10369;
w11470 <= not w11468 and not w11469;
w11471 <= not w11467 and w11470;
w11472 <= not w9805 and w11471;
w11473 <= not w6526 and w11471;
w11474 <= not w11472 and not w11473;
w11475 <= a(5) and not w11474;
w11476 <= not a(5) and w11474;
w11477 <= not w11475 and not w11476;
w11478 <= not w11466 and not w11477;
w11479 <= w6 and not w2399;
w11480 <= not w2506 and w9802;
w11481 <= not w2468 and w10369;
w11482 <= not w11480 and not w11481;
w11483 <= not w11479 and w11482;
w11484 <= w6581 and w9805;
w11485 <= w11483 and not w11484;
w11486 <= a(5) and not w11485;
w11487 <= not w11485 and not w11486;
w11488 <= a(5) and not w11486;
w11489 <= not w11487 and not w11488;
w11490 <= not w10828 and w10839;
w11491 <= not w10840 and not w11490;
w11492 <= not w11489 and w11491;
w11493 <= not w11489 and not w11492;
w11494 <= w11491 and not w11492;
w11495 <= not w11493 and not w11494;
w11496 <= w10825 and not w10827;
w11497 <= not w10828 and not w11496;
w11498 <= w6 and not w2468;
w11499 <= not w2609 and w9802;
w11500 <= not w2506 and w10369;
w11501 <= not w11499 and not w11500;
w11502 <= not w11498 and w11501;
w11503 <= not w9805 and w11502;
w11504 <= not w6630 and w11502;
w11505 <= not w11503 and not w11504;
w11506 <= a(5) and not w11505;
w11507 <= not a(5) and w11505;
w11508 <= not w11506 and not w11507;
w11509 <= w11497 and not w11508;
w11510 <= not w2764 and w10369;
w11511 <= w6 and not w2671;
w11512 <= not w11510 and not w11511;
w11513 <= not w7404 and w9805;
w11514 <= w11512 and not w11513;
w11515 <= a(5) and not w11514;
w11516 <= a(5) and not w11515;
w11517 <= not w11514 and not w11515;
w11518 <= not w11516 and not w11517;
w11519 <= not w5 and not w2764;
w11520 <= a(5) and not w11519;
w11521 <= not w11518 and w11520;
w11522 <= w6 and not w2609;
w11523 <= not w2764 and w9802;
w11524 <= not w2671 and w10369;
w11525 <= not w11523 and not w11524;
w11526 <= not w11522 and w11525;
w11527 <= not w9805 and w11526;
w11528 <= not w6733 and w11526;
w11529 <= not w11527 and not w11528;
w11530 <= a(5) and not w11529;
w11531 <= not a(5) and w11529;
w11532 <= not w11530 and not w11531;
w11533 <= w11521 and not w11532;
w11534 <= w10826 and w11533;
w11535 <= w11533 and not w11534;
w11536 <= w10826 and not w11534;
w11537 <= not w11535 and not w11536;
w11538 <= w6 and not w2506;
w11539 <= not w2671 and w9802;
w11540 <= not w2609 and w10369;
w11541 <= not w11539 and not w11540;
w11542 <= not w11538 and w11541;
w11543 <= w6741 and w9805;
w11544 <= w11542 and not w11543;
w11545 <= a(5) and not w11544;
w11546 <= a(5) and not w11545;
w11547 <= not w11544 and not w11545;
w11548 <= not w11546 and not w11547;
w11549 <= not w11537 and not w11548;
w11550 <= not w11534 and not w11549;
w11551 <= not w11497 and w11508;
w11552 <= not w11509 and not w11551;
w11553 <= not w11550 and w11552;
w11554 <= not w11509 and not w11553;
w11555 <= not w11495 and not w11554;
w11556 <= not w11492 and not w11555;
w11557 <= w11466 and w11477;
w11558 <= not w11478 and not w11557;
w11559 <= not w11556 and w11558;
w11560 <= not w11478 and not w11559;
w11561 <= not w11463 and not w11560;
w11562 <= not w11460 and not w11561;
w11563 <= w11434 and not w11446;
w11564 <= not w11445 and not w11446;
w11565 <= not w11563 and not w11564;
w11566 <= not w11562 and not w11565;
w11567 <= not w11446 and not w11566;
w11568 <= w11420 and not w11432;
w11569 <= not w11431 and not w11432;
w11570 <= not w11568 and not w11569;
w11571 <= not w11567 and not w11570;
w11572 <= not w11432 and not w11571;
w11573 <= not w11406 and w11417;
w11574 <= not w11418 and not w11573;
w11575 <= not w11572 and w11574;
w11576 <= not w11418 and not w11575;
w11577 <= not w11404 and not w11576;
w11578 <= not w11401 and not w11577;
w11579 <= not w11386 and not w11578;
w11580 <= not w11383 and not w11579;
w11581 <= not w11368 and not w11580;
w11582 <= not w11365 and not w11581;
w11583 <= w11339 and not w11351;
w11584 <= not w11350 and not w11351;
w11585 <= not w11583 and not w11584;
w11586 <= not w11582 and not w11585;
w11587 <= not w11351 and not w11586;
w11588 <= w11325 and not w11337;
w11589 <= not w11336 and not w11337;
w11590 <= not w11588 and not w11589;
w11591 <= not w11587 and not w11590;
w11592 <= not w11337 and not w11591;
w11593 <= not w11311 and w11322;
w11594 <= not w11323 and not w11593;
w11595 <= not w11592 and w11594;
w11596 <= not w11323 and not w11595;
w11597 <= not w11309 and not w11596;
w11598 <= not w11306 and not w11597;
w11599 <= not w11291 and not w11598;
w11600 <= not w11288 and not w11599;
w11601 <= not w11273 and not w11600;
w11602 <= not w11270 and not w11601;
w11603 <= w11244 and not w11256;
w11604 <= not w11255 and not w11256;
w11605 <= not w11603 and not w11604;
w11606 <= not w11602 and not w11605;
w11607 <= not w11256 and not w11606;
w11608 <= w11230 and not w11242;
w11609 <= not w11241 and not w11242;
w11610 <= not w11608 and not w11609;
w11611 <= not w11607 and not w11610;
w11612 <= not w11242 and not w11611;
w11613 <= not w11216 and w11227;
w11614 <= not w11228 and not w11613;
w11615 <= not w11612 and w11614;
w11616 <= not w11228 and not w11615;
w11617 <= not w11214 and not w11616;
w11618 <= not w11211 and not w11617;
w11619 <= not w11196 and not w11618;
w11620 <= not w11193 and not w11619;
w11621 <= not w11178 and not w11620;
w11622 <= not w11175 and not w11621;
w11623 <= w11149 and not w11161;
w11624 <= not w11160 and not w11161;
w11625 <= not w11623 and not w11624;
w11626 <= not w11622 and not w11625;
w11627 <= not w11161 and not w11626;
w11628 <= not w11135 and w11146;
w11629 <= not w11147 and not w11628;
w11630 <= not w11627 and w11629;
w11631 <= not w11147 and not w11630;
w11632 <= not w11133 and not w11631;
w11633 <= not w11130 and not w11632;
w11634 <= not w11115 and not w11633;
w11635 <= not w11112 and not w11634;
w11636 <= not w11097 and not w11635;
w11637 <= not w11094 and not w11636;
w11638 <= not w11079 and not w11637;
w11639 <= not w11076 and not w11638;
w11640 <= not w11061 and not w11639;
w11641 <= not w11058 and not w11640;
w11642 <= not w11043 and not w11641;
w11643 <= not w11040 and not w11642;
w11644 <= not w11025 and not w11643;
w11645 <= w11025 and w11643;
w11646 <= not w11644 and not w11645;
w11647 <= w11043 and w11641;
w11648 <= not w11642 and not w11647;
w11649 <= not w3812 and w10990;
w11650 <= not a(0) and a(1);
w11651 <= not w4450 and w11650;
w11652 <= not w11649 and not w11651;
w11653 <= not w10992 and w11652;
w11654 <= not w4544 and w11652;
w11655 <= not w11653 and not w11654;
w11656 <= a(2) and not w11655;
w11657 <= not a(2) and w11655;
w11658 <= not w11656 and not w11657;
w11659 <= w11648 and not w11658;
w11660 <= w11061 and w11639;
w11661 <= not w11640 and not w11660;
w11662 <= a(0) and w10988;
w11663 <= not w4450 and w11662;
w11664 <= not w3980 and w10990;
w11665 <= not w3812 and w11650;
w11666 <= not w11664 and not w11665;
w11667 <= not w11663 and w11666;
w11668 <= not w10992 and w11667;
w11669 <= not w4650 and w11667;
w11670 <= not w11668 and not w11669;
w11671 <= a(2) and not w11670;
w11672 <= not a(2) and w11670;
w11673 <= not w11671 and not w11672;
w11674 <= w11661 and not w11673;
w11675 <= w11079 and w11637;
w11676 <= not w11638 and not w11675;
w11677 <= not w3812 and w11662;
w11678 <= not w3899 and w10990;
w11679 <= not w3980 and w11650;
w11680 <= not w11678 and not w11679;
w11681 <= not w11677 and w11680;
w11682 <= not w10992 and w11681;
w11683 <= not w4002 and w11681;
w11684 <= not w11682 and not w11683;
w11685 <= a(2) and not w11684;
w11686 <= not a(2) and w11684;
w11687 <= not w11685 and not w11686;
w11688 <= w11676 and not w11687;
w11689 <= w11097 and w11635;
w11690 <= not w11636 and not w11689;
w11691 <= not w3980 and w11662;
w11692 <= not w3740 and w10990;
w11693 <= not w3899 and w11650;
w11694 <= not w11692 and not w11693;
w11695 <= not w11691 and w11694;
w11696 <= not w10992 and w11695;
w11697 <= not w4412 and w11695;
w11698 <= not w11696 and not w11697;
w11699 <= a(2) and not w11698;
w11700 <= not a(2) and w11698;
w11701 <= not w11699 and not w11700;
w11702 <= w11690 and not w11701;
w11703 <= w11115 and w11633;
w11704 <= not w11634 and not w11703;
w11705 <= not w3899 and w11662;
w11706 <= not w3391 and w10990;
w11707 <= not w3740 and w11650;
w11708 <= not w11706 and not w11707;
w11709 <= not w11705 and w11708;
w11710 <= not w10992 and w11709;
w11711 <= not w4493 and w11709;
w11712 <= not w11710 and not w11711;
w11713 <= a(2) and not w11712;
w11714 <= not a(2) and w11712;
w11715 <= not w11713 and not w11714;
w11716 <= w11704 and not w11715;
w11717 <= w11627 and not w11629;
w11718 <= not w11630 and not w11717;
w11719 <= w11612 and not w11614;
w11720 <= not w11615 and not w11719;
w11721 <= w11592 and not w11594;
w11722 <= not w11595 and not w11721;
w11723 <= w11572 and not w11574;
w11724 <= not w11575 and not w11723;
w11725 <= w11550 and not w11552;
w11726 <= not w11553 and not w11725;
w11727 <= not w11521 and w11532;
w11728 <= not w11533 and not w11727;
w11729 <= not w10992 and not w11662;
w11730 <= not w2764 and not w11729;
w11731 <= a(2) and w10992;
w11732 <= w6733 and w11731;
w11733 <= not w2609 and w11662;
w11734 <= not w2764 and w10990;
w11735 <= not w2671 and w11650;
w11736 <= not w11734 and not w11735;
w11737 <= not w11733 and w11736;
w11738 <= a(2) and not w11737;
w11739 <= not w7404 and w11731;
w11740 <= a(2) and w11650;
w11741 <= not w2764 and w11740;
w11742 <= a(2) and w11662;
w11743 <= not w2671 and w11742;
w11744 <= a(2) and not w11743;
w11745 <= not w11741 and w11744;
w11746 <= not w11739 and w11745;
w11747 <= not w11738 and w11746;
w11748 <= not w11732 and w11747;
w11749 <= not w11730 and w11748;
w11750 <= w11519 and w11749;
w11751 <= not w11519 and not w11749;
w11752 <= not w2506 and w11662;
w11753 <= not w2671 and w10990;
w11754 <= not w2609 and w11650;
w11755 <= not w11753 and not w11754;
w11756 <= not w11752 and w11755;
w11757 <= w6741 and w10992;
w11758 <= w11756 and not w11757;
w11759 <= not a(2) and not w11758;
w11760 <= a(2) and w11758;
w11761 <= not w11759 and not w11760;
w11762 <= not w11751 and not w11761;
w11763 <= not w11750 and not w11762;
w11764 <= not w2468 and w11662;
w11765 <= not w2609 and w10990;
w11766 <= not w2506 and w11650;
w11767 <= not w11765 and not w11766;
w11768 <= not w11764 and w11767;
w11769 <= not w10992 and w11768;
w11770 <= not w6630 and w11768;
w11771 <= not w11769 and not w11770;
w11772 <= a(2) and not w11771;
w11773 <= not a(2) and w11771;
w11774 <= not w11772 and not w11773;
w11775 <= w11763 and w11774;
w11776 <= w11518 and not w11520;
w11777 <= not w11521 and not w11776;
w11778 <= not w11775 and w11777;
w11779 <= not w11763 and not w11774;
w11780 <= not w11778 and not w11779;
w11781 <= w11728 and not w11780;
w11782 <= not w11728 and w11780;
w11783 <= not w2399 and w11662;
w11784 <= not w2506 and w10990;
w11785 <= not w2468 and w11650;
w11786 <= not w11784 and not w11785;
w11787 <= not w11783 and w11786;
w11788 <= w6581 and w10992;
w11789 <= w11787 and not w11788;
w11790 <= not a(2) and not w11789;
w11791 <= a(2) and w11789;
w11792 <= not w11790 and not w11791;
w11793 <= not w11782 and not w11792;
w11794 <= not w11781 and not w11793;
w11795 <= not w2323 and w11662;
w11796 <= not w2468 and w10990;
w11797 <= not w2399 and w11650;
w11798 <= not w11796 and not w11797;
w11799 <= not w11795 and w11798;
w11800 <= not w10992 and w11799;
w11801 <= not w6526 and w11799;
w11802 <= not w11800 and not w11801;
w11803 <= a(2) and not w11802;
w11804 <= not a(2) and w11802;
w11805 <= not w11803 and not w11804;
w11806 <= not w11794 and not w11805;
w11807 <= w11794 and w11805;
w11808 <= w11537 and w11548;
w11809 <= not w11549 and not w11808;
w11810 <= not w11807 and w11809;
w11811 <= not w11806 and not w11810;
w11812 <= w11726 and not w11811;
w11813 <= not w11726 and w11811;
w11814 <= not w2226 and w11662;
w11815 <= not w2399 and w10990;
w11816 <= not w2323 and w11650;
w11817 <= not w11815 and not w11816;
w11818 <= not w11814 and w11817;
w11819 <= w6476 and w10992;
w11820 <= w11818 and not w11819;
w11821 <= not a(2) and not w11820;
w11822 <= a(2) and w11820;
w11823 <= not w11821 and not w11822;
w11824 <= not w11813 and not w11823;
w11825 <= not w11812 and not w11824;
w11826 <= not w2124 and w11662;
w11827 <= not w2323 and w10990;
w11828 <= not w2226 and w11650;
w11829 <= not w11827 and not w11828;
w11830 <= not w11826 and w11829;
w11831 <= not w10992 and w11830;
w11832 <= not w6057 and w11830;
w11833 <= not w11831 and not w11832;
w11834 <= a(2) and not w11833;
w11835 <= not a(2) and w11833;
w11836 <= not w11834 and not w11835;
w11837 <= w11825 and w11836;
w11838 <= w11495 and w11554;
w11839 <= not w11555 and not w11838;
w11840 <= not w11837 and w11839;
w11841 <= not w11825 and not w11836;
w11842 <= not w11840 and not w11841;
w11843 <= not w2087 and w11662;
w11844 <= not w2226 and w10990;
w11845 <= not w2124 and w11650;
w11846 <= not w11844 and not w11845;
w11847 <= not w11843 and w11846;
w11848 <= not w10992 and w11847;
w11849 <= not w6427 and w11847;
w11850 <= not w11848 and not w11849;
w11851 <= a(2) and not w11850;
w11852 <= not a(2) and w11850;
w11853 <= not w11851 and not w11852;
w11854 <= w11842 and w11853;
w11855 <= w11556 and not w11558;
w11856 <= not w11559 and not w11855;
w11857 <= not w11854 and w11856;
w11858 <= not w11842 and not w11853;
w11859 <= not w11857 and not w11858;
w11860 <= not w1992 and w11662;
w11861 <= not w2124 and w10990;
w11862 <= not w2087 and w11650;
w11863 <= not w11861 and not w11862;
w11864 <= not w11860 and w11863;
w11865 <= not w10992 and w11864;
w11866 <= not w6414 and w11864;
w11867 <= not w11865 and not w11866;
w11868 <= a(2) and not w11867;
w11869 <= not a(2) and w11867;
w11870 <= not w11868 and not w11869;
w11871 <= w11859 and w11870;
w11872 <= w11463 and w11560;
w11873 <= not w11561 and not w11872;
w11874 <= not w11871 and w11873;
w11875 <= not w11859 and not w11870;
w11876 <= not w11874 and not w11875;
w11877 <= w11562 and not w11564;
w11878 <= not w11563 and w11877;
w11879 <= not w11566 and not w11878;
w11880 <= not w11876 and w11879;
w11881 <= w11876 and not w11879;
w11882 <= not w1927 and w11662;
w11883 <= not w2087 and w10990;
w11884 <= not w1992 and w11650;
w11885 <= not w11883 and not w11884;
w11886 <= not w11882 and w11885;
w11887 <= w6078 and w10992;
w11888 <= w11886 and not w11887;
w11889 <= not a(2) and not w11888;
w11890 <= a(2) and w11888;
w11891 <= not w11889 and not w11890;
w11892 <= not w11881 and not w11891;
w11893 <= not w11880 and not w11892;
w11894 <= w11567 and not w11569;
w11895 <= not w11568 and w11894;
w11896 <= not w11571 and not w11895;
w11897 <= not w11893 and w11896;
w11898 <= w11893 and not w11896;
w11899 <= not w1848 and w11662;
w11900 <= not w1992 and w10990;
w11901 <= not w1927 and w11650;
w11902 <= not w11900 and not w11901;
w11903 <= not w11899 and w11902;
w11904 <= w5769 and w10992;
w11905 <= w11903 and not w11904;
w11906 <= not a(2) and not w11905;
w11907 <= a(2) and w11905;
w11908 <= not w11906 and not w11907;
w11909 <= not w11898 and not w11908;
w11910 <= not w11897 and not w11909;
w11911 <= w11724 and not w11910;
w11912 <= not w11724 and w11910;
w11913 <= not w1812 and w11662;
w11914 <= not w1927 and w10990;
w11915 <= not w1848 and w11650;
w11916 <= not w11914 and not w11915;
w11917 <= not w11913 and w11916;
w11918 <= w5942 and w10992;
w11919 <= w11917 and not w11918;
w11920 <= not a(2) and not w11919;
w11921 <= a(2) and w11919;
w11922 <= not w11920 and not w11921;
w11923 <= not w11912 and not w11922;
w11924 <= not w11911 and not w11923;
w11925 <= not w1714 and w11662;
w11926 <= not w1848 and w10990;
w11927 <= not w1812 and w11650;
w11928 <= not w11926 and not w11927;
w11929 <= not w11925 and w11928;
w11930 <= not w10992 and w11929;
w11931 <= not w5786 and w11929;
w11932 <= not w11930 and not w11931;
w11933 <= a(2) and not w11932;
w11934 <= not a(2) and w11932;
w11935 <= not w11933 and not w11934;
w11936 <= w11924 and w11935;
w11937 <= w11404 and w11576;
w11938 <= not w11577 and not w11937;
w11939 <= not w11936 and w11938;
w11940 <= not w11924 and not w11935;
w11941 <= not w11939 and not w11940;
w11942 <= not w1600 and w11662;
w11943 <= not w1812 and w10990;
w11944 <= not w1714 and w11650;
w11945 <= not w11943 and not w11944;
w11946 <= not w11942 and w11945;
w11947 <= not w10992 and w11946;
w11948 <= not w5263 and w11946;
w11949 <= not w11947 and not w11948;
w11950 <= a(2) and not w11949;
w11951 <= not a(2) and w11949;
w11952 <= not w11950 and not w11951;
w11953 <= w11941 and w11952;
w11954 <= w11386 and w11578;
w11955 <= not w11579 and not w11954;
w11956 <= not w11953 and w11955;
w11957 <= not w11941 and not w11952;
w11958 <= not w11956 and not w11957;
w11959 <= not w1507 and w11662;
w11960 <= not w1714 and w10990;
w11961 <= not w1600 and w11650;
w11962 <= not w11960 and not w11961;
w11963 <= not w11959 and w11962;
w11964 <= not w10992 and w11963;
w11965 <= not w5496 and w11963;
w11966 <= not w11964 and not w11965;
w11967 <= a(2) and not w11966;
w11968 <= not a(2) and w11966;
w11969 <= not w11967 and not w11968;
w11970 <= w11958 and w11969;
w11971 <= w11368 and w11580;
w11972 <= not w11581 and not w11971;
w11973 <= not w11970 and w11972;
w11974 <= not w11958 and not w11969;
w11975 <= not w11973 and not w11974;
w11976 <= w11582 and not w11584;
w11977 <= not w11583 and w11976;
w11978 <= not w11586 and not w11977;
w11979 <= not w11975 and w11978;
w11980 <= w11975 and not w11978;
w11981 <= not w1407 and w11662;
w11982 <= not w1600 and w10990;
w11983 <= not w1507 and w11650;
w11984 <= not w11982 and not w11983;
w11985 <= not w11981 and w11984;
w11986 <= w5074 and w10992;
w11987 <= w11985 and not w11986;
w11988 <= not a(2) and not w11987;
w11989 <= a(2) and w11987;
w11990 <= not w11988 and not w11989;
w11991 <= not w11980 and not w11990;
w11992 <= not w11979 and not w11991;
w11993 <= w11587 and not w11589;
w11994 <= not w11588 and w11993;
w11995 <= not w11591 and not w11994;
w11996 <= not w11992 and w11995;
w11997 <= w11992 and not w11995;
w11998 <= not w1299 and w11662;
w11999 <= not w1507 and w10990;
w12000 <= not w1407 and w11650;
w12001 <= not w11999 and not w12000;
w12002 <= not w11998 and w12001;
w12003 <= w5049 and w10992;
w12004 <= w12002 and not w12003;
w12005 <= not a(2) and not w12004;
w12006 <= a(2) and w12004;
w12007 <= not w12005 and not w12006;
w12008 <= not w11997 and not w12007;
w12009 <= not w11996 and not w12008;
w12010 <= w11722 and not w12009;
w12011 <= not w11722 and w12009;
w12012 <= not w1170 and w11662;
w12013 <= not w1407 and w10990;
w12014 <= not w1299 and w11650;
w12015 <= not w12013 and not w12014;
w12016 <= not w12012 and w12015;
w12017 <= w4783 and w10992;
w12018 <= w12016 and not w12017;
w12019 <= not a(2) and not w12018;
w12020 <= a(2) and w12018;
w12021 <= not w12019 and not w12020;
w12022 <= not w12011 and not w12021;
w12023 <= not w12010 and not w12022;
w12024 <= not w1113 and w11662;
w12025 <= not w1299 and w10990;
w12026 <= not w1170 and w11650;
w12027 <= not w12025 and not w12026;
w12028 <= not w12024 and w12027;
w12029 <= not w10992 and w12028;
w12030 <= not w4796 and w12028;
w12031 <= not w12029 and not w12030;
w12032 <= a(2) and not w12031;
w12033 <= not a(2) and w12031;
w12034 <= not w12032 and not w12033;
w12035 <= w12023 and w12034;
w12036 <= w11309 and w11596;
w12037 <= not w11597 and not w12036;
w12038 <= not w12035 and w12037;
w12039 <= not w12023 and not w12034;
w12040 <= not w12038 and not w12039;
w12041 <= not w995 and w11662;
w12042 <= not w1170 and w10990;
w12043 <= not w1113 and w11650;
w12044 <= not w12042 and not w12043;
w12045 <= not w12041 and w12044;
w12046 <= not w10992 and w12045;
w12047 <= not w4364 and w12045;
w12048 <= not w12046 and not w12047;
w12049 <= a(2) and not w12048;
w12050 <= not a(2) and w12048;
w12051 <= not w12049 and not w12050;
w12052 <= w12040 and w12051;
w12053 <= w11291 and w11598;
w12054 <= not w11599 and not w12053;
w12055 <= not w12052 and w12054;
w12056 <= not w12040 and not w12051;
w12057 <= not w12055 and not w12056;
w12058 <= not w893 and w11662;
w12059 <= not w1113 and w10990;
w12060 <= not w995 and w11650;
w12061 <= not w12059 and not w12060;
w12062 <= not w12058 and w12061;
w12063 <= not w10992 and w12062;
w12064 <= not w4568 and w12062;
w12065 <= not w12063 and not w12064;
w12066 <= a(2) and not w12065;
w12067 <= not a(2) and w12065;
w12068 <= not w12066 and not w12067;
w12069 <= w12057 and w12068;
w12070 <= w11273 and w11600;
w12071 <= not w11601 and not w12070;
w12072 <= not w12069 and w12071;
w12073 <= not w12057 and not w12068;
w12074 <= not w12072 and not w12073;
w12075 <= w11602 and not w11604;
w12076 <= not w11603 and w12075;
w12077 <= not w11606 and not w12076;
w12078 <= not w12074 and w12077;
w12079 <= w12074 and not w12077;
w12080 <= not w802 and w11662;
w12081 <= not w995 and w10990;
w12082 <= not w893 and w11650;
w12083 <= not w12081 and not w12082;
w12084 <= not w12080 and w12083;
w12085 <= w4139 and w10992;
w12086 <= w12084 and not w12085;
w12087 <= not a(2) and not w12086;
w12088 <= a(2) and w12086;
w12089 <= not w12087 and not w12088;
w12090 <= not w12079 and not w12089;
w12091 <= not w12078 and not w12090;
w12092 <= w11607 and not w11609;
w12093 <= not w11608 and w12092;
w12094 <= not w11611 and not w12093;
w12095 <= not w12091 and w12094;
w12096 <= w12091 and not w12094;
w12097 <= not w645 and w11662;
w12098 <= not w893 and w10990;
w12099 <= not w802 and w11650;
w12100 <= not w12098 and not w12099;
w12101 <= not w12097 and w12100;
w12102 <= w4114 and w10992;
w12103 <= w12101 and not w12102;
w12104 <= not a(2) and not w12103;
w12105 <= a(2) and w12103;
w12106 <= not w12104 and not w12105;
w12107 <= not w12096 and not w12106;
w12108 <= not w12095 and not w12107;
w12109 <= w11720 and not w12108;
w12110 <= not w11720 and w12108;
w12111 <= not w522 and w11662;
w12112 <= not w802 and w10990;
w12113 <= not w645 and w11650;
w12114 <= not w12112 and not w12113;
w12115 <= not w12111 and w12114;
w12116 <= w3266 and w10992;
w12117 <= w12115 and not w12116;
w12118 <= not a(2) and not w12117;
w12119 <= a(2) and w12117;
w12120 <= not w12118 and not w12119;
w12121 <= not w12110 and not w12120;
w12122 <= not w12109 and not w12121;
w12123 <= not w327 and w11662;
w12124 <= not w645 and w10990;
w12125 <= not w522 and w11650;
w12126 <= not w12124 and not w12125;
w12127 <= not w12123 and w12126;
w12128 <= not w10992 and w12127;
w12129 <= not w3282 and w12127;
w12130 <= not w12128 and not w12129;
w12131 <= a(2) and not w12130;
w12132 <= not a(2) and w12130;
w12133 <= not w12131 and not w12132;
w12134 <= w12122 and w12133;
w12135 <= w11214 and w11616;
w12136 <= not w11617 and not w12135;
w12137 <= not w12134 and w12136;
w12138 <= not w12122 and not w12133;
w12139 <= not w12137 and not w12138;
w12140 <= not w2947 and w11662;
w12141 <= not w522 and w10990;
w12142 <= not w327 and w11650;
w12143 <= not w12141 and not w12142;
w12144 <= not w12140 and w12143;
w12145 <= not w10992 and w12144;
w12146 <= not w2953 and w12144;
w12147 <= not w12145 and not w12146;
w12148 <= a(2) and not w12147;
w12149 <= not a(2) and w12147;
w12150 <= not w12148 and not w12149;
w12151 <= w12139 and w12150;
w12152 <= w11196 and w11618;
w12153 <= not w11619 and not w12152;
w12154 <= not w12151 and w12153;
w12155 <= not w12139 and not w12150;
w12156 <= not w12154 and not w12155;
w12157 <= not w3474 and w11662;
w12158 <= not w327 and w10990;
w12159 <= not w2947 and w11650;
w12160 <= not w12158 and not w12159;
w12161 <= not w12157 and w12160;
w12162 <= not w10992 and w12161;
w12163 <= not w3650 and w12161;
w12164 <= not w12162 and not w12163;
w12165 <= a(2) and not w12164;
w12166 <= not a(2) and w12164;
w12167 <= not w12165 and not w12166;
w12168 <= w12156 and w12167;
w12169 <= w11178 and w11620;
w12170 <= not w11621 and not w12169;
w12171 <= not w12168 and w12170;
w12172 <= not w12156 and not w12167;
w12173 <= not w12171 and not w12172;
w12174 <= w11622 and not w11624;
w12175 <= not w11623 and w12174;
w12176 <= not w11626 and not w12175;
w12177 <= not w12173 and w12176;
w12178 <= w12173 and not w12176;
w12179 <= not w3540 and w11662;
w12180 <= not w2947 and w10990;
w12181 <= not w3474 and w11650;
w12182 <= not w12180 and not w12181;
w12183 <= not w12179 and w12182;
w12184 <= w4019 and w10992;
w12185 <= w12183 and not w12184;
w12186 <= not a(2) and not w12185;
w12187 <= a(2) and w12185;
w12188 <= not w12186 and not w12187;
w12189 <= not w12178 and not w12188;
w12190 <= not w12177 and not w12189;
w12191 <= w11718 and not w12190;
w12192 <= not w11718 and w12190;
w12193 <= not w3391 and w11662;
w12194 <= not w3474 and w10990;
w12195 <= not w3540 and w11650;
w12196 <= not w12194 and not w12195;
w12197 <= not w12193 and w12196;
w12198 <= w3562 and w10992;
w12199 <= w12197 and not w12198;
w12200 <= not a(2) and not w12199;
w12201 <= a(2) and w12199;
w12202 <= not w12200 and not w12201;
w12203 <= not w12192 and not w12202;
w12204 <= not w12191 and not w12203;
w12205 <= not w3740 and w11662;
w12206 <= not w3540 and w10990;
w12207 <= not w3391 and w11650;
w12208 <= not w12206 and not w12207;
w12209 <= not w12205 and w12208;
w12210 <= not w10992 and w12209;
w12211 <= not w3753 and w12209;
w12212 <= not w12210 and not w12211;
w12213 <= a(2) and not w12212;
w12214 <= not a(2) and w12212;
w12215 <= not w12213 and not w12214;
w12216 <= w12204 and w12215;
w12217 <= w11133 and w11631;
w12218 <= not w11632 and not w12217;
w12219 <= not w12216 and w12218;
w12220 <= not w12204 and not w12215;
w12221 <= not w12219 and not w12220;
w12222 <= w11704 and not w11716;
w12223 <= not w11715 and not w11716;
w12224 <= not w12222 and not w12223;
w12225 <= not w12221 and not w12224;
w12226 <= not w11716 and not w12225;
w12227 <= not w11690 and w11701;
w12228 <= not w11702 and not w12227;
w12229 <= not w12226 and w12228;
w12230 <= not w11702 and not w12229;
w12231 <= not w11676 and w11687;
w12232 <= not w11688 and not w12231;
w12233 <= not w12230 and w12232;
w12234 <= not w11688 and not w12233;
w12235 <= not w11661 and w11673;
w12236 <= not w11674 and not w12235;
w12237 <= not w12234 and w12236;
w12238 <= not w11674 and not w12237;
w12239 <= not w11648 and w11658;
w12240 <= not w11659 and not w12239;
w12241 <= not w12238 and w12240;
w12242 <= not w11659 and not w12241;
w12243 <= w11646 and not w12242;
w12244 <= not w11644 and not w12243;
w12245 <= w11018 and not w11021;
w12246 <= not w11022 and not w12245;
w12247 <= not w12244 and w12246;
w12248 <= not w11022 and not w12247;
w12249 <= w10982 and not w10984;
w12250 <= not w10985 and not w12249;
w12251 <= not w12248 and w12250;
w12252 <= not w10985 and not w12251;
w12253 <= w10388 and not w12252;
w12254 <= not w10386 and not w12253;
w12255 <= w9818 and not w9821;
w12256 <= not w9822 and not w12255;
w12257 <= not w12254 and w12256;
w12258 <= not w9822 and not w12257;
w12259 <= w9298 and not w9300;
w12260 <= not w9301 and not w12259;
w12261 <= not w12258 and w12260;
w12262 <= not w9301 and not w12261;
w12263 <= w8814 and not w12262;
w12264 <= not w8812 and not w12263;
w12265 <= w8372 and not w12264;
w12266 <= not w8370 and not w12265;
w12267 <= w7950 and not w7952;
w12268 <= not w7953 and not w12267;
w12269 <= not w12266 and w12268;
w12270 <= not w7953 and not w12269;
w12271 <= w7586 and not w12270;
w12272 <= not w7584 and not w12271;
w12273 <= w7242 and not w7245;
w12274 <= not w7246 and not w12273;
w12275 <= not w12272 and w12274;
w12276 <= not w7246 and not w12275;
w12277 <= w7068 and not w7070;
w12278 <= not w7071 and not w12277;
w12279 <= not w12276 and w12278;
w12280 <= not w7071 and not w12279;
w12281 <= w6905 and not w12280;
w12282 <= not w6903 and not w12281;
w12283 <= w6357 and not w12282;
w12284 <= not w6355 and not w12283;
w12285 <= w6202 and not w12284;
w12286 <= not w6200 and not w12285;
w12287 <= w5887 and not w12286;
w12288 <= not w5885 and not w12287;
w12289 <= w5614 and not w5616;
w12290 <= not w5617 and not w12289;
w12291 <= not w12288 and w12290;
w12292 <= not w5617 and not w12291;
w12293 <= w5465 and not w12292;
w12294 <= not w5463 and not w12293;
w12295 <= w5355 and not w12294;
w12296 <= not w5353 and not w12295;
w12297 <= w4889 and not w12296;
w12298 <= not w4887 and not w12297;
w12299 <= w4663 and not w4665;
w12300 <= not w4666 and not w12299;
w12301 <= not w12298 and w12300;
w12302 <= not w4666 and not w12301;
w12303 <= w4557 and not w12302;
w12304 <= not w4557 and w12302;
w12305 <= not w12303 and not w12304;
w12306 <= not w4556 and not w12303;
w12307 <= not w4477 and not w4480;
w12308 <= w3392 and not w3899;
w12309 <= not w3391 and w3477;
w12310 <= w3541 and not w3740;
w12311 <= not w12309 and not w12310;
w12312 <= not w12308 and w12311;
w12313 <= w3303 and w4493;
w12314 <= w12312 and not w12313;
w12315 <= a(29) and not w12314;
w12316 <= a(29) and not w12315;
w12317 <= not w12314 and not w12315;
w12318 <= not w12316 and not w12317;
w12319 <= not w3655 and not w3659;
w12320 <= w223 and w2211;
w12321 <= not w58 and w12320;
w12322 <= not w166 and w12321;
w12323 <= not w430 and w443;
w12324 <= not w302 and w12323;
w12325 <= not w140 and w12324;
w12326 <= w2519 and w12325;
w12327 <= w12322 and w12326;
w12328 <= w2517 and w12327;
w12329 <= not w106 and w12328;
w12330 <= not w56 and w12329;
w12331 <= not w98 and w12330;
w12332 <= not w335 and not w1138;
w12333 <= w1485 and w12332;
w12334 <= not w46 and w12333;
w12335 <= not w224 and w12334;
w12336 <= not w361 and w12335;
w12337 <= not w867 and w12336;
w12338 <= not w405 and w12337;
w12339 <= not w206 and w12338;
w12340 <= w468 and w1006;
w12341 <= not w129 and w12340;
w12342 <= not w138 and w12341;
w12343 <= not w82 and w12342;
w12344 <= not w338 and w12343;
w12345 <= not w225 and w2281;
w12346 <= not w387 and w12345;
w12347 <= not w241 and w12346;
w12348 <= w1579 and w12347;
w12349 <= w12344 and w12348;
w12350 <= w1431 and w12349;
w12351 <= w2896 and w12350;
w12352 <= w746 and w12351;
w12353 <= w709 and w12352;
w12354 <= w1188 and w12353;
w12355 <= w1929 and w12354;
w12356 <= w820 and w12355;
w12357 <= not w211 and w12356;
w12358 <= not w782 and w12357;
w12359 <= not w290 and w12358;
w12360 <= not w26 and w12359;
w12361 <= not w359 and w12360;
w12362 <= not w386 and w12361;
w12363 <= not w16 and w12362;
w12364 <= not w77 and not w236;
w12365 <= not w499 and w12364;
w12366 <= not w568 and w12365;
w12367 <= w188 and w657;
w12368 <= w1093 and w12367;
w12369 <= w12366 and w12368;
w12370 <= w12363 and w12369;
w12371 <= w12339 and w12370;
w12372 <= w6704 and w12371;
w12373 <= w12331 and w12372;
w12374 <= w3098 and w12373;
w12375 <= not w1241 and w12374;
w12376 <= not w167 and w12375;
w12377 <= not w506 and w12376;
w12378 <= not w591 and w12377;
w12379 <= not w292 and w12378;
w12380 <= not w306 and w12379;
w12381 <= not w54 and w12380;
w12382 <= not w504 and w12381;
w12383 <= not w364 and w12382;
w12384 <= not w3637 and not w12383;
w12385 <= w3637 and w12383;
w12386 <= not w12384 and not w12385;
w12387 <= not a(23) and w12386;
w12388 <= not a(23) and not w12387;
w12389 <= not w12384 and not w12387;
w12390 <= not w12385 and w12389;
w12391 <= not w12388 and not w12390;
w12392 <= w2955 and not w3540;
w12393 <= w2963 and not w3474;
w12394 <= not w2947 and w2958;
w12395 <= w10 and w4019;
w12396 <= not w12394 and not w12395;
w12397 <= not w12393 and w12396;
w12398 <= not w12392 and w12397;
w12399 <= not w12391 and not w12398;
w12400 <= w12391 and w12398;
w12401 <= not w12399 and not w12400;
w12402 <= not w3643 and w12401;
w12403 <= w3643 and not w12401;
w12404 <= not w12402 and not w12403;
w12405 <= not w12319 and w12404;
w12406 <= w12319 and not w12404;
w12407 <= not w12405 and not w12406;
w12408 <= not w12318 and w12407;
w12409 <= w12407 and not w12408;
w12410 <= not w12318 and not w12408;
w12411 <= not w12409 and not w12410;
w12412 <= not w3760 and not w4009;
w12413 <= w3819 and not w4450;
w12414 <= w3902 and not w3980;
w12415 <= not w3812 and w3981;
w12416 <= not w12414 and not w12415;
w12417 <= not w12413 and w12416;
w12418 <= not w3985 and w12417;
w12419 <= not w4650 and w12417;
w12420 <= not w12418 and not w12419;
w12421 <= a(26) and not w12420;
w12422 <= not a(26) and w12420;
w12423 <= not w12421 and not w12422;
w12424 <= not w12412 and not w12423;
w12425 <= not w12412 and not w12424;
w12426 <= not w12423 and not w12424;
w12427 <= not w12425 and not w12426;
w12428 <= not w12411 and not w12427;
w12429 <= w12411 and not w12426;
w12430 <= not w12425 and w12429;
w12431 <= not w12428 and not w12430;
w12432 <= not w12307 and w12431;
w12433 <= w12307 and not w12431;
w12434 <= not w12432 and not w12433;
w12435 <= not w12306 and w12434;
w12436 <= w12306 and not w12434;
w12437 <= not w12435 and not w12436;
w12438 <= w12305 and w12437;
w12439 <= w12298 and not w12300;
w12440 <= not w12301 and not w12439;
w12441 <= w12305 and w12440;
w12442 <= not w4889 and w12296;
w12443 <= not w12297 and not w12442;
w12444 <= w12440 and w12443;
w12445 <= not w5465 and w12292;
w12446 <= not w12293 and not w12445;
w12447 <= not w5355 and w12294;
w12448 <= not w12295 and not w12447;
w12449 <= w12446 and w12448;
w12450 <= w12288 and not w12290;
w12451 <= not w12291 and not w12450;
w12452 <= w12446 and w12451;
w12453 <= not w5887 and w12286;
w12454 <= not w12287 and not w12453;
w12455 <= w12451 and w12454;
w12456 <= not w6202 and w12284;
w12457 <= not w12285 and not w12456;
w12458 <= w12454 and w12457;
w12459 <= not w6357 and w12282;
w12460 <= not w12283 and not w12459;
w12461 <= w12457 and w12460;
w12462 <= not w6905 and w12280;
w12463 <= not w12281 and not w12462;
w12464 <= w12460 and w12463;
w12465 <= w12276 and not w12278;
w12466 <= not w12279 and not w12465;
w12467 <= w12463 and w12466;
w12468 <= w12272 and not w12274;
w12469 <= not w12275 and not w12468;
w12470 <= w12466 and w12469;
w12471 <= not w7586 and w12270;
w12472 <= not w12271 and not w12471;
w12473 <= w12469 and w12472;
w12474 <= w12266 and not w12268;
w12475 <= not w12269 and not w12474;
w12476 <= w12472 and w12475;
w12477 <= not w8372 and w12264;
w12478 <= not w12265 and not w12477;
w12479 <= w12475 and w12478;
w12480 <= not w8814 and w12262;
w12481 <= not w12263 and not w12480;
w12482 <= w12478 and w12481;
w12483 <= w12258 and not w12260;
w12484 <= not w12261 and not w12483;
w12485 <= w12481 and w12484;
w12486 <= w12254 and not w12256;
w12487 <= not w12257 and not w12486;
w12488 <= w12484 and w12487;
w12489 <= not w10388 and w12252;
w12490 <= not w12253 and not w12489;
w12491 <= w12487 and w12490;
w12492 <= w12248 and not w12250;
w12493 <= not w12251 and not w12492;
w12494 <= w12490 and w12493;
w12495 <= w12244 and not w12246;
w12496 <= not w12247 and not w12495;
w12497 <= w12493 and w12496;
w12498 <= not w11646 and w12242;
w12499 <= not w12243 and not w12498;
w12500 <= w12496 and w12499;
w12501 <= w12238 and not w12240;
w12502 <= not w12241 and not w12501;
w12503 <= w12499 and w12502;
w12504 <= not w12499 and not w12502;
w12505 <= w12234 and not w12236;
w12506 <= not w12237 and not w12505;
w12507 <= w12502 and w12506;
w12508 <= w12230 and not w12232;
w12509 <= not w12233 and not w12508;
w12510 <= w12506 and w12509;
w12511 <= w12226 and not w12228;
w12512 <= not w12229 and not w12511;
w12513 <= w12509 and w12512;
w12514 <= not w12221 and not w12225;
w12515 <= not w12224 and not w12225;
w12516 <= not w12514 and not w12515;
w12517 <= w12512 and not w12516;
w12518 <= not w12509 and w12517;
w12519 <= not w12513 and not w12518;
w12520 <= not w12506 and not w12509;
w12521 <= not w12510 and not w12520;
w12522 <= not w12519 and w12521;
w12523 <= not w12510 and not w12522;
w12524 <= not w12502 and not w12506;
w12525 <= not w12507 and not w12524;
w12526 <= not w12523 and w12525;
w12527 <= not w12507 and not w12526;
w12528 <= not w12503 and not w12527;
w12529 <= not w12504 and w12528;
w12530 <= not w12503 and not w12529;
w12531 <= not w12496 and not w12499;
w12532 <= not w12530 and not w12531;
w12533 <= not w12500 and w12532;
w12534 <= not w12500 and not w12533;
w12535 <= not w12493 and not w12496;
w12536 <= not w12497 and not w12535;
w12537 <= not w12534 and w12536;
w12538 <= not w12497 and not w12537;
w12539 <= not w12490 and not w12493;
w12540 <= not w12538 and not w12539;
w12541 <= not w12494 and w12540;
w12542 <= not w12494 and not w12541;
w12543 <= not w12487 and not w12490;
w12544 <= not w12542 and not w12543;
w12545 <= not w12491 and w12544;
w12546 <= not w12491 and not w12545;
w12547 <= not w12484 and not w12487;
w12548 <= not w12488 and not w12547;
w12549 <= not w12546 and w12548;
w12550 <= not w12488 and not w12549;
w12551 <= not w12481 and not w12484;
w12552 <= not w12550 and not w12551;
w12553 <= not w12485 and w12552;
w12554 <= not w12485 and not w12553;
w12555 <= not w12478 and not w12481;
w12556 <= not w12482 and not w12555;
w12557 <= not w12554 and w12556;
w12558 <= not w12482 and not w12557;
w12559 <= not w12475 and not w12478;
w12560 <= not w12558 and not w12559;
w12561 <= not w12479 and w12560;
w12562 <= not w12479 and not w12561;
w12563 <= not w12472 and not w12475;
w12564 <= not w12562 and not w12563;
w12565 <= not w12476 and w12564;
w12566 <= not w12476 and not w12565;
w12567 <= not w12469 and not w12472;
w12568 <= not w12566 and not w12567;
w12569 <= not w12473 and w12568;
w12570 <= not w12473 and not w12569;
w12571 <= not w12466 and not w12469;
w12572 <= not w12470 and not w12571;
w12573 <= not w12570 and w12572;
w12574 <= not w12470 and not w12573;
w12575 <= not w12463 and not w12466;
w12576 <= not w12574 and not w12575;
w12577 <= not w12467 and w12576;
w12578 <= not w12467 and not w12577;
w12579 <= not w12460 and not w12463;
w12580 <= not w12464 and not w12579;
w12581 <= not w12578 and w12580;
w12582 <= not w12464 and not w12581;
w12583 <= not w12457 and not w12460;
w12584 <= not w12461 and not w12583;
w12585 <= not w12582 and w12584;
w12586 <= not w12461 and not w12585;
w12587 <= not w12454 and not w12457;
w12588 <= not w12458 and not w12587;
w12589 <= not w12586 and w12588;
w12590 <= not w12458 and not w12589;
w12591 <= not w12451 and not w12454;
w12592 <= not w12590 and not w12591;
w12593 <= not w12455 and w12592;
w12594 <= not w12455 and not w12593;
w12595 <= not w12446 and not w12451;
w12596 <= not w12594 and not w12595;
w12597 <= not w12452 and w12596;
w12598 <= not w12452 and not w12597;
w12599 <= not w12446 and not w12448;
w12600 <= not w12449 and not w12599;
w12601 <= not w12598 and w12600;
w12602 <= not w12449 and not w12601;
w12603 <= not w12443 and not w12448;
w12604 <= w12443 and w12448;
w12605 <= not w12603 and not w12604;
w12606 <= not w12602 and w12605;
w12607 <= not w12604 and not w12606;
w12608 <= not w12440 and not w12443;
w12609 <= not w12607 and not w12608;
w12610 <= not w12444 and w12609;
w12611 <= not w12444 and not w12610;
w12612 <= not w12305 and not w12440;
w12613 <= not w12611 and not w12612;
w12614 <= not w12441 and w12613;
w12615 <= not w12441 and not w12614;
w12616 <= not w12305 and not w12437;
w12617 <= not w12615 and not w12616;
w12618 <= not w12438 and w12617;
w12619 <= not w12438 and not w12618;
w12620 <= not w12432 and not w12435;
w12621 <= not w12424 and not w12428;
w12622 <= not w3812 and w3902;
w12623 <= w3981 and not w4450;
w12624 <= not w12622 and not w12623;
w12625 <= w3985 and w4544;
w12626 <= w12624 and not w12625;
w12627 <= a(26) and not w12626;
w12628 <= not w12626 and not w12627;
w12629 <= a(26) and not w12627;
w12630 <= not w12628 and not w12629;
w12631 <= not w12405 and not w12408;
w12632 <= w10 and w3562;
w12633 <= w2955 and not w3391;
w12634 <= w2958 and not w3474;
w12635 <= w2963 and not w3540;
w12636 <= not w12634 and not w12635;
w12637 <= not w12633 and w12636;
w12638 <= not w12632 and w12637;
w12639 <= not w104 and not w129;
w12640 <= not w738 and w12639;
w12641 <= not w1036 and w12640;
w12642 <= not w354 and w12641;
w12643 <= not w329 and w12642;
w12644 <= not w592 and w12643;
w12645 <= not w96 and w12644;
w12646 <= not w167 and not w328;
w12647 <= not w136 and w12646;
w12648 <= w2296 and w12647;
w12649 <= w1814 and w12648;
w12650 <= w5989 and w12649;
w12651 <= w5741 and w12650;
w12652 <= w1484 and w12651;
w12653 <= w2442 and w12652;
w12654 <= w1512 and w12653;
w12655 <= w2508 and w12654;
w12656 <= w12645 and w12655;
w12657 <= w55 and w12656;
w12658 <= w4721 and w12657;
w12659 <= w291 and w12658;
w12660 <= w51 and w12659;
w12661 <= not w89 and w12660;
w12662 <= not w650 and w12661;
w12663 <= not w37 and w12662;
w12664 <= not w212 and w12663;
w12665 <= not w205 and w12664;
w12666 <= not w12389 and w12665;
w12667 <= w12389 and not w12665;
w12668 <= not w12666 and not w12667;
w12669 <= not w12638 and w12668;
w12670 <= not w12638 and not w12669;
w12671 <= w12668 and not w12669;
w12672 <= not w12670 and not w12671;
w12673 <= not w12399 and not w12402;
w12674 <= w12672 and w12673;
w12675 <= not w12672 and not w12673;
w12676 <= not w12674 and not w12675;
w12677 <= w3392 and not w3980;
w12678 <= w3477 and not w3740;
w12679 <= w3541 and not w3899;
w12680 <= not w12678 and not w12679;
w12681 <= not w12677 and w12680;
w12682 <= not w3303 and w12681;
w12683 <= not w4412 and w12681;
w12684 <= not w12682 and not w12683;
w12685 <= a(29) and not w12684;
w12686 <= not a(29) and w12684;
w12687 <= not w12685 and not w12686;
w12688 <= w12676 and not w12687;
w12689 <= not w12676 and w12687;
w12690 <= not w12688 and not w12689;
w12691 <= not w12631 and w12690;
w12692 <= not w12631 and not w12691;
w12693 <= w12690 and not w12691;
w12694 <= not w12692 and not w12693;
w12695 <= not w12630 and not w12694;
w12696 <= w12630 and not w12693;
w12697 <= not w12692 and w12696;
w12698 <= not w12695 and not w12697;
w12699 <= not w12621 and w12698;
w12700 <= w12621 and not w12698;
w12701 <= not w12699 and not w12700;
w12702 <= not w12620 and w12701;
w12703 <= w12620 and not w12701;
w12704 <= not w12702 and not w12703;
w12705 <= not w12437 and not w12704;
w12706 <= w12437 and w12704;
w12707 <= not w12705 and not w12706;
w12708 <= not w12619 and w12707;
w12709 <= not w12706 and not w12708;
w12710 <= not w12699 and not w12702;
w12711 <= not w12691 and not w12695;
w12712 <= w10 and w3753;
w12713 <= w2955 and not w3740;
w12714 <= w2958 and not w3540;
w12715 <= w2963 and not w3391;
w12716 <= not w12714 and not w12715;
w12717 <= not w12713 and w12716;
w12718 <= not w12712 and w12717;
w12719 <= not w159 and not w240;
w12720 <= not w649 and w12719;
w12721 <= w588 and w12720;
w12722 <= w2508 and w12721;
w12723 <= w2517 and w12722;
w12724 <= not w211 and w12723;
w12725 <= not w395 and w12724;
w12726 <= not w867 and w12725;
w12727 <= not w208 and w12726;
w12728 <= not w160 and w12727;
w12729 <= not w647 and w12728;
w12730 <= not w166 and w12729;
w12731 <= w496 and w5743;
w12732 <= w1411 and w12731;
w12733 <= w903 and w12732;
w12734 <= w2105 and w12733;
w12735 <= w217 and w12734;
w12736 <= w1182 and w12735;
w12737 <= not w141 and w12736;
w12738 <= not w608 and w12737;
w12739 <= not w466 and w12738;
w12740 <= not w1039 and w12739;
w12741 <= not w397 and not w602;
w12742 <= not w86 and w12741;
w12743 <= not w997 and w12742;
w12744 <= not w386 and w12743;
w12745 <= not w60 and w12744;
w12746 <= not w338 and not w441;
w12747 <= not w536 and w12746;
w12748 <= w1462 and w12747;
w12749 <= w12745 and w12748;
w12750 <= w12740 and w12749;
w12751 <= w4729 and w12750;
w12752 <= w137 and w12751;
w12753 <= not w125 and w12752;
w12754 <= not w190 and w12753;
w12755 <= not w174 and w12754;
w12756 <= not w56 and w12755;
w12757 <= not w337 and w12756;
w12758 <= not w222 and w12757;
w12759 <= not w237 and w12758;
w12760 <= not w178 and w12759;
w12761 <= not w454 and w12760;
w12762 <= not w206 and w12761;
w12763 <= not w364 and w12762;
w12764 <= not w269 and not w370;
w12765 <= not w187 and w12764;
w12766 <= w3762 and w12765;
w12767 <= w6019 and w12766;
w12768 <= w12763 and w12767;
w12769 <= w12730 and w12768;
w12770 <= w1414 and w12769;
w12771 <= w94 and w12770;
w12772 <= w1602 and w12771;
w12773 <= w505 and w12772;
w12774 <= not w219 and w12773;
w12775 <= not w126 and w12774;
w12776 <= not w387 and w12775;
w12777 <= not w409 and w12776;
w12778 <= not w12665 and w12777;
w12779 <= w12665 and not w12777;
w12780 <= not w12718 and not w12779;
w12781 <= not w12778 and w12780;
w12782 <= not w12718 and not w12781;
w12783 <= not w12779 and not w12781;
w12784 <= not w12778 and w12783;
w12785 <= not w12782 and not w12784;
w12786 <= not w12666 and not w12669;
w12787 <= w12785 and w12786;
w12788 <= not w12785 and not w12786;
w12789 <= not w12787 and not w12788;
w12790 <= not w12675 and not w12688;
w12791 <= w12789 and not w12790;
w12792 <= not w12789 and w12790;
w12793 <= not w12791 and not w12792;
w12794 <= w3985 and w4457;
w12795 <= w3902 and not w4450;
w12796 <= not w12794 and not w12795;
w12797 <= a(26) and not w12796;
w12798 <= not w12796 and not w12797;
w12799 <= a(26) and not w12797;
w12800 <= not w12798 and not w12799;
w12801 <= w3392 and not w3812;
w12802 <= w3477 and not w3899;
w12803 <= w3541 and not w3980;
w12804 <= not w12802 and not w12803;
w12805 <= not w12801 and w12804;
w12806 <= w3303 and w4002;
w12807 <= w12805 and not w12806;
w12808 <= a(29) and not w12807;
w12809 <= a(29) and not w12808;
w12810 <= not w12807 and not w12808;
w12811 <= not w12809 and not w12810;
w12812 <= not w12800 and not w12811;
w12813 <= not w12800 and not w12812;
w12814 <= not w12811 and not w12812;
w12815 <= not w12813 and not w12814;
w12816 <= w12793 and not w12815;
w12817 <= not w12793 and w12815;
w12818 <= not w12816 and not w12817;
w12819 <= not w12711 and w12818;
w12820 <= w12711 and not w12818;
w12821 <= not w12819 and not w12820;
w12822 <= not w12710 and w12821;
w12823 <= w12710 and not w12821;
w12824 <= not w12822 and not w12823;
w12825 <= not w12704 and not w12824;
w12826 <= w12704 and w12824;
w12827 <= not w12825 and not w12826;
w12828 <= not w12709 and w12827;
w12829 <= w12709 and not w12827;
w12830 <= not w12828 and not w12829;
w12831 <= w10 and w12830;
w12832 <= w2955 and w12824;
w12833 <= w2958 and w12437;
w12834 <= w2963 and w12704;
w12835 <= not w12833 and not w12834;
w12836 <= not w12832 and w12835;
w12837 <= not w12831 and w12836;
w12838 <= not w211 and not w602;
w12839 <= not w125 and w12838;
w12840 <= not w1036 and w12839;
w12841 <= not w331 and w12840;
w12842 <= not w388 and w12841;
w12843 <= not w357 and w12842;
w12844 <= not w67 and w12843;
w12845 <= w165 and not w241;
w12846 <= not w207 and w12845;
w12847 <= w1546 and w4262;
w12848 <= w12846 and w12847;
w12849 <= not w90 and w12848;
w12850 <= not w337 and w12849;
w12851 <= not w1039 and w12850;
w12852 <= not w818 and w12851;
w12853 <= not w272 and w12852;
w12854 <= not w123 and w12853;
w12855 <= not w174 and w2027;
w12856 <= not w760 and w12855;
w12857 <= not w536 and w12856;
w12858 <= not w502 and w12857;
w12859 <= not w228 and w12858;
w12860 <= w1929 and w6455;
w12861 <= w1717 and w12860;
w12862 <= not w46 and w12861;
w12863 <= not w177 and w12862;
w12864 <= not w262 and w12863;
w12865 <= not w82 and w12864;
w12866 <= not w330 and w12865;
w12867 <= not w21 and w12866;
w12868 <= w575 and w4975;
w12869 <= w12867 and w12868;
w12870 <= w12859 and w12869;
w12871 <= w2378 and w12870;
w12872 <= not w71 and w12871;
w12873 <= not w821 and w12872;
w12874 <= not w293 and w12873;
w12875 <= not w290 and not w946;
w12876 <= not w106 and w12875;
w12877 <= w308 and w12876;
w12878 <= w1172 and w12877;
w12879 <= not w499 and w12878;
w12880 <= w573 and w2165;
w12881 <= w1184 and w12880;
w12882 <= w2403 and w12881;
w12883 <= w12879 and w12882;
w12884 <= w12874 and w12883;
w12885 <= w2558 and w12884;
w12886 <= w12854 and w12885;
w12887 <= w12844 and w12886;
w12888 <= w1064 and w12887;
w12889 <= w4230 and w12888;
w12890 <= not w265 and w12889;
w12891 <= not w189 and w12890;
w12892 <= not w227 and w12891;
w12893 <= not w26 and w12892;
w12894 <= w2619 and w3373;
w12895 <= w465 and w12894;
w12896 <= w1860 and w12895;
w12897 <= w724 and w12896;
w12898 <= w1189 and w12897;
w12899 <= w1762 and w12898;
w12900 <= w1096 and w12899;
w12901 <= not w782 and w12900;
w12902 <= not w554 and w12901;
w12903 <= not w90 and w12902;
w12904 <= not w572 and w12903;
w12905 <= not w915 and w12904;
w12906 <= not w329 and w12905;
w12907 <= not w160 and w12906;
w12908 <= not w267 and w12907;
w12909 <= not w216 and not w361;
w12910 <= not w124 and w12909;
w12911 <= not w396 and w12910;
w12912 <= not w166 and w12911;
w12913 <= w3920 and w4269;
w12914 <= w12912 and w12913;
w12915 <= w1151 and w12914;
w12916 <= w5159 and w12915;
w12917 <= w1904 and w12916;
w12918 <= w12908 and w12917;
w12919 <= w1458 and w12918;
w12920 <= w2568 and w12919;
w12921 <= w1760 and w12920;
w12922 <= w1187 and w12921;
w12923 <= not w177 and w12922;
w12924 <= not w290 and w12923;
w12925 <= not w430 and w12924;
w12926 <= not w181 and w12925;
w12927 <= w6641 and w12926;
w12928 <= not w310 and w12927;
w12929 <= not w172 and w12928;
w12930 <= not w499 and w12929;
w12931 <= w12893 and not w12930;
w12932 <= not w12893 and w12930;
w12933 <= w12619 and not w12707;
w12934 <= not w12708 and not w12933;
w12935 <= w10 and w12934;
w12936 <= w2955 and w12704;
w12937 <= w2958 and w12305;
w12938 <= w2963 and w12437;
w12939 <= not w12937 and not w12938;
w12940 <= not w12936 and w12939;
w12941 <= not w12935 and w12940;
w12942 <= not w12931 and not w12941;
w12943 <= not w12932 and w12942;
w12944 <= not w12931 and not w12943;
w12945 <= not w104 and w173;
w12946 <= not w449 and w12945;
w12947 <= not w54 and w12946;
w12948 <= not w288 and not w782;
w12949 <= not w261 and w12948;
w12950 <= not w354 and not w624;
w12951 <= not w428 and w12950;
w12952 <= w12949 and w12951;
w12953 <= w1628 and w12952;
w12954 <= w12947 and w12953;
w12955 <= w12730 and w12954;
w12956 <= w1446 and w12955;
w12957 <= w2717 and w12956;
w12958 <= w2442 and w12957;
w12959 <= w1762 and w12958;
w12960 <= w1183 and w12959;
w12961 <= not w236 and w12960;
w12962 <= not w213 and w12961;
w12963 <= not w50 and w12962;
w12964 <= not w26 and w12963;
w12965 <= not w439 and w12964;
w12966 <= not w371 and w12965;
w12967 <= w1491 and w4086;
w12968 <= w832 and w12967;
w12969 <= w526 and w12968;
w12970 <= not w591 and w12969;
w12971 <= not w529 and w12970;
w12972 <= not w352 and w12971;
w12973 <= not w462 and w12972;
w12974 <= not w100 and w12973;
w12975 <= not w607 and w12974;
w12976 <= not w228 and w12975;
w12977 <= w1955 and w6599;
w12978 <= w528 and w12977;
w12979 <= w6542 and w12978;
w12980 <= w12763 and w12979;
w12981 <= w12976 and w12980;
w12982 <= w1456 and w12981;
w12983 <= w12966 and w12982;
w12984 <= w964 and w12983;
w12985 <= w226 and w12984;
w12986 <= w1074 and w12985;
w12987 <= w761 and w12986;
w12988 <= w1324 and w12987;
w12989 <= w276 and w12988;
w12990 <= not w1037 and w12989;
w12991 <= not w1062 and w12990;
w12992 <= w3766 and w12991;
w12993 <= w128 and w12992;
w12994 <= not w387 and w12993;
w12995 <= w1190 and w1716;
w12996 <= w3919 and w12995;
w12997 <= not w524 and w12996;
w12998 <= not w384 and w12997;
w12999 <= w2200 and w3841;
w13000 <= w3515 and w12999;
w13001 <= w5168 and w13000;
w13002 <= w3952 and w13001;
w13003 <= w12998 and w13002;
w13004 <= w4437 and w13003;
w13005 <= w3783 and w13004;
w13006 <= w2673 and w13005;
w13007 <= w2518 and w13006;
w13008 <= not w177 and w13007;
w13009 <= not w453 and w13008;
w13010 <= w3504 and w3841;
w13011 <= w3767 and w3969;
w13012 <= w13010 and w13011;
w13013 <= w3804 and w13012;
w13014 <= not w263 and w13013;
w13015 <= not w471 and w13014;
w13016 <= not w502 and w13015;
w13017 <= w13009 and w13016;
w13018 <= not w12994 and w13017;
w13019 <= w3505 and w3767;
w13020 <= w474 and w13019;
w13021 <= w903 and w13020;
w13022 <= not w388 and w13021;
w13023 <= w3884 and w13022;
w13024 <= w3791 and w13023;
w13025 <= w4428 and w13024;
w13026 <= w600 and w13025;
w13027 <= w1696 and w13026;
w13028 <= not w536 and w13027;
w13029 <= not w608 and w13028;
w13030 <= not w34 and w13029;
w13031 <= w13009 and not w13030;
w13032 <= not w13009 and w13030;
w13033 <= w10 and w4457;
w13034 <= w2958 and not w4450;
w13035 <= not w13033 and not w13034;
w13036 <= not w13031 and not w13035;
w13037 <= not w13032 and w13036;
w13038 <= not w13031 and not w13037;
w13039 <= not w13009 and not w13016;
w13040 <= not w13017 and not w13039;
w13041 <= not w13038 and not w13040;
w13042 <= not w13038 and not w13041;
w13043 <= not w13040 and not w13041;
w13044 <= not w13042 and not w13043;
w13045 <= not w13035 and not w13037;
w13046 <= not w13032 and w13038;
w13047 <= not w13045 and not w13046;
w13048 <= not w218 and not w1241;
w13049 <= not w184 and w13048;
w13050 <= w12332 and w13049;
w13051 <= w4151 and w13050;
w13052 <= w1851 and w13051;
w13053 <= not w240 and w13052;
w13054 <= not w338 and w13053;
w13055 <= not w181 and w13054;
w13056 <= not w454 and w13055;
w13057 <= not w60 and w13056;
w13058 <= not w228 and w13057;
w13059 <= w465 and w3505;
w13060 <= w2675 and w13059;
w13061 <= not w167 and w13060;
w13062 <= not w224 and w13061;
w13063 <= not w84 and w13062;
w13064 <= not w161 and w13063;
w13065 <= not w425 and w13064;
w13066 <= not w431 and w13065;
w13067 <= not w92 and w13066;
w13068 <= not w558 and w13067;
w13069 <= not w21 and w13068;
w13070 <= not w706 and w13069;
w13071 <= not w102 and w13070;
w13072 <= not w100 and w13071;
w13073 <= not w93 and w13072;
w13074 <= w1098 and w2479;
w13075 <= w13073 and w13074;
w13076 <= w1670 and w13075;
w13077 <= w1137 and w13076;
w13078 <= w13058 and w13077;
w13079 <= w5020 and w13078;
w13080 <= w2570 and w13079;
w13081 <= w1301 and w13080;
w13082 <= w665 and w13081;
w13083 <= w1187 and w13082;
w13084 <= w2401 and w13083;
w13085 <= w913 and w13084;
w13086 <= not w58 and w13085;
w13087 <= not w782 and w13086;
w13088 <= not w219 and w13087;
w13089 <= not w302 and w13088;
w13090 <= not w227 and w13089;
w13091 <= not w209 and w13090;
w13092 <= not w460 and w13091;
w13093 <= not w607 and w13092;
w13094 <= w3864 and w4999;
w13095 <= w820 and w13094;
w13096 <= not w79 and w13095;
w13097 <= w1360 and w1675;
w13098 <= w1184 and w13097;
w13099 <= w13096 and w13098;
w13100 <= w13022 and w13099;
w13101 <= w3882 and w13100;
w13102 <= w12998 and w13101;
w13103 <= w3944 and w13102;
w13104 <= w981 and w13103;
w13105 <= not w502 and w13104;
w13106 <= not w460 and w13105;
w13107 <= not w228 and w13106;
w13108 <= not w13093 and not w13107;
w13109 <= w13093 and w13107;
w13110 <= not w13108 and not w13109;
w13111 <= not a(29) and w13110;
w13112 <= not w13108 and not w13111;
w13113 <= w13009 and not w13112;
w13114 <= w10 and w4544;
w13115 <= w2958 and not w3812;
w13116 <= w2963 and not w4450;
w13117 <= not w13115 and not w13116;
w13118 <= not w13114 and w13117;
w13119 <= not w13009 and w13112;
w13120 <= not w13113 and not w13119;
w13121 <= not w13118 and w13120;
w13122 <= not w13113 and not w13121;
w13123 <= not w13047 and not w13122;
w13124 <= w13047 and w13122;
w13125 <= not w13123 and not w13124;
w13126 <= not w13118 and not w13121;
w13127 <= w13120 and not w13121;
w13128 <= not w13126 and not w13127;
w13129 <= not a(29) and not w13111;
w13130 <= not w13109 and w13112;
w13131 <= not w13129 and not w13130;
w13132 <= w1073 and w3235;
w13133 <= w710 and w13132;
w13134 <= w223 and w13133;
w13135 <= w406 and w13134;
w13136 <= w1661 and w13135;
w13137 <= w975 and w13136;
w13138 <= not w687 and w13137;
w13139 <= not w289 and w13138;
w13140 <= not w337 and w13139;
w13141 <= not w440 and w13140;
w13142 <= not w401 and w13141;
w13143 <= not w896 and w13142;
w13144 <= not w267 and w13143;
w13145 <= not w30 and w13144;
w13146 <= w556 and w3394;
w13147 <= w761 and w13146;
w13148 <= not w648 and w13147;
w13149 <= not w86 and w13148;
w13150 <= not w263 and w13149;
w13151 <= not w352 and w13150;
w13152 <= not w302 and w13151;
w13153 <= not w26 and w13152;
w13154 <= not w67 and w13153;
w13155 <= not w135 and w13154;
w13156 <= not w590 and w13155;
w13157 <= w3050 and w5722;
w13158 <= w559 and w13157;
w13159 <= w429 and w13158;
w13160 <= w2922 and w13159;
w13161 <= w13156 and w13160;
w13162 <= w13145 and w13161;
w13163 <= w6642 and w13162;
w13164 <= w4167 and w13163;
w13165 <= w1189 and w13164;
w13166 <= w1466 and w13165;
w13167 <= not w159 and w13166;
w13168 <= not w650 and w13167;
w13169 <= not w503 and w13168;
w13170 <= not w427 and w13169;
w13171 <= not w439 and w13170;
w13172 <= not w388 and w13171;
w13173 <= not w105 and w13172;
w13174 <= w13093 and not w13173;
w13175 <= not w13093 and w13173;
w13176 <= w4732 and w12347;
w13177 <= w1761 and w13176;
w13178 <= w353 and w13177;
w13179 <= not w287 and w13178;
w13180 <= not w79 and w13179;
w13181 <= not w260 and w13180;
w13182 <= not w384 and w13181;
w13183 <= not w81 and not w648;
w13184 <= not w62 and w13183;
w13185 <= w626 and w13184;
w13186 <= w6019 and w13185;
w13187 <= w6018 and w13186;
w13188 <= w1227 and w13187;
w13189 <= w3479 and w13188;
w13190 <= w220 and w13189;
w13191 <= w1760 and w13190;
w13192 <= w1301 and w13191;
w13193 <= not w171 and w13192;
w13194 <= not w1241 and w13193;
w13195 <= not w1037 and w13194;
w13196 <= not w222 and w13195;
w13197 <= not w425 and w13196;
w13198 <= not w127 and w13197;
w13199 <= not w181 and w13198;
w13200 <= not w601 and w13199;
w13201 <= not w301 and w525;
w13202 <= not w60 and w13201;
w13203 <= not w363 and w13202;
w13204 <= w3580 and w6039;
w13205 <= w1492 and w13204;
w13206 <= w13203 and w13205;
w13207 <= w2707 and w13206;
w13208 <= w13200 and w13207;
w13209 <= w13182 and w13208;
w13210 <= w2025 and w13209;
w13211 <= w1265 and w13210;
w13212 <= w2341 and w13211;
w13213 <= w91 and w13212;
w13214 <= w214 and w13213;
w13215 <= not w167 and w13214;
w13216 <= not w262 and w13215;
w13217 <= not w80 and w13216;
w13218 <= not w100 and w13217;
w13219 <= not w12665 and not w13218;
w13220 <= w12665 and w13218;
w13221 <= not w13219 and not w13220;
w13222 <= not a(26) and w13221;
w13223 <= not w13219 and not w13222;
w13224 <= w13173 and not w13223;
w13225 <= w10 and w4412;
w13226 <= w2955 and not w3980;
w13227 <= w2958 and not w3740;
w13228 <= w2963 and not w3899;
w13229 <= not w13227 and not w13228;
w13230 <= not w13226 and w13229;
w13231 <= not w13225 and w13230;
w13232 <= not w13173 and w13223;
w13233 <= not w13224 and not w13232;
w13234 <= not w13231 and w13233;
w13235 <= not w13224 and not w13234;
w13236 <= not w13174 and not w13235;
w13237 <= not w13175 and w13236;
w13238 <= not w13174 and not w13237;
w13239 <= not w13131 and not w13238;
w13240 <= w10 and w4650;
w13241 <= w2955 and not w4450;
w13242 <= w2958 and not w3980;
w13243 <= w2963 and not w3812;
w13244 <= not w13242 and not w13243;
w13245 <= not w13241 and w13244;
w13246 <= not w13240 and w13245;
w13247 <= w13131 and w13238;
w13248 <= not w13239 and not w13247;
w13249 <= not w13246 and w13248;
w13250 <= not w13239 and not w13249;
w13251 <= not w13128 and not w13250;
w13252 <= w13128 and w13250;
w13253 <= not w13251 and not w13252;
w13254 <= w3477 and not w4450;
w13255 <= w3303 and w4457;
w13256 <= not w13254 and not w13255;
w13257 <= a(29) and not w13256;
w13258 <= not w13256 and not w13257;
w13259 <= a(29) and not w13257;
w13260 <= not w13258 and not w13259;
w13261 <= w10 and w4002;
w13262 <= w2955 and not w3812;
w13263 <= w2958 and not w3899;
w13264 <= w2963 and not w3980;
w13265 <= not w13263 and not w13264;
w13266 <= not w13262 and w13265;
w13267 <= not w13261 and w13266;
w13268 <= not w13260 and not w13267;
w13269 <= not w13260 and not w13268;
w13270 <= not w13267 and not w13268;
w13271 <= not w13269 and not w13270;
w13272 <= not w13235 and not w13237;
w13273 <= not w13175 and w13238;
w13274 <= not w13272 and not w13273;
w13275 <= not w13271 and not w13274;
w13276 <= not w13268 and not w13275;
w13277 <= w13246 and not w13248;
w13278 <= not w13249 and not w13277;
w13279 <= not w13276 and w13278;
w13280 <= not w13231 and not w13234;
w13281 <= w13233 and not w13234;
w13282 <= not w13280 and not w13281;
w13283 <= not a(26) and not w13222;
w13284 <= not w13220 and w13223;
w13285 <= not w13283 and not w13284;
w13286 <= not w12783 and not w13285;
w13287 <= w10 and w4493;
w13288 <= w2955 and not w3899;
w13289 <= w2958 and not w3391;
w13290 <= w2963 and not w3740;
w13291 <= not w13289 and not w13290;
w13292 <= not w13288 and w13291;
w13293 <= not w13287 and w13292;
w13294 <= w12783 and w13285;
w13295 <= not w13286 and not w13294;
w13296 <= not w13293 and w13295;
w13297 <= not w13286 and not w13296;
w13298 <= not w13282 and not w13297;
w13299 <= w13282 and w13297;
w13300 <= not w13298 and not w13299;
w13301 <= w3477 and not w3812;
w13302 <= w3541 and not w4450;
w13303 <= not w13301 and not w13302;
w13304 <= w3303 and w4544;
w13305 <= w13303 and not w13304;
w13306 <= a(29) and not w13305;
w13307 <= a(29) and not w13306;
w13308 <= not w13305 and not w13306;
w13309 <= not w13307 and not w13308;
w13310 <= w13300 and not w13309;
w13311 <= not w13298 and not w13310;
w13312 <= not w13271 and w13274;
w13313 <= w13271 and not w13274;
w13314 <= not w13312 and not w13313;
w13315 <= not w13311 and not w13314;
w13316 <= w13300 and not w13310;
w13317 <= not w13309 and not w13310;
w13318 <= not w13316 and not w13317;
w13319 <= not w12788 and not w12791;
w13320 <= not w13293 and not w13296;
w13321 <= w13295 and not w13296;
w13322 <= not w13320 and not w13321;
w13323 <= not w13319 and not w13322;
w13324 <= not w13319 and not w13323;
w13325 <= not w13322 and not w13323;
w13326 <= not w13324 and not w13325;
w13327 <= w3392 and not w4450;
w13328 <= w3477 and not w3980;
w13329 <= w3541 and not w3812;
w13330 <= not w13328 and not w13329;
w13331 <= not w13327 and w13330;
w13332 <= w3303 and w4650;
w13333 <= w13331 and not w13332;
w13334 <= a(29) and not w13333;
w13335 <= a(29) and not w13334;
w13336 <= not w13333 and not w13334;
w13337 <= not w13335 and not w13336;
w13338 <= not w13326 and not w13337;
w13339 <= not w13323 and not w13338;
w13340 <= not w13318 and not w13339;
w13341 <= w13318 and w13339;
w13342 <= not w13340 and not w13341;
w13343 <= not w13326 and not w13338;
w13344 <= not w13337 and not w13338;
w13345 <= not w13343 and not w13344;
w13346 <= not w12812 and not w12816;
w13347 <= not w13345 and not w13346;
w13348 <= not w13345 and not w13347;
w13349 <= not w13346 and not w13347;
w13350 <= not w13348 and not w13349;
w13351 <= not w12819 and not w12822;
w13352 <= not w13350 and not w13351;
w13353 <= not w13347 and not w13352;
w13354 <= w13342 and not w13353;
w13355 <= not w13340 and not w13354;
w13356 <= w13311 and w13314;
w13357 <= not w13315 and not w13356;
w13358 <= not w13355 and w13357;
w13359 <= not w13315 and not w13358;
w13360 <= w13276 and not w13278;
w13361 <= not w13279 and not w13360;
w13362 <= not w13359 and w13361;
w13363 <= not w13279 and not w13362;
w13364 <= w13253 and not w13363;
w13365 <= not w13251 and not w13364;
w13366 <= w13125 and not w13365;
w13367 <= not w13123 and not w13366;
w13368 <= not w13044 and not w13367;
w13369 <= not w13041 and not w13368;
w13370 <= w12994 and not w13017;
w13371 <= not w13369 and not w13370;
w13372 <= not w13018 and w13371;
w13373 <= not w12994 and w13372;
w13374 <= not w5342 and not w5431;
w13375 <= not w4870 and w13374;
w13376 <= not w4873 and w13375;
w13377 <= not w13373 and not w13376;
w13378 <= a(20) and not w13377;
w13379 <= not a(20) and w13377;
w13380 <= not w13378 and not w13379;
w13381 <= w271 and w4937;
w13382 <= w2530 and w13381;
w13383 <= w3370 and w13382;
w13384 <= w1829 and w13383;
w13385 <= w1180 and w13384;
w13386 <= w176 and w13385;
w13387 <= w229 and w13386;
w13388 <= w1187 and w13387;
w13389 <= not w164 and w13388;
w13390 <= not w167 and w13389;
w13391 <= not w219 and w13390;
w13392 <= not w647 and w13391;
w13393 <= not w497 and w13392;
w13394 <= w629 and w3127;
w13395 <= w2741 and w13394;
w13396 <= w923 and w13395;
w13397 <= w740 and w13396;
w13398 <= w13393 and w13397;
w13399 <= w1643 and w13398;
w13400 <= w556 and w13399;
w13401 <= w385 and w13400;
w13402 <= w804 and w13401;
w13403 <= not w492 and w13402;
w13404 <= not w190 and w13403;
w13405 <= not w187 and w13404;
w13406 <= not w818 and w13405;
w13407 <= not w504 and w13406;
w13408 <= not w706 and w13407;
w13409 <= not w810 and w13408;
w13410 <= w12893 and w13409;
w13411 <= not w12893 and not w13409;
w13412 <= not w13410 and not w13411;
w13413 <= w13380 and w13412;
w13414 <= not w13380 and not w13412;
w13415 <= not w13413 and not w13414;
w13416 <= not w12944 and w13415;
w13417 <= w12944 and not w13415;
w13418 <= not w13416 and not w13417;
w13419 <= not w12837 and w13418;
w13420 <= not w13416 and not w13419;
w13421 <= not w13411 and not w13413;
w13422 <= w12966 and not w13421;
w13423 <= not w12966 and w13421;
w13424 <= not w13422 and not w13423;
w13425 <= w13350 and w13351;
w13426 <= not w13352 and not w13425;
w13427 <= w2955 and w13426;
w13428 <= w2963 and w12824;
w13429 <= w2958 and w12704;
w13430 <= not w12826 and not w12828;
w13431 <= w12824 and w13426;
w13432 <= not w12824 and not w13426;
w13433 <= not w13430 and not w13432;
w13434 <= not w13431 and w13433;
w13435 <= not w13430 and not w13434;
w13436 <= not w13431 and not w13434;
w13437 <= not w13432 and w13436;
w13438 <= not w13435 and not w13437;
w13439 <= w10 and not w13438;
w13440 <= not w13429 and not w13439;
w13441 <= not w13428 and w13440;
w13442 <= not w13427 and w13441;
w13443 <= w13424 and not w13442;
w13444 <= not w13424 and w13442;
w13445 <= not w13443 and not w13444;
w13446 <= not w13420 and w13445;
w13447 <= w13420 and not w13445;
w13448 <= not w13446 and not w13447;
w13449 <= w13359 and not w13361;
w13450 <= not w13362 and not w13449;
w13451 <= w3392 and w13450;
w13452 <= not w13342 and w13353;
w13453 <= not w13354 and not w13452;
w13454 <= w3477 and w13453;
w13455 <= w13355 and not w13357;
w13456 <= not w13358 and not w13455;
w13457 <= w3541 and w13456;
w13458 <= not w13454 and not w13457;
w13459 <= not w13451 and w13458;
w13460 <= not w3303 and w13459;
w13461 <= w13453 and w13456;
w13462 <= w13426 and w13453;
w13463 <= not w13426 and not w13453;
w13464 <= not w13462 and not w13463;
w13465 <= not w13436 and w13464;
w13466 <= not w13462 and not w13465;
w13467 <= not w13453 and not w13456;
w13468 <= not w13466 and not w13467;
w13469 <= not w13461 and w13468;
w13470 <= not w13461 and not w13469;
w13471 <= not w13450 and not w13456;
w13472 <= w13450 and w13456;
w13473 <= not w13471 and not w13472;
w13474 <= not w13470 and w13473;
w13475 <= w13470 and not w13473;
w13476 <= not w13474 and not w13475;
w13477 <= w13459 and not w13476;
w13478 <= not w13460 and not w13477;
w13479 <= a(29) and not w13478;
w13480 <= not a(29) and w13478;
w13481 <= not w13479 and not w13480;
w13482 <= w13448 and not w13481;
w13483 <= not w13446 and not w13482;
w13484 <= not w13422 and not w13443;
w13485 <= w3727 and w4723;
w13486 <= w924 and w13485;
w13487 <= w2306 and w13486;
w13488 <= w3479 and w13487;
w13489 <= w220 and w13488;
w13490 <= not w333 and w13489;
w13491 <= not w997 and w13490;
w13492 <= not w554 and w13491;
w13493 <= not w405 and w13492;
w13494 <= not w206 and w13493;
w13495 <= not w60 and w13494;
w13496 <= w3484 and w5669;
w13497 <= w12325 and w13496;
w13498 <= w3324 and w13497;
w13499 <= w12874 and w13498;
w13500 <= w13495 and w13499;
w13501 <= w4228 and w13500;
w13502 <= w1956 and w13501;
w13503 <= w831 and w13502;
w13504 <= w3821 and w13503;
w13505 <= not w782 and w13504;
w13506 <= not w110 and w13505;
w13507 <= not w221 and w13506;
w13508 <= not w498 and w13507;
w13509 <= not w303 and w13508;
w13510 <= not w12966 and w13509;
w13511 <= w12966 and not w13509;
w13512 <= not w13484 and not w13511;
w13513 <= not w13510 and w13512;
w13514 <= not w13484 and not w13513;
w13515 <= not w13510 and not w13513;
w13516 <= not w13511 and w13515;
w13517 <= not w13514 and not w13516;
w13518 <= w13436 and not w13464;
w13519 <= not w13465 and not w13518;
w13520 <= w10 and w13519;
w13521 <= w2955 and w13453;
w13522 <= w2958 and w12824;
w13523 <= w2963 and w13426;
w13524 <= not w13522 and not w13523;
w13525 <= not w13521 and w13524;
w13526 <= not w13520 and w13525;
w13527 <= not w13517 and not w13526;
w13528 <= not w13517 and not w13527;
w13529 <= not w13526 and not w13527;
w13530 <= not w13528 and not w13529;
w13531 <= not w13253 and w13363;
w13532 <= not w13364 and not w13531;
w13533 <= w3392 and w13532;
w13534 <= w3477 and w13456;
w13535 <= w3541 and w13450;
w13536 <= not w13534 and not w13535;
w13537 <= not w13533 and w13536;
w13538 <= not w3303 and w13537;
w13539 <= not w13472 and not w13474;
w13540 <= w13450 and w13532;
w13541 <= not w13450 and not w13532;
w13542 <= not w13539 and not w13541;
w13543 <= not w13540 and w13542;
w13544 <= not w13539 and not w13543;
w13545 <= not w13540 and not w13543;
w13546 <= not w13541 and w13545;
w13547 <= not w13544 and not w13546;
w13548 <= w13537 and w13547;
w13549 <= not w13538 and not w13548;
w13550 <= a(29) and not w13549;
w13551 <= not a(29) and w13549;
w13552 <= not w13550 and not w13551;
w13553 <= not w13530 and not w13552;
w13554 <= w13530 and w13552;
w13555 <= not w13553 and not w13554;
w13556 <= not w13483 and w13555;
w13557 <= w13483 and not w13555;
w13558 <= not w13556 and not w13557;
w13559 <= not w13369 and not w13372;
w13560 <= not w13370 and not w13372;
w13561 <= not w13018 and w13560;
w13562 <= not w13559 and not w13561;
w13563 <= w3819 and not w13562;
w13564 <= not w13125 and w13365;
w13565 <= not w13366 and not w13564;
w13566 <= w3902 and w13565;
w13567 <= w13044 and w13367;
w13568 <= not w13368 and not w13567;
w13569 <= w3981 and w13568;
w13570 <= not w13566 and not w13569;
w13571 <= not w13563 and w13570;
w13572 <= w13565 and w13568;
w13573 <= w13532 and w13565;
w13574 <= not w13532 and not w13565;
w13575 <= not w13573 and not w13574;
w13576 <= not w13545 and w13575;
w13577 <= not w13573 and not w13576;
w13578 <= not w13565 and not w13568;
w13579 <= not w13572 and not w13578;
w13580 <= not w13577 and w13579;
w13581 <= not w13572 and not w13580;
w13582 <= not w13562 and w13568;
w13583 <= w13562 and not w13568;
w13584 <= not w13581 and not w13583;
w13585 <= not w13582 and w13584;
w13586 <= not w13581 and not w13585;
w13587 <= not w13582 and not w13585;
w13588 <= not w13583 and w13587;
w13589 <= not w13586 and not w13588;
w13590 <= w3985 and not w13589;
w13591 <= w13571 and not w13590;
w13592 <= a(26) and not w13591;
w13593 <= a(26) and not w13592;
w13594 <= not w13591 and not w13592;
w13595 <= not w13593 and not w13594;
w13596 <= w13558 and not w13595;
w13597 <= w13558 and not w13596;
w13598 <= not w13595 and not w13596;
w13599 <= not w13597 and not w13598;
w13600 <= w13418 and not w13419;
w13601 <= not w12837 and not w13419;
w13602 <= not w13600 and not w13601;
w13603 <= not w12941 and not w12943;
w13604 <= not w12932 and w12944;
w13605 <= not w13603 and not w13604;
w13606 <= not w265 and not w287;
w13607 <= not w1007 and w2744;
w13608 <= not w782 and w13607;
w13609 <= not w492 and w13608;
w13610 <= not w352 and w13609;
w13611 <= not w503 and w13610;
w13612 <= not w140 and w13611;
w13613 <= w1372 and w2155;
w13614 <= w2422 and w13613;
w13615 <= w2280 and w13614;
w13616 <= w13612 and w13615;
w13617 <= w707 and w13616;
w13618 <= w3043 and w13617;
w13619 <= w5199 and w13618;
w13620 <= w4721 and w13619;
w13621 <= w1759 and w13620;
w13622 <= w2518 and w13621;
w13623 <= w2401 and w13622;
w13624 <= not w124 and w13623;
w13625 <= w13606 and w13624;
w13626 <= not w591 and w13625;
w13627 <= not w427 and w13626;
w13628 <= not w136 and w13627;
w13629 <= not w405 and w13628;
w13630 <= not w21 and w13629;
w13631 <= not w591 and not w744;
w13632 <= not w80 and w13631;
w13633 <= not w424 and w13632;
w13634 <= w356 and not w574;
w13635 <= not w527 and w13634;
w13636 <= w2688 and w13635;
w13637 <= w6607 and w13636;
w13638 <= w13073 and w13637;
w13639 <= w13633 and w13638;
w13640 <= w12854 and w13639;
w13641 <= w4750 and w13640;
w13642 <= w2540 and w13641;
w13643 <= w1510 and w13642;
w13644 <= w2341 and w13643;
w13645 <= w137 and w13644;
w13646 <= w1315 and w13645;
w13647 <= not w71 and w13646;
w13648 <= not w262 and w13647;
w13649 <= not w328 and w13648;
w13650 <= not w205 and w13649;
w13651 <= not w13630 and not w13650;
w13652 <= not w5874 and not w6168;
w13653 <= not w5598 and w13652;
w13654 <= not w5601 and w13653;
w13655 <= not w13373 and not w13654;
w13656 <= a(17) and not w13655;
w13657 <= not a(17) and w13655;
w13658 <= not w13656 and not w13657;
w13659 <= w13630 and w13650;
w13660 <= not w13651 and not w13659;
w13661 <= w13658 and w13660;
w13662 <= not w13651 and not w13661;
w13663 <= w12893 and not w13662;
w13664 <= not w12893 and w13662;
w13665 <= not w13663 and not w13664;
w13666 <= w2955 and w12437;
w13667 <= w2963 and w12305;
w13668 <= w2958 and w12440;
w13669 <= not w12615 and not w12618;
w13670 <= not w12616 and w12619;
w13671 <= not w13669 and not w13670;
w13672 <= w10 and not w13671;
w13673 <= not w13668 and not w13672;
w13674 <= not w13667 and w13673;
w13675 <= not w13666 and w13674;
w13676 <= w13665 and not w13675;
w13677 <= not w13663 and not w13676;
w13678 <= not w13605 and not w13677;
w13679 <= w13605 and w13677;
w13680 <= not w13678 and not w13679;
w13681 <= not w12611 and not w12614;
w13682 <= not w12612 and w12615;
w13683 <= not w13681 and not w13682;
w13684 <= w10 and not w13683;
w13685 <= w2955 and w12305;
w13686 <= w2958 and w12443;
w13687 <= w2963 and w12440;
w13688 <= not w13686 and not w13687;
w13689 <= not w13685 and w13688;
w13690 <= not w13684 and w13689;
w13691 <= not w13658 and not w13660;
w13692 <= not w13661 and not w13691;
w13693 <= not w13690 and w13692;
w13694 <= w1188 and w2674;
w13695 <= w2025 and w13694;
w13696 <= w173 and w13695;
w13697 <= not w362 and w13696;
w13698 <= not w270 and w13697;
w13699 <= not w215 and w13698;
w13700 <= not w174 and w13699;
w13701 <= not w395 and w13700;
w13702 <= not w592 and w13701;
w13703 <= not w21 and w13702;
w13704 <= not w552 and not w1241;
w13705 <= not w687 and w13704;
w13706 <= not w537 and w13705;
w13707 <= not w221 and w13706;
w13708 <= not w467 and w13707;
w13709 <= not w65 and not w79;
w13710 <= w3095 and w13709;
w13711 <= w13708 and w13710;
w13712 <= w4260 and w13711;
w13713 <= w5955 and w13712;
w13714 <= w1301 and w13713;
w13715 <= not w602 and w13714;
w13716 <= not w167 and w13715;
w13717 <= not w430 and w13716;
w13718 <= not w370 and w13717;
w13719 <= not w183 and w13718;
w13720 <= not w26 and w13719;
w13721 <= not w207 and w13720;
w13722 <= not w821 and w13721;
w13723 <= w2618 and w13722;
w13724 <= not w103 and w13723;
w13725 <= w1243 and w13724;
w13726 <= w1877 and w13725;
w13727 <= w5726 and w13726;
w13728 <= w2731 and w13727;
w13729 <= w13703 and w13728;
w13730 <= w1510 and w13729;
w13731 <= w2419 and w13730;
w13732 <= w94 and w13731;
w13733 <= w1096 and w13732;
w13734 <= not w164 and w13733;
w13735 <= not w264 and w13734;
w13736 <= not w288 and w13735;
w13737 <= not w574 and w13736;
w13738 <= not w502 and w13737;
w13739 <= not w647 and w13738;
w13740 <= not w239 and w13739;
w13741 <= w13630 and not w13740;
w13742 <= not w71 and w5017;
w13743 <= not w819 and w13742;
w13744 <= w5206 and w13743;
w13745 <= w2976 and w13744;
w13746 <= w2651 and w13745;
w13747 <= w3424 and w13746;
w13748 <= w4302 and w13747;
w13749 <= w1015 and w13748;
w13750 <= not w453 and w13749;
w13751 <= not w537 and w13750;
w13752 <= not w81 and w13751;
w13753 <= w823 and w13752;
w13754 <= not w608 and w13753;
w13755 <= not w499 and w13754;
w13756 <= not w60 and w13755;
w13757 <= w358 and w1301;
w13758 <= not w86 and w13757;
w13759 <= not w472 and w13758;
w13760 <= not w310 and w13759;
w13761 <= not w157 and w13760;
w13762 <= w708 and w1463;
w13763 <= w1281 and w13762;
w13764 <= w4233 and w13763;
w13765 <= w3003 and w13764;
w13766 <= w369 and w13765;
w13767 <= w13761 and w13766;
w13768 <= w1749 and w13767;
w13769 <= w6449 and w13768;
w13770 <= w709 and w13769;
w13771 <= w1773 and w13770;
w13772 <= not w167 and w13771;
w13773 <= not w572 and w13772;
w13774 <= not w163 and w13773;
w13775 <= not w237 and w13774;
w13776 <= not w233 and w13775;
w13777 <= not w230 and w13776;
w13778 <= not w62 and w13777;
w13779 <= not w13756 and not w13778;
w13780 <= not w6886 and not w7036;
w13781 <= not w6337 and w13780;
w13782 <= not w6332 and w13781;
w13783 <= not w13373 and not w13782;
w13784 <= a(14) and not w13783;
w13785 <= not a(14) and w13783;
w13786 <= not w13784 and not w13785;
w13787 <= w13756 and w13778;
w13788 <= not w13779 and not w13787;
w13789 <= w13786 and w13788;
w13790 <= not w13779 and not w13789;
w13791 <= w13740 and not w13790;
w13792 <= not w13740 and w13790;
w13793 <= not w13791 and not w13792;
w13794 <= w2955 and w12443;
w13795 <= w2963 and w12448;
w13796 <= w2958 and w12446;
w13797 <= w12602 and not w12605;
w13798 <= not w12606 and not w13797;
w13799 <= w10 and w13798;
w13800 <= not w13796 and not w13799;
w13801 <= not w13795 and w13800;
w13802 <= not w13794 and w13801;
w13803 <= w13793 and not w13802;
w13804 <= not w13791 and not w13803;
w13805 <= not w13630 and w13740;
w13806 <= not w13804 and not w13805;
w13807 <= not w13741 and w13806;
w13808 <= not w13741 and not w13807;
w13809 <= w13692 and not w13693;
w13810 <= not w13690 and not w13693;
w13811 <= not w13809 and not w13810;
w13812 <= not w13808 and not w13811;
w13813 <= not w13693 and not w13812;
w13814 <= not w13665 and w13675;
w13815 <= not w13676 and not w13814;
w13816 <= not w13813 and w13815;
w13817 <= w13813 and not w13815;
w13818 <= not w13816 and not w13817;
w13819 <= w3392 and w13426;
w13820 <= w3477 and w12704;
w13821 <= w3541 and w12824;
w13822 <= not w13820 and not w13821;
w13823 <= not w13819 and w13822;
w13824 <= not w3303 and w13823;
w13825 <= w13438 and w13823;
w13826 <= not w13824 and not w13825;
w13827 <= a(29) and not w13826;
w13828 <= not a(29) and w13826;
w13829 <= not w13827 and not w13828;
w13830 <= w13818 and not w13829;
w13831 <= not w13816 and not w13830;
w13832 <= w13680 and not w13831;
w13833 <= not w13678 and not w13832;
w13834 <= not w13602 and not w13833;
w13835 <= w13602 and w13833;
w13836 <= not w13834 and not w13835;
w13837 <= w3392 and w13456;
w13838 <= w3477 and w13426;
w13839 <= w3541 and w13453;
w13840 <= not w13838 and not w13839;
w13841 <= not w13837 and w13840;
w13842 <= not w13466 and not w13469;
w13843 <= not w13467 and w13470;
w13844 <= not w13842 and not w13843;
w13845 <= w3303 and not w13844;
w13846 <= w13841 and not w13845;
w13847 <= a(29) and not w13846;
w13848 <= a(29) and not w13847;
w13849 <= not w13846 and not w13847;
w13850 <= not w13848 and not w13849;
w13851 <= w13836 and not w13850;
w13852 <= not w13834 and not w13851;
w13853 <= not w13448 and w13481;
w13854 <= not w13482 and not w13853;
w13855 <= not w13852 and w13854;
w13856 <= w13852 and not w13854;
w13857 <= not w13855 and not w13856;
w13858 <= w3819 and w13568;
w13859 <= w3902 and w13532;
w13860 <= w3981 and w13565;
w13861 <= not w13859 and not w13860;
w13862 <= not w13858 and w13861;
w13863 <= w13577 and not w13579;
w13864 <= not w13580 and not w13863;
w13865 <= w3985 and w13864;
w13866 <= w13862 and not w13865;
w13867 <= a(26) and not w13866;
w13868 <= a(26) and not w13867;
w13869 <= not w13866 and not w13867;
w13870 <= not w13868 and not w13869;
w13871 <= w13857 and not w13870;
w13872 <= not w13855 and not w13871;
w13873 <= not w4539 and not w4629;
w13874 <= not w13373 and not w13873;
w13875 <= w12994 and w13560;
w13876 <= not w13373 and not w13875;
w13877 <= w4468 and w13876;
w13878 <= not w13874 and not w13877;
w13879 <= not w4471 and w13878;
w13880 <= not w13562 and w13876;
w13881 <= w13562 and not w13876;
w13882 <= not w13880 and not w13881;
w13883 <= not w13587 and w13882;
w13884 <= not w13880 and not w13883;
w13885 <= w13875 and not w13884;
w13886 <= not w13876 and not w13885;
w13887 <= w13878 and w13886;
w13888 <= not w13879 and not w13887;
w13889 <= a(23) and not w13888;
w13890 <= not a(23) and w13888;
w13891 <= not w13889 and not w13890;
w13892 <= not w13872 and not w13891;
w13893 <= w13872 and w13891;
w13894 <= not w13892 and not w13893;
w13895 <= not w13599 and w13894;
w13896 <= not w13599 and not w13895;
w13897 <= w13894 and not w13895;
w13898 <= not w13896 and not w13897;
w13899 <= w13857 and not w13871;
w13900 <= not w13870 and not w13871;
w13901 <= not w13899 and not w13900;
w13902 <= w13836 and not w13851;
w13903 <= not w13850 and not w13851;
w13904 <= not w13902 and not w13903;
w13905 <= w3819 and w13565;
w13906 <= w3902 and w13450;
w13907 <= w3981 and w13532;
w13908 <= not w13906 and not w13907;
w13909 <= not w13905 and w13908;
w13910 <= w13545 and not w13575;
w13911 <= not w13576 and not w13910;
w13912 <= w3985 and w13911;
w13913 <= w13909 and not w13912;
w13914 <= a(26) and not w13913;
w13915 <= a(26) and not w13914;
w13916 <= not w13913 and not w13914;
w13917 <= not w13915 and not w13916;
w13918 <= not w13904 and not w13917;
w13919 <= not w13904 and not w13918;
w13920 <= not w13917 and not w13918;
w13921 <= not w13919 and not w13920;
w13922 <= not w13680 and w13831;
w13923 <= not w13832 and not w13922;
w13924 <= w3392 and w13453;
w13925 <= w3477 and w12824;
w13926 <= w3541 and w13426;
w13927 <= not w13925 and not w13926;
w13928 <= not w13924 and w13927;
w13929 <= w3303 and w13519;
w13930 <= w13928 and not w13929;
w13931 <= a(29) and not w13930;
w13932 <= a(29) and not w13931;
w13933 <= not w13930 and not w13931;
w13934 <= not w13932 and not w13933;
w13935 <= w13923 and not w13934;
w13936 <= w13923 and not w13935;
w13937 <= not w13934 and not w13935;
w13938 <= not w13936 and not w13937;
w13939 <= w3819 and w13532;
w13940 <= w3902 and w13456;
w13941 <= w3981 and w13450;
w13942 <= not w13940 and not w13941;
w13943 <= not w13939 and w13942;
w13944 <= w3985 and not w13547;
w13945 <= w13943 and not w13944;
w13946 <= a(26) and not w13945;
w13947 <= a(26) and not w13946;
w13948 <= not w13945 and not w13946;
w13949 <= not w13947 and not w13948;
w13950 <= not w13938 and not w13949;
w13951 <= not w13935 and not w13950;
w13952 <= not w13921 and not w13951;
w13953 <= not w13918 and not w13952;
w13954 <= not w13901 and not w13953;
w13955 <= w13901 and w13953;
w13956 <= not w13954 and not w13955;
w13957 <= w4629 and not w13373;
w13958 <= w4468 and not w13562;
w13959 <= w4539 and w13876;
w13960 <= not w13958 and not w13959;
w13961 <= not w13957 and w13960;
w13962 <= not w13875 and w13884;
w13963 <= not w13885 and not w13962;
w13964 <= w4471 and w13963;
w13965 <= w13961 and not w13964;
w13966 <= a(23) and not w13965;
w13967 <= a(23) and not w13966;
w13968 <= not w13965 and not w13966;
w13969 <= not w13967 and not w13968;
w13970 <= w13956 and not w13969;
w13971 <= not w13954 and not w13970;
w13972 <= not w13898 and not w13971;
w13973 <= w13898 and w13971;
w13974 <= not w13972 and not w13973;
w13975 <= w13956 and not w13970;
w13976 <= not w13969 and not w13970;
w13977 <= not w13975 and not w13976;
w13978 <= not w13938 and not w13950;
w13979 <= not w13949 and not w13950;
w13980 <= not w13978 and not w13979;
w13981 <= not w13804 and not w13807;
w13982 <= not w13805 and w13808;
w13983 <= not w13981 and not w13982;
w13984 <= not w12607 and not w12610;
w13985 <= not w12608 and w12611;
w13986 <= not w13984 and not w13985;
w13987 <= w10 and not w13986;
w13988 <= w2955 and w12440;
w13989 <= w2958 and w12448;
w13990 <= w2963 and w12443;
w13991 <= not w13989 and not w13990;
w13992 <= not w13988 and w13991;
w13993 <= not w13987 and w13992;
w13994 <= not w13983 and not w13993;
w13995 <= not w13983 and not w13994;
w13996 <= not w13993 and not w13994;
w13997 <= not w13995 and not w13996;
w13998 <= w3392 and w12704;
w13999 <= w3477 and w12305;
w14000 <= w3541 and w12437;
w14001 <= not w13999 and not w14000;
w14002 <= not w13998 and w14001;
w14003 <= not w3303 and w14002;
w14004 <= not w12934 and w14002;
w14005 <= not w14003 and not w14004;
w14006 <= a(29) and not w14005;
w14007 <= not a(29) and w14005;
w14008 <= not w14006 and not w14007;
w14009 <= not w13997 and not w14008;
w14010 <= not w13994 and not w14009;
w14011 <= not w13811 and not w13812;
w14012 <= not w13808 and not w13812;
w14013 <= not w14011 and not w14012;
w14014 <= not w14010 and not w14013;
w14015 <= not w14010 and not w14014;
w14016 <= not w14013 and not w14014;
w14017 <= not w14015 and not w14016;
w14018 <= w3392 and w12824;
w14019 <= w3477 and w12437;
w14020 <= w3541 and w12704;
w14021 <= not w14019 and not w14020;
w14022 <= not w14018 and w14021;
w14023 <= w3303 and w12830;
w14024 <= w14022 and not w14023;
w14025 <= a(29) and not w14024;
w14026 <= a(29) and not w14025;
w14027 <= not w14024 and not w14025;
w14028 <= not w14026 and not w14027;
w14029 <= not w14017 and not w14028;
w14030 <= not w14014 and not w14029;
w14031 <= not w13818 and w13829;
w14032 <= not w13830 and not w14031;
w14033 <= not w14030 and w14032;
w14034 <= w14030 and not w14032;
w14035 <= not w14033 and not w14034;
w14036 <= w3819 and w13450;
w14037 <= w3902 and w13453;
w14038 <= w3981 and w13456;
w14039 <= not w14037 and not w14038;
w14040 <= not w14036 and w14039;
w14041 <= w3985 and w13476;
w14042 <= w14040 and not w14041;
w14043 <= a(26) and not w14042;
w14044 <= a(26) and not w14043;
w14045 <= not w14042 and not w14043;
w14046 <= not w14044 and not w14045;
w14047 <= w14035 and not w14046;
w14048 <= not w14033 and not w14047;
w14049 <= not w13980 and not w14048;
w14050 <= w13980 and w14048;
w14051 <= not w14049 and not w14050;
w14052 <= w4629 and not w13562;
w14053 <= w4468 and w13565;
w14054 <= w4539 and w13568;
w14055 <= not w14053 and not w14054;
w14056 <= not w14052 and w14055;
w14057 <= w4471 and not w13589;
w14058 <= w14056 and not w14057;
w14059 <= a(23) and not w14058;
w14060 <= a(23) and not w14059;
w14061 <= not w14058 and not w14059;
w14062 <= not w14060 and not w14061;
w14063 <= w14051 and not w14062;
w14064 <= not w14049 and not w14063;
w14065 <= w4629 and w13876;
w14066 <= w4468 and w13568;
w14067 <= w4539 and not w13562;
w14068 <= not w14066 and not w14067;
w14069 <= not w14065 and w14068;
w14070 <= w13587 and not w13882;
w14071 <= not w13883 and not w14070;
w14072 <= w4471 and w14071;
w14073 <= w14069 and not w14072;
w14074 <= a(23) and not w14073;
w14075 <= a(23) and not w14074;
w14076 <= not w14073 and not w14074;
w14077 <= not w14075 and not w14076;
w14078 <= not w14064 and not w14077;
w14079 <= w13921 and w13951;
w14080 <= not w13952 and not w14079;
w14081 <= not w14064 and not w14078;
w14082 <= not w14077 and not w14078;
w14083 <= not w14081 and not w14082;
w14084 <= w14080 and not w14083;
w14085 <= not w14078 and not w14084;
w14086 <= not w13977 and not w14085;
w14087 <= not w13977 and not w14086;
w14088 <= not w14085 and not w14086;
w14089 <= not w14087 and not w14088;
w14090 <= w14035 and not w14047;
w14091 <= not w14046 and not w14047;
w14092 <= not w14090 and not w14091;
w14093 <= not w14017 and not w14029;
w14094 <= not w14028 and not w14029;
w14095 <= not w14093 and not w14094;
w14096 <= w3819 and w13456;
w14097 <= w3902 and w13426;
w14098 <= w3981 and w13453;
w14099 <= not w14097 and not w14098;
w14100 <= not w14096 and w14099;
w14101 <= w3985 and not w13844;
w14102 <= w14100 and not w14101;
w14103 <= a(26) and not w14102;
w14104 <= a(26) and not w14103;
w14105 <= not w14102 and not w14103;
w14106 <= not w14104 and not w14105;
w14107 <= not w14095 and not w14106;
w14108 <= not w14095 and not w14107;
w14109 <= not w14106 and not w14107;
w14110 <= not w14108 and not w14109;
w14111 <= w12598 and not w12600;
w14112 <= not w12601 and not w14111;
w14113 <= w10 and w14112;
w14114 <= w2955 and w12448;
w14115 <= w2958 and w12451;
w14116 <= w2963 and w12446;
w14117 <= not w14115 and not w14116;
w14118 <= not w14114 and w14117;
w14119 <= not w14113 and w14118;
w14120 <= not w77 and not w441;
w14121 <= not w357 and w14120;
w14122 <= not w538 and w14121;
w14123 <= not w65 and w14122;
w14124 <= not w267 and w14123;
w14125 <= w1044 and w3458;
w14126 <= w5712 and w14125;
w14127 <= w14124 and w14126;
w14128 <= w1957 and w14127;
w14129 <= w557 and w14128;
w14130 <= w809 and w14129;
w14131 <= w709 and w14130;
w14132 <= w807 and w14131;
w14133 <= w291 and w14132;
w14134 <= not w1241 and w14133;
w14135 <= not w338 and w14134;
w14136 <= not w96 and w14135;
w14137 <= not w590 and w14136;
w14138 <= w577 and w3100;
w14139 <= w2325 and w14138;
w14140 <= w924 and w14139;
w14141 <= w1717 and w14140;
w14142 <= not w946 and w14141;
w14143 <= not w782 and w14142;
w14144 <= not w266 and w14143;
w14145 <= not w67 and w14144;
w14146 <= w464 and w14145;
w14147 <= w3616 and w14146;
w14148 <= w2231 and w14147;
w14149 <= w14137 and w14148;
w14150 <= w981 and w14149;
w14151 <= w385 and w14150;
w14152 <= w872 and w14151;
w14153 <= w2023 and w14152;
w14154 <= w4036 and w14153;
w14155 <= w1457 and w14154;
w14156 <= not w71 and w14155;
w14157 <= not w997 and w14156;
w14158 <= not w237 and w14157;
w14159 <= not w127 and w14158;
w14160 <= not w365 and w14159;
w14161 <= not w136 and w14160;
w14162 <= not w592 and w14161;
w14163 <= not w93 and w14162;
w14164 <= w13756 and not w14163;
w14165 <= not w13756 and w14163;
w14166 <= not w12594 and not w12597;
w14167 <= not w12595 and w12598;
w14168 <= not w14166 and not w14167;
w14169 <= w10 and not w14168;
w14170 <= w2955 and w12446;
w14171 <= w2958 and w12454;
w14172 <= w2963 and w12451;
w14173 <= not w14171 and not w14172;
w14174 <= not w14170 and w14173;
w14175 <= not w14169 and w14174;
w14176 <= not w14164 and not w14175;
w14177 <= not w14165 and w14176;
w14178 <= not w14164 and not w14177;
w14179 <= not w13786 and not w13788;
w14180 <= not w13789 and not w14179;
w14181 <= not w14178 and w14180;
w14182 <= w14178 and not w14180;
w14183 <= not w14181 and not w14182;
w14184 <= not w14119 and w14183;
w14185 <= not w14181 and not w14184;
w14186 <= not w13793 and w13802;
w14187 <= not w13803 and not w14186;
w14188 <= not w14185 and w14187;
w14189 <= w14185 and not w14187;
w14190 <= not w14188 and not w14189;
w14191 <= w3392 and w12437;
w14192 <= w3477 and w12440;
w14193 <= w3541 and w12305;
w14194 <= not w14192 and not w14193;
w14195 <= not w14191 and w14194;
w14196 <= not w3303 and w14195;
w14197 <= w13671 and w14195;
w14198 <= not w14196 and not w14197;
w14199 <= a(29) and not w14198;
w14200 <= not a(29) and w14198;
w14201 <= not w14199 and not w14200;
w14202 <= w14190 and not w14201;
w14203 <= not w14188 and not w14202;
w14204 <= w13997 and w14008;
w14205 <= not w14009 and not w14204;
w14206 <= not w14203 and w14205;
w14207 <= w14203 and not w14205;
w14208 <= not w14206 and not w14207;
w14209 <= w3819 and w13453;
w14210 <= w3902 and w12824;
w14211 <= w3981 and w13426;
w14212 <= not w14210 and not w14211;
w14213 <= not w14209 and w14212;
w14214 <= w3985 and w13519;
w14215 <= w14213 and not w14214;
w14216 <= a(26) and not w14215;
w14217 <= a(26) and not w14216;
w14218 <= not w14215 and not w14216;
w14219 <= not w14217 and not w14218;
w14220 <= w14208 and not w14219;
w14221 <= not w14206 and not w14220;
w14222 <= not w14110 and not w14221;
w14223 <= not w14107 and not w14222;
w14224 <= not w14092 and not w14223;
w14225 <= w14092 and w14223;
w14226 <= not w14224 and not w14225;
w14227 <= w4629 and w13568;
w14228 <= w4468 and w13532;
w14229 <= w4539 and w13565;
w14230 <= not w14228 and not w14229;
w14231 <= not w14227 and w14230;
w14232 <= w4471 and w13864;
w14233 <= w14231 and not w14232;
w14234 <= a(23) and not w14233;
w14235 <= a(23) and not w14234;
w14236 <= not w14233 and not w14234;
w14237 <= not w14235 and not w14236;
w14238 <= w14226 and not w14237;
w14239 <= not w14224 and not w14238;
w14240 <= not w13373 and not w13374;
w14241 <= w4870 and w13876;
w14242 <= not w14240 and not w14241;
w14243 <= not w4873 and w14242;
w14244 <= w13886 and w14242;
w14245 <= not w14243 and not w14244;
w14246 <= a(20) and not w14245;
w14247 <= not a(20) and w14245;
w14248 <= not w14246 and not w14247;
w14249 <= not w14239 and not w14248;
w14250 <= w14051 and not w14063;
w14251 <= not w14062 and not w14063;
w14252 <= not w14250 and not w14251;
w14253 <= w14239 and w14248;
w14254 <= not w14249 and not w14253;
w14255 <= not w14252 and w14254;
w14256 <= not w14249 and not w14255;
w14257 <= not w14080 and w14083;
w14258 <= not w14084 and not w14257;
w14259 <= not w14256 and w14258;
w14260 <= not w14252 and not w14255;
w14261 <= w14254 and not w14255;
w14262 <= not w14260 and not w14261;
w14263 <= w14226 and not w14238;
w14264 <= not w14237 and not w14238;
w14265 <= not w14263 and not w14264;
w14266 <= w14110 and w14221;
w14267 <= not w14222 and not w14266;
w14268 <= w4629 and w13565;
w14269 <= w4468 and w13450;
w14270 <= w4539 and w13532;
w14271 <= not w14269 and not w14270;
w14272 <= not w14268 and w14271;
w14273 <= w4471 and w13911;
w14274 <= w14272 and not w14273;
w14275 <= a(23) and not w14274;
w14276 <= a(23) and not w14275;
w14277 <= not w14274 and not w14275;
w14278 <= not w14276 and not w14277;
w14279 <= w14267 and not w14278;
w14280 <= w14267 and not w14279;
w14281 <= not w14278 and not w14279;
w14282 <= not w14280 and not w14281;
w14283 <= w14208 and not w14220;
w14284 <= not w14219 and not w14220;
w14285 <= not w14283 and not w14284;
w14286 <= w14183 and not w14184;
w14287 <= not w14119 and not w14184;
w14288 <= not w14286 and not w14287;
w14289 <= w3392 and w12305;
w14290 <= w3477 and w12443;
w14291 <= w3541 and w12440;
w14292 <= not w14290 and not w14291;
w14293 <= not w14289 and w14292;
w14294 <= w3303 and not w13683;
w14295 <= w14293 and not w14294;
w14296 <= a(29) and not w14295;
w14297 <= a(29) and not w14296;
w14298 <= not w14295 and not w14296;
w14299 <= not w14297 and not w14298;
w14300 <= not w14288 and not w14299;
w14301 <= not w14288 and not w14300;
w14302 <= not w14299 and not w14300;
w14303 <= not w14301 and not w14302;
w14304 <= not w14175 and not w14177;
w14305 <= not w14165 and w14178;
w14306 <= not w14304 and not w14305;
w14307 <= w1206 and w1537;
w14308 <= w2633 and w14307;
w14309 <= not w58 and w14308;
w14310 <= not w492 and w14309;
w14311 <= not w506 and w14310;
w14312 <= not w448 and w14311;
w14313 <= not w425 and w14312;
w14314 <= not w237 and w14313;
w14315 <= not w126 and w14314;
w14316 <= not w307 and w14315;
w14317 <= not w213 and w4999;
w14318 <= not w183 and w14317;
w14319 <= not w338 and w14318;
w14320 <= not w99 and w14319;
w14321 <= not w301 and w14320;
w14322 <= w1931 and w13049;
w14323 <= w4065 and w14322;
w14324 <= w1957 and w14323;
w14325 <= w14321 and w14324;
w14326 <= w2707 and w14325;
w14327 <= w6032 and w14326;
w14328 <= w14316 and w14327;
w14329 <= w2518 and w14328;
w14330 <= w1302 and w14329;
w14331 <= w1324 and w14330;
w14332 <= not w355 and w14331;
w14333 <= not w216 and w14332;
w14334 <= w4229 and w14333;
w14335 <= not w328 and w14334;
w14336 <= not w207 and w14335;
w14337 <= not w607 and w14336;
w14338 <= not w306 and w14337;
w14339 <= w1075 and w2145;
w14340 <= not w554 and w14339;
w14341 <= not w92 and w14340;
w14342 <= not w60 and w14341;
w14343 <= w824 and w2298;
w14344 <= w2479 and w14343;
w14345 <= w1020 and w14344;
w14346 <= w5681 and w14345;
w14347 <= w1054 and w14346;
w14348 <= w203 and w14347;
w14349 <= w3340 and w14348;
w14350 <= w3407 and w14349;
w14351 <= w14342 and w14350;
w14352 <= w868 and w14351;
w14353 <= w4230 and w14352;
w14354 <= not w103 and w14353;
w14355 <= not w335 and w14354;
w14356 <= not w141 and w14355;
w14357 <= not w80 and w14356;
w14358 <= not w14338 and not w14357;
w14359 <= not w7567 and not w7918;
w14360 <= not w7226 and w14359;
w14361 <= not w7229 and w14360;
w14362 <= not w13373 and not w14361;
w14363 <= a(11) and not w14362;
w14364 <= not a(11) and w14362;
w14365 <= not w14363 and not w14364;
w14366 <= w14338 and w14357;
w14367 <= not w14358 and not w14366;
w14368 <= w14365 and w14367;
w14369 <= not w14358 and not w14368;
w14370 <= w13756 and not w14369;
w14371 <= not w13756 and w14369;
w14372 <= not w14370 and not w14371;
w14373 <= w2955 and w12451;
w14374 <= w2963 and w12454;
w14375 <= w2958 and w12457;
w14376 <= not w12590 and not w12593;
w14377 <= not w12591 and w12594;
w14378 <= not w14376 and not w14377;
w14379 <= w10 and not w14378;
w14380 <= not w14375 and not w14379;
w14381 <= not w14374 and w14380;
w14382 <= not w14373 and w14381;
w14383 <= w14372 and not w14382;
w14384 <= not w14370 and not w14383;
w14385 <= not w14306 and not w14384;
w14386 <= w14306 and w14384;
w14387 <= not w14385 and not w14386;
w14388 <= w12586 and not w12588;
w14389 <= not w12589 and not w14388;
w14390 <= w10 and w14389;
w14391 <= w2955 and w12454;
w14392 <= w2958 and w12460;
w14393 <= w2963 and w12457;
w14394 <= not w14392 and not w14393;
w14395 <= not w14391 and w14394;
w14396 <= not w14390 and w14395;
w14397 <= not w14365 and not w14367;
w14398 <= not w14368 and not w14397;
w14399 <= not w14396 and w14398;
w14400 <= w14398 and not w14399;
w14401 <= not w14396 and not w14399;
w14402 <= not w14400 and not w14401;
w14403 <= w1139 and w2089;
w14404 <= w600 and w14403;
w14405 <= not w552 and w14404;
w14406 <= not w104 and w14405;
w14407 <= not w602 and w14406;
w14408 <= not w337 and w14407;
w14409 <= not w425 and w14408;
w14410 <= not w309 and w14409;
w14411 <= not w67 and w14410;
w14412 <= not w536 and not w1036;
w14413 <= not w186 and w14412;
w14414 <= not w205 and w14413;
w14415 <= w445 and not w744;
w14416 <= not w503 and w14415;
w14417 <= not w359 and w14416;
w14418 <= w1360 and w3484;
w14419 <= w2588 and w14418;
w14420 <= w14417 and w14419;
w14421 <= w133 and w14420;
w14422 <= w1875 and w14421;
w14423 <= w14414 and w14422;
w14424 <= w1227 and w14423;
w14425 <= w1265 and w14424;
w14426 <= w762 and w14425;
w14427 <= w1315 and w14426;
w14428 <= w1204 and w14427;
w14429 <= not w332 and w14428;
w14430 <= not w1181 and w14429;
w14431 <= not w213 and w14430;
w14432 <= not w30 and w14431;
w14433 <= not w60 and w14432;
w14434 <= w609 and w1581;
w14435 <= w3920 and w14434;
w14436 <= w142 and w14435;
w14437 <= w14433 and w14436;
w14438 <= w4182 and w14437;
w14439 <= w14411 and w14438;
w14440 <= w557 and w14439;
w14441 <= w2674 and w14440;
w14442 <= w94 and w14441;
w14443 <= w291 and w14442;
w14444 <= not w164 and w14443;
w14445 <= not w555 and w14444;
w14446 <= not w183 and w14445;
w14447 <= not w351 and w14446;
w14448 <= not w172 and w14447;
w14449 <= not w54 and w14448;
w14450 <= w14338 and not w14449;
w14451 <= not w14338 and w14449;
w14452 <= not w53 and w389;
w14453 <= not w100 and w14452;
w14454 <= w2283 and w14453;
w14455 <= w1511 and w14454;
w14456 <= not w506 and w14455;
w14457 <= not w529 and w14456;
w14458 <= not w67 and w14457;
w14459 <= not w945 and w14458;
w14460 <= not w205 and w14459;
w14461 <= w278 and w13635;
w14462 <= w1005 and w14461;
w14463 <= w3344 and w14462;
w14464 <= not w997 and w14463;
w14465 <= not w744 and w14464;
w14466 <= not w266 and w14465;
w14467 <= not w624 and w14466;
w14468 <= not w608 and w14467;
w14469 <= not w409 and w14468;
w14470 <= w432 and w1250;
w14471 <= w4067 and w14470;
w14472 <= w2127 and w14471;
w14473 <= w385 and w14472;
w14474 <= w162 and w14473;
w14475 <= not w738 and w14474;
w14476 <= not w370 and w14475;
w14477 <= not w396 and w14476;
w14478 <= not w241 and w14477;
w14479 <= not w172 and w14478;
w14480 <= w1961 and w2930;
w14481 <= w3447 and w14480;
w14482 <= w2252 and w14481;
w14483 <= w3048 and w14482;
w14484 <= w14479 and w14483;
w14485 <= w14469 and w14484;
w14486 <= w14460 and w14485;
w14487 <= w2568 and w14486;
w14488 <= w2378 and w14487;
w14489 <= w655 and w14488;
w14490 <= w291 and w14489;
w14491 <= w1115 and w14490;
w14492 <= not w129 and w14491;
w14493 <= not w269 and w14492;
w14494 <= not w60 and w14493;
w14495 <= not w529 and not w651;
w14496 <= not w266 and w14495;
w14497 <= not w1181 and w14496;
w14498 <= not w224 and w14497;
w14499 <= not w462 and w14498;
w14500 <= not w136 and w14499;
w14501 <= w1630 and w1947;
w14502 <= w1537 and w14501;
w14503 <= w745 and w14502;
w14504 <= not w86 and w14503;
w14505 <= not w221 and w14504;
w14506 <= not w431 and w14505;
w14507 <= not w207 and w14506;
w14508 <= w1831 and w2228;
w14509 <= w628 and w14508;
w14510 <= w4971 and w14509;
w14511 <= w1627 and w14510;
w14512 <= w13200 and w14511;
w14513 <= w14507 and w14512;
w14514 <= w1035 and w14513;
w14515 <= w55 and w14514;
w14516 <= w14500 and w14515;
w14517 <= w294 and w14516;
w14518 <= not w362 and w14517;
w14519 <= not w332 and w14518;
w14520 <= not w141 and w14519;
w14521 <= not w440 and w14520;
w14522 <= not w105 and w14521;
w14523 <= not w428 and w14522;
w14524 <= not w14494 and not w14523;
w14525 <= not w8795 and not w9266;
w14526 <= not w8353 and w14525;
w14527 <= not w8356 and w14526;
w14528 <= not w13373 and not w14527;
w14529 <= a(8) and not w14528;
w14530 <= not a(8) and w14528;
w14531 <= not w14529 and not w14530;
w14532 <= w14494 and w14523;
w14533 <= not w14524 and not w14532;
w14534 <= w14531 and w14533;
w14535 <= not w14524 and not w14534;
w14536 <= w14338 and not w14535;
w14537 <= not w14338 and w14535;
w14538 <= not w14536 and not w14537;
w14539 <= w2955 and w12460;
w14540 <= w2963 and w12463;
w14541 <= w2958 and w12466;
w14542 <= w12578 and not w12580;
w14543 <= not w12581 and not w14542;
w14544 <= w10 and w14543;
w14545 <= not w14541 and not w14544;
w14546 <= not w14540 and w14545;
w14547 <= not w14539 and w14546;
w14548 <= w14538 and not w14547;
w14549 <= not w14536 and not w14548;
w14550 <= not w14450 and not w14549;
w14551 <= not w14451 and w14550;
w14552 <= not w14450 and not w14551;
w14553 <= not w14402 and not w14552;
w14554 <= not w14399 and not w14553;
w14555 <= not w14372 and w14382;
w14556 <= not w14383 and not w14555;
w14557 <= not w14554 and w14556;
w14558 <= w14554 and not w14556;
w14559 <= not w14557 and not w14558;
w14560 <= w3392 and w12443;
w14561 <= w3477 and w12446;
w14562 <= w3541 and w12448;
w14563 <= not w14561 and not w14562;
w14564 <= not w14560 and w14563;
w14565 <= not w3303 and w14564;
w14566 <= not w13798 and w14564;
w14567 <= not w14565 and not w14566;
w14568 <= a(29) and not w14567;
w14569 <= not a(29) and w14567;
w14570 <= not w14568 and not w14569;
w14571 <= w14559 and not w14570;
w14572 <= not w14557 and not w14571;
w14573 <= w14387 and not w14572;
w14574 <= not w14385 and not w14573;
w14575 <= not w14303 and not w14574;
w14576 <= not w14300 and not w14575;
w14577 <= not w14190 and w14201;
w14578 <= not w14202 and not w14577;
w14579 <= not w14576 and w14578;
w14580 <= w14576 and not w14578;
w14581 <= not w14579 and not w14580;
w14582 <= w3819 and w13426;
w14583 <= w3902 and w12704;
w14584 <= w3981 and w12824;
w14585 <= not w14583 and not w14584;
w14586 <= not w14582 and w14585;
w14587 <= w3985 and not w13438;
w14588 <= w14586 and not w14587;
w14589 <= a(26) and not w14588;
w14590 <= a(26) and not w14589;
w14591 <= not w14588 and not w14589;
w14592 <= not w14590 and not w14591;
w14593 <= w14581 and not w14592;
w14594 <= not w14579 and not w14593;
w14595 <= not w14285 and not w14594;
w14596 <= w14285 and w14594;
w14597 <= not w14595 and not w14596;
w14598 <= w4629 and w13532;
w14599 <= w4468 and w13456;
w14600 <= w4539 and w13450;
w14601 <= not w14599 and not w14600;
w14602 <= not w14598 and w14601;
w14603 <= w4471 and not w13547;
w14604 <= w14602 and not w14603;
w14605 <= a(23) and not w14604;
w14606 <= a(23) and not w14605;
w14607 <= not w14604 and not w14605;
w14608 <= not w14606 and not w14607;
w14609 <= w14597 and not w14608;
w14610 <= not w14595 and not w14609;
w14611 <= not w14282 and not w14610;
w14612 <= not w14279 and not w14611;
w14613 <= not w14265 and not w14612;
w14614 <= w14265 and w14612;
w14615 <= not w14613 and not w14614;
w14616 <= w5431 and not w13373;
w14617 <= w4870 and not w13562;
w14618 <= w5342 and w13876;
w14619 <= not w14617 and not w14618;
w14620 <= not w14616 and w14619;
w14621 <= w4873 and w13963;
w14622 <= w14620 and not w14621;
w14623 <= a(20) and not w14622;
w14624 <= a(20) and not w14623;
w14625 <= not w14622 and not w14623;
w14626 <= not w14624 and not w14625;
w14627 <= w14615 and not w14626;
w14628 <= not w14613 and not w14627;
w14629 <= not w14262 and not w14628;
w14630 <= w14262 and w14628;
w14631 <= not w14629 and not w14630;
w14632 <= w14615 and not w14627;
w14633 <= not w14626 and not w14627;
w14634 <= not w14632 and not w14633;
w14635 <= w14597 and not w14609;
w14636 <= not w14608 and not w14609;
w14637 <= not w14635 and not w14636;
w14638 <= w14581 and not w14593;
w14639 <= not w14592 and not w14593;
w14640 <= not w14638 and not w14639;
w14641 <= w14303 and w14574;
w14642 <= not w14575 and not w14641;
w14643 <= w3819 and w12824;
w14644 <= w3902 and w12437;
w14645 <= w3981 and w12704;
w14646 <= not w14644 and not w14645;
w14647 <= not w14643 and w14646;
w14648 <= w3985 and w12830;
w14649 <= w14647 and not w14648;
w14650 <= a(26) and not w14649;
w14651 <= a(26) and not w14650;
w14652 <= not w14649 and not w14650;
w14653 <= not w14651 and not w14652;
w14654 <= w14642 and not w14653;
w14655 <= w14642 and not w14654;
w14656 <= not w14653 and not w14654;
w14657 <= not w14655 and not w14656;
w14658 <= not w14387 and w14572;
w14659 <= not w14573 and not w14658;
w14660 <= w3392 and w12440;
w14661 <= w3477 and w12448;
w14662 <= w3541 and w12443;
w14663 <= not w14661 and not w14662;
w14664 <= not w14660 and w14663;
w14665 <= w3303 and not w13986;
w14666 <= w14664 and not w14665;
w14667 <= a(29) and not w14666;
w14668 <= a(29) and not w14667;
w14669 <= not w14666 and not w14667;
w14670 <= not w14668 and not w14669;
w14671 <= w14659 and not w14670;
w14672 <= w14659 and not w14671;
w14673 <= not w14670 and not w14671;
w14674 <= not w14672 and not w14673;
w14675 <= w3819 and w12704;
w14676 <= w3902 and w12305;
w14677 <= w3981 and w12437;
w14678 <= not w14676 and not w14677;
w14679 <= not w14675 and w14678;
w14680 <= w3985 and w12934;
w14681 <= w14679 and not w14680;
w14682 <= a(26) and not w14681;
w14683 <= a(26) and not w14682;
w14684 <= not w14681 and not w14682;
w14685 <= not w14683 and not w14684;
w14686 <= not w14674 and not w14685;
w14687 <= not w14671 and not w14686;
w14688 <= not w14657 and not w14687;
w14689 <= not w14654 and not w14688;
w14690 <= not w14640 and not w14689;
w14691 <= w14640 and w14689;
w14692 <= not w14690 and not w14691;
w14693 <= w4629 and w13450;
w14694 <= w4468 and w13453;
w14695 <= w4539 and w13456;
w14696 <= not w14694 and not w14695;
w14697 <= not w14693 and w14696;
w14698 <= w4471 and w13476;
w14699 <= w14697 and not w14698;
w14700 <= a(23) and not w14699;
w14701 <= a(23) and not w14700;
w14702 <= not w14699 and not w14700;
w14703 <= not w14701 and not w14702;
w14704 <= w14692 and not w14703;
w14705 <= not w14690 and not w14704;
w14706 <= not w14637 and not w14705;
w14707 <= w14637 and w14705;
w14708 <= not w14706 and not w14707;
w14709 <= w5431 and not w13562;
w14710 <= w4870 and w13565;
w14711 <= w5342 and w13568;
w14712 <= not w14710 and not w14711;
w14713 <= not w14709 and w14712;
w14714 <= w4873 and not w13589;
w14715 <= w14713 and not w14714;
w14716 <= a(20) and not w14715;
w14717 <= a(20) and not w14716;
w14718 <= not w14715 and not w14716;
w14719 <= not w14717 and not w14718;
w14720 <= w14708 and not w14719;
w14721 <= not w14706 and not w14720;
w14722 <= w5431 and w13876;
w14723 <= w4870 and w13568;
w14724 <= w5342 and not w13562;
w14725 <= not w14723 and not w14724;
w14726 <= not w14722 and w14725;
w14727 <= w4873 and w14071;
w14728 <= w14726 and not w14727;
w14729 <= a(20) and not w14728;
w14730 <= a(20) and not w14729;
w14731 <= not w14728 and not w14729;
w14732 <= not w14730 and not w14731;
w14733 <= not w14721 and not w14732;
w14734 <= w14282 and w14610;
w14735 <= not w14611 and not w14734;
w14736 <= not w14721 and not w14733;
w14737 <= not w14732 and not w14733;
w14738 <= not w14736 and not w14737;
w14739 <= w14735 and not w14738;
w14740 <= not w14733 and not w14739;
w14741 <= not w14634 and not w14740;
w14742 <= not w14634 and not w14741;
w14743 <= not w14740 and not w14741;
w14744 <= not w14742 and not w14743;
w14745 <= w14692 and not w14704;
w14746 <= not w14703 and not w14704;
w14747 <= not w14745 and not w14746;
w14748 <= w14657 and w14687;
w14749 <= not w14688 and not w14748;
w14750 <= w4629 and w13456;
w14751 <= w4468 and w13426;
w14752 <= w4539 and w13453;
w14753 <= not w14751 and not w14752;
w14754 <= not w14750 and w14753;
w14755 <= w4471 and not w13844;
w14756 <= w14754 and not w14755;
w14757 <= a(23) and not w14756;
w14758 <= a(23) and not w14757;
w14759 <= not w14756 and not w14757;
w14760 <= not w14758 and not w14759;
w14761 <= w14749 and not w14760;
w14762 <= w14749 and not w14761;
w14763 <= not w14760 and not w14761;
w14764 <= not w14762 and not w14763;
w14765 <= not w14674 and not w14686;
w14766 <= not w14685 and not w14686;
w14767 <= not w14765 and not w14766;
w14768 <= not w14549 and not w14551;
w14769 <= not w14451 and w14552;
w14770 <= not w14768 and not w14769;
w14771 <= w12582 and not w12584;
w14772 <= not w12585 and not w14771;
w14773 <= w10 and w14772;
w14774 <= w2955 and w12457;
w14775 <= w2958 and w12463;
w14776 <= w2963 and w12460;
w14777 <= not w14775 and not w14776;
w14778 <= not w14774 and w14777;
w14779 <= not w14773 and w14778;
w14780 <= not w14770 and not w14779;
w14781 <= not w14770 and not w14780;
w14782 <= not w14779 and not w14780;
w14783 <= not w14781 and not w14782;
w14784 <= w3392 and w12446;
w14785 <= w3477 and w12454;
w14786 <= w3541 and w12451;
w14787 <= not w14785 and not w14786;
w14788 <= not w14784 and w14787;
w14789 <= not w3303 and w14788;
w14790 <= w14168 and w14788;
w14791 <= not w14789 and not w14790;
w14792 <= a(29) and not w14791;
w14793 <= not a(29) and w14791;
w14794 <= not w14792 and not w14793;
w14795 <= not w14783 and not w14794;
w14796 <= not w14780 and not w14795;
w14797 <= not w14402 and not w14553;
w14798 <= not w14552 and not w14553;
w14799 <= not w14797 and not w14798;
w14800 <= not w14796 and not w14799;
w14801 <= not w14796 and not w14800;
w14802 <= not w14799 and not w14800;
w14803 <= not w14801 and not w14802;
w14804 <= w3392 and w12448;
w14805 <= w3477 and w12451;
w14806 <= w3541 and w12446;
w14807 <= not w14805 and not w14806;
w14808 <= not w14804 and w14807;
w14809 <= w3303 and w14112;
w14810 <= w14808 and not w14809;
w14811 <= a(29) and not w14810;
w14812 <= a(29) and not w14811;
w14813 <= not w14810 and not w14811;
w14814 <= not w14812 and not w14813;
w14815 <= not w14803 and not w14814;
w14816 <= not w14800 and not w14815;
w14817 <= not w14559 and w14570;
w14818 <= not w14571 and not w14817;
w14819 <= not w14816 and w14818;
w14820 <= w14816 and not w14818;
w14821 <= not w14819 and not w14820;
w14822 <= w3819 and w12437;
w14823 <= w3902 and w12440;
w14824 <= w3981 and w12305;
w14825 <= not w14823 and not w14824;
w14826 <= not w14822 and w14825;
w14827 <= w3985 and not w13671;
w14828 <= w14826 and not w14827;
w14829 <= a(26) and not w14828;
w14830 <= a(26) and not w14829;
w14831 <= not w14828 and not w14829;
w14832 <= not w14830 and not w14831;
w14833 <= w14821 and not w14832;
w14834 <= not w14819 and not w14833;
w14835 <= not w14767 and not w14834;
w14836 <= w14767 and w14834;
w14837 <= not w14835 and not w14836;
w14838 <= w4629 and w13453;
w14839 <= w4468 and w12824;
w14840 <= w4539 and w13426;
w14841 <= not w14839 and not w14840;
w14842 <= not w14838 and w14841;
w14843 <= w4471 and w13519;
w14844 <= w14842 and not w14843;
w14845 <= a(23) and not w14844;
w14846 <= a(23) and not w14845;
w14847 <= not w14844 and not w14845;
w14848 <= not w14846 and not w14847;
w14849 <= w14837 and not w14848;
w14850 <= not w14835 and not w14849;
w14851 <= not w14764 and not w14850;
w14852 <= not w14761 and not w14851;
w14853 <= not w14747 and not w14852;
w14854 <= w14747 and w14852;
w14855 <= not w14853 and not w14854;
w14856 <= w5431 and w13568;
w14857 <= w4870 and w13532;
w14858 <= w5342 and w13565;
w14859 <= not w14857 and not w14858;
w14860 <= not w14856 and w14859;
w14861 <= w4873 and w13864;
w14862 <= w14860 and not w14861;
w14863 <= a(20) and not w14862;
w14864 <= a(20) and not w14863;
w14865 <= not w14862 and not w14863;
w14866 <= not w14864 and not w14865;
w14867 <= w14855 and not w14866;
w14868 <= not w14853 and not w14867;
w14869 <= not w13373 and not w13652;
w14870 <= w5598 and w13876;
w14871 <= not w14869 and not w14870;
w14872 <= not w5601 and w14871;
w14873 <= w13886 and w14871;
w14874 <= not w14872 and not w14873;
w14875 <= a(17) and not w14874;
w14876 <= not a(17) and w14874;
w14877 <= not w14875 and not w14876;
w14878 <= not w14868 and not w14877;
w14879 <= w14708 and not w14720;
w14880 <= not w14719 and not w14720;
w14881 <= not w14879 and not w14880;
w14882 <= w14868 and w14877;
w14883 <= not w14878 and not w14882;
w14884 <= not w14881 and w14883;
w14885 <= not w14878 and not w14884;
w14886 <= not w14735 and w14738;
w14887 <= not w14739 and not w14886;
w14888 <= not w14885 and w14887;
w14889 <= not w14881 and not w14884;
w14890 <= w14883 and not w14884;
w14891 <= not w14889 and not w14890;
w14892 <= w14855 and not w14867;
w14893 <= not w14866 and not w14867;
w14894 <= not w14892 and not w14893;
w14895 <= w14764 and w14850;
w14896 <= not w14851 and not w14895;
w14897 <= w5431 and w13565;
w14898 <= w4870 and w13450;
w14899 <= w5342 and w13532;
w14900 <= not w14898 and not w14899;
w14901 <= not w14897 and w14900;
w14902 <= w4873 and w13911;
w14903 <= w14901 and not w14902;
w14904 <= a(20) and not w14903;
w14905 <= a(20) and not w14904;
w14906 <= not w14903 and not w14904;
w14907 <= not w14905 and not w14906;
w14908 <= w14896 and not w14907;
w14909 <= w14896 and not w14908;
w14910 <= not w14907 and not w14908;
w14911 <= not w14909 and not w14910;
w14912 <= w14837 and not w14849;
w14913 <= not w14848 and not w14849;
w14914 <= not w14912 and not w14913;
w14915 <= w14821 and not w14833;
w14916 <= not w14832 and not w14833;
w14917 <= not w14915 and not w14916;
w14918 <= not w14803 and not w14815;
w14919 <= not w14814 and not w14815;
w14920 <= not w14918 and not w14919;
w14921 <= w3819 and w12305;
w14922 <= w3902 and w12443;
w14923 <= w3981 and w12440;
w14924 <= not w14922 and not w14923;
w14925 <= not w14921 and w14924;
w14926 <= w3985 and not w13683;
w14927 <= w14925 and not w14926;
w14928 <= a(26) and not w14927;
w14929 <= a(26) and not w14928;
w14930 <= not w14927 and not w14928;
w14931 <= not w14929 and not w14930;
w14932 <= not w14920 and not w14931;
w14933 <= not w14920 and not w14932;
w14934 <= not w14931 and not w14932;
w14935 <= not w14933 and not w14934;
w14936 <= not w12574 and not w12577;
w14937 <= not w12575 and w12578;
w14938 <= not w14936 and not w14937;
w14939 <= w10 and not w14938;
w14940 <= w2955 and w12463;
w14941 <= w2958 and w12469;
w14942 <= w2963 and w12466;
w14943 <= not w14941 and not w14942;
w14944 <= not w14940 and w14943;
w14945 <= not w14939 and w14944;
w14946 <= not w602 and w1074;
w14947 <= not w821 and w14946;
w14948 <= w191 and w5108;
w14949 <= w14947 and w14948;
w14950 <= w2028 and w14949;
w14951 <= w1893 and w14950;
w14952 <= w3500 and w14951;
w14953 <= w2673 and w14952;
w14954 <= w122 and w14953;
w14955 <= w2105 and w14954;
w14956 <= w406 and w14955;
w14957 <= w1792 and w14956;
w14958 <= not w362 and w14957;
w14959 <= not w224 and w14958;
w14960 <= not w216 and w14959;
w14961 <= not w492 and w14960;
w14962 <= not w172 and w14961;
w14963 <= not w136 and w14962;
w14964 <= w14494 and not w14963;
w14965 <= not w14494 and w14963;
w14966 <= w10988 and w10989;
w14967 <= not w13373 and not w14966;
w14968 <= a(2) and not w14967;
w14969 <= not a(2) and w14967;
w14970 <= not w14968 and not w14969;
w14971 <= w1673 and w3580;
w14972 <= w1005 and w14971;
w14973 <= w3483 and w14972;
w14974 <= w374 and w14973;
w14975 <= w443 and w14974;
w14976 <= not w103 and w14975;
w14977 <= not w337 and w14976;
w14978 <= not w896 and w14977;
w14979 <= not w105 and w14978;
w14980 <= not w945 and w14979;
w14981 <= not w424 and w14980;
w14982 <= not w706 and w14981;
w14983 <= w2586 and w14414;
w14984 <= not w236 and w14983;
w14985 <= not w164 and w14984;
w14986 <= w3129 and w13762;
w14987 <= w305 and w14986;
w14988 <= w2176 and w14987;
w14989 <= w14985 and w14988;
w14990 <= w12745 and w14989;
w14991 <= w2526 and w14990;
w14992 <= w229 and w14991;
w14993 <= w1716 and w14992;
w14994 <= w14982 and w14993;
w14995 <= w1324 and w14994;
w14996 <= not w352 and w14995;
w14997 <= w72 and w3127;
w14998 <= w6037 and w14997;
w14999 <= w6602 and w14998;
w15000 <= w14316 and w14999;
w15001 <= w12339 and w15000;
w15002 <= w14996 and w15001;
w15003 <= w1458 and w15002;
w15004 <= w182 and w15003;
w15005 <= w3187 and w15004;
w15006 <= not w555 and w15005;
w15007 <= not w287 and w15006;
w15008 <= not w53 and w15007;
w15009 <= not w467 and w15008;
w15010 <= w14970 and not w15009;
w15011 <= not w6 and not w10369;
w15012 <= not w9802 and w15011;
w15013 <= not w9805 and w15012;
w15014 <= not w13373 and not w15013;
w15015 <= not a(5) and w15014;
w15016 <= w14970 and w15009;
w15017 <= not w14970 and not w15009;
w15018 <= not w15016 and not w15017;
w15019 <= a(5) and not w15014;
w15020 <= not w15018 and not w15019;
w15021 <= not w15015 and w15020;
w15022 <= not w15010 and not w15021;
w15023 <= w14494 and not w15022;
w15024 <= not w14494 and w15022;
w15025 <= not w15023 and not w15024;
w15026 <= w2955 and w12469;
w15027 <= w2963 and w12472;
w15028 <= w2958 and w12475;
w15029 <= not w12566 and not w12569;
w15030 <= not w12567 and w12570;
w15031 <= not w15029 and not w15030;
w15032 <= w10 and not w15031;
w15033 <= not w15028 and not w15032;
w15034 <= not w15027 and w15033;
w15035 <= not w15026 and w15034;
w15036 <= w15025 and not w15035;
w15037 <= not w15023 and not w15036;
w15038 <= not w14964 and not w15037;
w15039 <= not w14965 and w15038;
w15040 <= not w14964 and not w15039;
w15041 <= not w14531 and not w14533;
w15042 <= not w14534 and not w15041;
w15043 <= not w15040 and w15042;
w15044 <= w15040 and not w15042;
w15045 <= not w15043 and not w15044;
w15046 <= not w14945 and w15045;
w15047 <= not w15043 and not w15046;
w15048 <= not w14538 and w14547;
w15049 <= not w14548 and not w15048;
w15050 <= not w15047 and w15049;
w15051 <= w15047 and not w15049;
w15052 <= not w15050 and not w15051;
w15053 <= w3392 and w12451;
w15054 <= w3477 and w12457;
w15055 <= w3541 and w12454;
w15056 <= not w15054 and not w15055;
w15057 <= not w15053 and w15056;
w15058 <= not w3303 and w15057;
w15059 <= w14378 and w15057;
w15060 <= not w15058 and not w15059;
w15061 <= a(29) and not w15060;
w15062 <= not a(29) and w15060;
w15063 <= not w15061 and not w15062;
w15064 <= w15052 and not w15063;
w15065 <= not w15050 and not w15064;
w15066 <= w14783 and w14794;
w15067 <= not w14795 and not w15066;
w15068 <= not w15065 and w15067;
w15069 <= w15065 and not w15067;
w15070 <= not w15068 and not w15069;
w15071 <= w3819 and w12440;
w15072 <= w3902 and w12448;
w15073 <= w3981 and w12443;
w15074 <= not w15072 and not w15073;
w15075 <= not w15071 and w15074;
w15076 <= w3985 and not w13986;
w15077 <= w15075 and not w15076;
w15078 <= a(26) and not w15077;
w15079 <= a(26) and not w15078;
w15080 <= not w15077 and not w15078;
w15081 <= not w15079 and not w15080;
w15082 <= w15070 and not w15081;
w15083 <= not w15068 and not w15082;
w15084 <= not w14935 and not w15083;
w15085 <= not w14932 and not w15084;
w15086 <= not w14917 and not w15085;
w15087 <= w14917 and w15085;
w15088 <= not w15086 and not w15087;
w15089 <= w4629 and w13426;
w15090 <= w4468 and w12704;
w15091 <= w4539 and w12824;
w15092 <= not w15090 and not w15091;
w15093 <= not w15089 and w15092;
w15094 <= w4471 and not w13438;
w15095 <= w15093 and not w15094;
w15096 <= a(23) and not w15095;
w15097 <= a(23) and not w15096;
w15098 <= not w15095 and not w15096;
w15099 <= not w15097 and not w15098;
w15100 <= w15088 and not w15099;
w15101 <= not w15086 and not w15100;
w15102 <= not w14914 and not w15101;
w15103 <= w14914 and w15101;
w15104 <= not w15102 and not w15103;
w15105 <= w5431 and w13532;
w15106 <= w4870 and w13456;
w15107 <= w5342 and w13450;
w15108 <= not w15106 and not w15107;
w15109 <= not w15105 and w15108;
w15110 <= w4873 and not w13547;
w15111 <= w15109 and not w15110;
w15112 <= a(20) and not w15111;
w15113 <= a(20) and not w15112;
w15114 <= not w15111 and not w15112;
w15115 <= not w15113 and not w15114;
w15116 <= w15104 and not w15115;
w15117 <= not w15102 and not w15116;
w15118 <= not w14911 and not w15117;
w15119 <= not w14908 and not w15118;
w15120 <= not w14894 and not w15119;
w15121 <= w14894 and w15119;
w15122 <= not w15120 and not w15121;
w15123 <= w6168 and not w13373;
w15124 <= w5598 and not w13562;
w15125 <= w5874 and w13876;
w15126 <= not w15124 and not w15125;
w15127 <= not w15123 and w15126;
w15128 <= w5601 and w13963;
w15129 <= w15127 and not w15128;
w15130 <= a(17) and not w15129;
w15131 <= a(17) and not w15130;
w15132 <= not w15129 and not w15130;
w15133 <= not w15131 and not w15132;
w15134 <= w15122 and not w15133;
w15135 <= not w15120 and not w15134;
w15136 <= not w14891 and not w15135;
w15137 <= w14891 and w15135;
w15138 <= not w15136 and not w15137;
w15139 <= w15122 and not w15134;
w15140 <= not w15133 and not w15134;
w15141 <= not w15139 and not w15140;
w15142 <= w15104 and not w15116;
w15143 <= not w15115 and not w15116;
w15144 <= not w15142 and not w15143;
w15145 <= w15088 and not w15100;
w15146 <= not w15099 and not w15100;
w15147 <= not w15145 and not w15146;
w15148 <= w14935 and w15083;
w15149 <= not w15084 and not w15148;
w15150 <= w4629 and w12824;
w15151 <= w4468 and w12437;
w15152 <= w4539 and w12704;
w15153 <= not w15151 and not w15152;
w15154 <= not w15150 and w15153;
w15155 <= w4471 and w12830;
w15156 <= w15154 and not w15155;
w15157 <= a(23) and not w15156;
w15158 <= a(23) and not w15157;
w15159 <= not w15156 and not w15157;
w15160 <= not w15158 and not w15159;
w15161 <= w15149 and not w15160;
w15162 <= w15149 and not w15161;
w15163 <= not w15160 and not w15161;
w15164 <= not w15162 and not w15163;
w15165 <= w15070 and not w15082;
w15166 <= not w15081 and not w15082;
w15167 <= not w15165 and not w15166;
w15168 <= w15045 and not w15046;
w15169 <= not w14945 and not w15046;
w15170 <= not w15168 and not w15169;
w15171 <= w3392 and w12454;
w15172 <= w3477 and w12460;
w15173 <= w3541 and w12457;
w15174 <= not w15172 and not w15173;
w15175 <= not w15171 and w15174;
w15176 <= w3303 and w14389;
w15177 <= w15175 and not w15176;
w15178 <= a(29) and not w15177;
w15179 <= a(29) and not w15178;
w15180 <= not w15177 and not w15178;
w15181 <= not w15179 and not w15180;
w15182 <= not w15170 and not w15181;
w15183 <= not w15170 and not w15182;
w15184 <= not w15181 and not w15182;
w15185 <= not w15183 and not w15184;
w15186 <= not w15037 and not w15039;
w15187 <= not w14965 and w15040;
w15188 <= not w15186 and not w15187;
w15189 <= w12570 and not w12572;
w15190 <= not w12573 and not w15189;
w15191 <= w10 and w15190;
w15192 <= w2955 and w12466;
w15193 <= w2958 and w12472;
w15194 <= w2963 and w12469;
w15195 <= not w15193 and not w15194;
w15196 <= not w15192 and w15195;
w15197 <= not w15191 and w15196;
w15198 <= not w15188 and not w15197;
w15199 <= not w15188 and not w15198;
w15200 <= not w15197 and not w15198;
w15201 <= not w15199 and not w15200;
w15202 <= w1120 and w2284;
w15203 <= w1829 and w15202;
w15204 <= w3678 and w15203;
w15205 <= w3610 and w15204;
w15206 <= w5720 and w15205;
w15207 <= w2713 and w15206;
w15208 <= w1115 and w15207;
w15209 <= not w404 and w15208;
w15210 <= not w1036 and w15209;
w15211 <= not w448 and w15210;
w15212 <= not w233 and w15211;
w15213 <= not w307 and w15212;
w15214 <= not w92 and w15213;
w15215 <= not w1039 and w15214;
w15216 <= not w527 and w15215;
w15217 <= not w230 and w15216;
w15218 <= not w460 and w15217;
w15219 <= not w14970 and not w15218;
w15220 <= w569 and w13709;
w15221 <= not w263 and w15220;
w15222 <= w12947 and w15221;
w15223 <= w1644 and w15222;
w15224 <= w14996 and w15223;
w15225 <= w438 and w15224;
w15226 <= w447 and w15225;
w15227 <= w1850 and w15226;
w15228 <= w1118 and w15227;
w15229 <= w220 and w15228;
w15230 <= w665 and w15229;
w15231 <= w1718 and w15230;
w15232 <= w137 and w15231;
w15233 <= w4036 and w15232;
w15234 <= not w681 and w15233;
w15235 <= not w174 and w15234;
w15236 <= not w127 and w15235;
w15237 <= not w388 and w15236;
w15238 <= not w818 and w15237;
w15239 <= not w821 and w15238;
w15240 <= not w272 and w15239;
w15241 <= not w14970 and not w15240;
w15242 <= w1492 and w2144;
w15243 <= not w355 and w15242;
w15244 <= not w213 and w15243;
w15245 <= not w370 and w15244;
w15246 <= not w524 and w15245;
w15247 <= not w504 and w15246;
w15248 <= w300 and w1264;
w15249 <= w2403 and w15248;
w15250 <= w12366 and w15249;
w15251 <= w5020 and w15250;
w15252 <= w1660 and w15251;
w15253 <= w15247 and w15252;
w15254 <= w2281 and w15253;
w15255 <= not w86 and w15254;
w15256 <= not w210 and w15255;
w15257 <= not w373 and w15256;
w15258 <= not w1138 and w15257;
w15259 <= not w558 and w15258;
w15260 <= w1627 and w15259;
w15261 <= not w289 and w15260;
w15262 <= not w103 and w15261;
w15263 <= not w231 and w15262;
w15264 <= not w1039 and w15263;
w15265 <= not w467 and w15264;
w15266 <= not w1241 and w3315;
w15267 <= not w681 and w15266;
w15268 <= not w167 and w15267;
w15269 <= not w87 and w15268;
w15270 <= not w138 and w15269;
w15271 <= not w180 and w15270;
w15272 <= not w867 and w15271;
w15273 <= w410 and w1465;
w15274 <= w2744 and w15273;
w15275 <= w1694 and w15274;
w15276 <= w15272 and w15275;
w15277 <= w12908 and w15276;
w15278 <= w15265 and w15277;
w15279 <= w14414 and w15278;
w15280 <= w1172 and w15279;
w15281 <= not w46 and w15280;
w15282 <= not w85 and w15281;
w15283 <= not w506 and w15282;
w15284 <= not w53 and w15283;
w15285 <= not w42 and w15284;
w15286 <= not w221 and w15285;
w15287 <= not w527 and w15286;
w15288 <= not w14970 and not w15287;
w15289 <= not w12550 and not w12553;
w15290 <= not w12551 and w12554;
w15291 <= not w15289 and not w15290;
w15292 <= w10 and not w15291;
w15293 <= w2955 and w12481;
w15294 <= w2958 and w12487;
w15295 <= w2963 and w12484;
w15296 <= not w15294 and not w15295;
w15297 <= not w15293 and w15296;
w15298 <= not w15292 and w15297;
w15299 <= w14970 and w15287;
w15300 <= not w15298 and not w15299;
w15301 <= not w15288 and w15300;
w15302 <= not w15288 and not w15301;
w15303 <= w14970 and w15240;
w15304 <= not w15302 and not w15303;
w15305 <= not w15241 and w15304;
w15306 <= not w15241 and not w15305;
w15307 <= w14970 and w15218;
w15308 <= not w15306 and not w15307;
w15309 <= not w15219 and w15308;
w15310 <= not w15219 and not w15309;
w15311 <= not w15018 and not w15021;
w15312 <= not w15019 and not w15021;
w15313 <= not w15015 and w15312;
w15314 <= not w15311 and not w15313;
w15315 <= not w15310 and w15314;
w15316 <= w15310 and not w15314;
w15317 <= not w15315 and not w15316;
w15318 <= not w12562 and not w12565;
w15319 <= not w12563 and w12566;
w15320 <= not w15318 and not w15319;
w15321 <= w10 and not w15320;
w15322 <= w2955 and w12472;
w15323 <= w2958 and w12478;
w15324 <= w2963 and w12475;
w15325 <= not w15323 and not w15324;
w15326 <= not w15322 and w15325;
w15327 <= not w15321 and w15326;
w15328 <= not w15317 and not w15327;
w15329 <= not w15310 and not w15314;
w15330 <= not w15328 and not w15329;
w15331 <= not w15025 and w15035;
w15332 <= not w15036 and not w15331;
w15333 <= not w15330 and w15332;
w15334 <= w15330 and not w15332;
w15335 <= not w15333 and not w15334;
w15336 <= w3392 and w12460;
w15337 <= w3477 and w12466;
w15338 <= w3541 and w12463;
w15339 <= not w15337 and not w15338;
w15340 <= not w15336 and w15339;
w15341 <= not w3303 and w15340;
w15342 <= not w14543 and w15340;
w15343 <= not w15341 and not w15342;
w15344 <= a(29) and not w15343;
w15345 <= not a(29) and w15343;
w15346 <= not w15344 and not w15345;
w15347 <= w15335 and not w15346;
w15348 <= not w15333 and not w15347;
w15349 <= not w15201 and not w15348;
w15350 <= not w15198 and not w15349;
w15351 <= not w15185 and not w15350;
w15352 <= not w15182 and not w15351;
w15353 <= not w15052 and w15063;
w15354 <= not w15064 and not w15353;
w15355 <= not w15352 and w15354;
w15356 <= w15352 and not w15354;
w15357 <= not w15355 and not w15356;
w15358 <= w3819 and w12443;
w15359 <= w3902 and w12446;
w15360 <= w3981 and w12448;
w15361 <= not w15359 and not w15360;
w15362 <= not w15358 and w15361;
w15363 <= w3985 and w13798;
w15364 <= w15362 and not w15363;
w15365 <= a(26) and not w15364;
w15366 <= a(26) and not w15365;
w15367 <= not w15364 and not w15365;
w15368 <= not w15366 and not w15367;
w15369 <= w15357 and not w15368;
w15370 <= not w15355 and not w15369;
w15371 <= not w15167 and not w15370;
w15372 <= w15167 and w15370;
w15373 <= not w15371 and not w15372;
w15374 <= w4629 and w12704;
w15375 <= w4468 and w12305;
w15376 <= w4539 and w12437;
w15377 <= not w15375 and not w15376;
w15378 <= not w15374 and w15377;
w15379 <= w4471 and w12934;
w15380 <= w15378 and not w15379;
w15381 <= a(23) and not w15380;
w15382 <= a(23) and not w15381;
w15383 <= not w15380 and not w15381;
w15384 <= not w15382 and not w15383;
w15385 <= w15373 and not w15384;
w15386 <= not w15371 and not w15385;
w15387 <= not w15164 and not w15386;
w15388 <= not w15161 and not w15387;
w15389 <= not w15147 and not w15388;
w15390 <= w15147 and w15388;
w15391 <= not w15389 and not w15390;
w15392 <= w5431 and w13450;
w15393 <= w4870 and w13453;
w15394 <= w5342 and w13456;
w15395 <= not w15393 and not w15394;
w15396 <= not w15392 and w15395;
w15397 <= w4873 and w13476;
w15398 <= w15396 and not w15397;
w15399 <= a(20) and not w15398;
w15400 <= a(20) and not w15399;
w15401 <= not w15398 and not w15399;
w15402 <= not w15400 and not w15401;
w15403 <= w15391 and not w15402;
w15404 <= not w15389 and not w15403;
w15405 <= not w15144 and not w15404;
w15406 <= w15144 and w15404;
w15407 <= not w15405 and not w15406;
w15408 <= w6168 and not w13562;
w15409 <= w5598 and w13565;
w15410 <= w5874 and w13568;
w15411 <= not w15409 and not w15410;
w15412 <= not w15408 and w15411;
w15413 <= w5601 and not w13589;
w15414 <= w15412 and not w15413;
w15415 <= a(17) and not w15414;
w15416 <= a(17) and not w15415;
w15417 <= not w15414 and not w15415;
w15418 <= not w15416 and not w15417;
w15419 <= w15407 and not w15418;
w15420 <= not w15405 and not w15419;
w15421 <= w6168 and w13876;
w15422 <= w5598 and w13568;
w15423 <= w5874 and not w13562;
w15424 <= not w15422 and not w15423;
w15425 <= not w15421 and w15424;
w15426 <= w5601 and w14071;
w15427 <= w15425 and not w15426;
w15428 <= a(17) and not w15427;
w15429 <= a(17) and not w15428;
w15430 <= not w15427 and not w15428;
w15431 <= not w15429 and not w15430;
w15432 <= not w15420 and not w15431;
w15433 <= w14911 and w15117;
w15434 <= not w15118 and not w15433;
w15435 <= not w15420 and not w15432;
w15436 <= not w15431 and not w15432;
w15437 <= not w15435 and not w15436;
w15438 <= w15434 and not w15437;
w15439 <= not w15432 and not w15438;
w15440 <= not w15141 and not w15439;
w15441 <= not w15141 and not w15440;
w15442 <= not w15439 and not w15440;
w15443 <= not w15441 and not w15442;
w15444 <= w15391 and not w15403;
w15445 <= not w15402 and not w15403;
w15446 <= not w15444 and not w15445;
w15447 <= w15164 and w15386;
w15448 <= not w15387 and not w15447;
w15449 <= w5431 and w13456;
w15450 <= w4870 and w13426;
w15451 <= w5342 and w13453;
w15452 <= not w15450 and not w15451;
w15453 <= not w15449 and w15452;
w15454 <= w4873 and not w13844;
w15455 <= w15453 and not w15454;
w15456 <= a(20) and not w15455;
w15457 <= a(20) and not w15456;
w15458 <= not w15455 and not w15456;
w15459 <= not w15457 and not w15458;
w15460 <= w15448 and not w15459;
w15461 <= w15448 and not w15460;
w15462 <= not w15459 and not w15460;
w15463 <= not w15461 and not w15462;
w15464 <= w15373 and not w15385;
w15465 <= not w15384 and not w15385;
w15466 <= not w15464 and not w15465;
w15467 <= w15357 and not w15369;
w15468 <= not w15368 and not w15369;
w15469 <= not w15467 and not w15468;
w15470 <= w15185 and w15350;
w15471 <= not w15351 and not w15470;
w15472 <= w3819 and w12448;
w15473 <= w3902 and w12451;
w15474 <= w3981 and w12446;
w15475 <= not w15473 and not w15474;
w15476 <= not w15472 and w15475;
w15477 <= w3985 and w14112;
w15478 <= w15476 and not w15477;
w15479 <= a(26) and not w15478;
w15480 <= a(26) and not w15479;
w15481 <= not w15478 and not w15479;
w15482 <= not w15480 and not w15481;
w15483 <= w15471 and not w15482;
w15484 <= w15471 and not w15483;
w15485 <= not w15482 and not w15483;
w15486 <= not w15484 and not w15485;
w15487 <= w15201 and w15348;
w15488 <= not w15349 and not w15487;
w15489 <= w3392 and w12457;
w15490 <= w3477 and w12463;
w15491 <= w3541 and w12460;
w15492 <= not w15490 and not w15491;
w15493 <= not w15489 and w15492;
w15494 <= w3303 and w14772;
w15495 <= w15493 and not w15494;
w15496 <= a(29) and not w15495;
w15497 <= a(29) and not w15496;
w15498 <= not w15495 and not w15496;
w15499 <= not w15497 and not w15498;
w15500 <= w15488 and not w15499;
w15501 <= w15488 and not w15500;
w15502 <= not w15499 and not w15500;
w15503 <= not w15501 and not w15502;
w15504 <= w3819 and w12446;
w15505 <= w3902 and w12454;
w15506 <= w3981 and w12451;
w15507 <= not w15505 and not w15506;
w15508 <= not w15504 and w15507;
w15509 <= w3985 and not w14168;
w15510 <= w15508 and not w15509;
w15511 <= a(26) and not w15510;
w15512 <= a(26) and not w15511;
w15513 <= not w15510 and not w15511;
w15514 <= not w15512 and not w15513;
w15515 <= not w15503 and not w15514;
w15516 <= not w15500 and not w15515;
w15517 <= not w15486 and not w15516;
w15518 <= not w15483 and not w15517;
w15519 <= not w15469 and not w15518;
w15520 <= w15469 and w15518;
w15521 <= not w15519 and not w15520;
w15522 <= w4629 and w12437;
w15523 <= w4468 and w12440;
w15524 <= w4539 and w12305;
w15525 <= not w15523 and not w15524;
w15526 <= not w15522 and w15525;
w15527 <= w4471 and not w13671;
w15528 <= w15526 and not w15527;
w15529 <= a(23) and not w15528;
w15530 <= a(23) and not w15529;
w15531 <= not w15528 and not w15529;
w15532 <= not w15530 and not w15531;
w15533 <= w15521 and not w15532;
w15534 <= not w15519 and not w15533;
w15535 <= not w15466 and not w15534;
w15536 <= w15466 and w15534;
w15537 <= not w15535 and not w15536;
w15538 <= w5431 and w13453;
w15539 <= w4870 and w12824;
w15540 <= w5342 and w13426;
w15541 <= not w15539 and not w15540;
w15542 <= not w15538 and w15541;
w15543 <= w4873 and w13519;
w15544 <= w15542 and not w15543;
w15545 <= a(20) and not w15544;
w15546 <= a(20) and not w15545;
w15547 <= not w15544 and not w15545;
w15548 <= not w15546 and not w15547;
w15549 <= w15537 and not w15548;
w15550 <= not w15535 and not w15549;
w15551 <= not w15463 and not w15550;
w15552 <= not w15460 and not w15551;
w15553 <= not w15446 and not w15552;
w15554 <= w15446 and w15552;
w15555 <= not w15553 and not w15554;
w15556 <= w6168 and w13568;
w15557 <= w5598 and w13532;
w15558 <= w5874 and w13565;
w15559 <= not w15557 and not w15558;
w15560 <= not w15556 and w15559;
w15561 <= w5601 and w13864;
w15562 <= w15560 and not w15561;
w15563 <= a(17) and not w15562;
w15564 <= a(17) and not w15563;
w15565 <= not w15562 and not w15563;
w15566 <= not w15564 and not w15565;
w15567 <= w15555 and not w15566;
w15568 <= not w15553 and not w15567;
w15569 <= not w13373 and not w13780;
w15570 <= w6337 and w13876;
w15571 <= not w15569 and not w15570;
w15572 <= not w6332 and w15571;
w15573 <= w13886 and w15571;
w15574 <= not w15572 and not w15573;
w15575 <= a(14) and not w15574;
w15576 <= not a(14) and w15574;
w15577 <= not w15575 and not w15576;
w15578 <= not w15568 and not w15577;
w15579 <= w15407 and not w15419;
w15580 <= not w15418 and not w15419;
w15581 <= not w15579 and not w15580;
w15582 <= w15568 and w15577;
w15583 <= not w15578 and not w15582;
w15584 <= not w15581 and w15583;
w15585 <= not w15578 and not w15584;
w15586 <= not w15434 and w15437;
w15587 <= not w15438 and not w15586;
w15588 <= not w15585 and w15587;
w15589 <= not w15581 and not w15584;
w15590 <= w15583 and not w15584;
w15591 <= not w15589 and not w15590;
w15592 <= w15555 and not w15567;
w15593 <= not w15566 and not w15567;
w15594 <= not w15592 and not w15593;
w15595 <= w15463 and w15550;
w15596 <= not w15551 and not w15595;
w15597 <= w6168 and w13565;
w15598 <= w5598 and w13450;
w15599 <= w5874 and w13532;
w15600 <= not w15598 and not w15599;
w15601 <= not w15597 and w15600;
w15602 <= w5601 and w13911;
w15603 <= w15601 and not w15602;
w15604 <= a(17) and not w15603;
w15605 <= a(17) and not w15604;
w15606 <= not w15603 and not w15604;
w15607 <= not w15605 and not w15606;
w15608 <= w15596 and not w15607;
w15609 <= w15596 and not w15608;
w15610 <= not w15607 and not w15608;
w15611 <= not w15609 and not w15610;
w15612 <= w15537 and not w15549;
w15613 <= not w15548 and not w15549;
w15614 <= not w15612 and not w15613;
w15615 <= w15521 and not w15533;
w15616 <= not w15532 and not w15533;
w15617 <= not w15615 and not w15616;
w15618 <= w15486 and w15516;
w15619 <= not w15517 and not w15618;
w15620 <= w4629 and w12305;
w15621 <= w4468 and w12443;
w15622 <= w4539 and w12440;
w15623 <= not w15621 and not w15622;
w15624 <= not w15620 and w15623;
w15625 <= w4471 and not w13683;
w15626 <= w15624 and not w15625;
w15627 <= a(23) and not w15626;
w15628 <= a(23) and not w15627;
w15629 <= not w15626 and not w15627;
w15630 <= not w15628 and not w15629;
w15631 <= w15619 and not w15630;
w15632 <= w15619 and not w15631;
w15633 <= not w15630 and not w15631;
w15634 <= not w15632 and not w15633;
w15635 <= not w15503 and not w15515;
w15636 <= not w15514 and not w15515;
w15637 <= not w15635 and not w15636;
w15638 <= not w15306 and not w15309;
w15639 <= not w15307 and w15310;
w15640 <= not w15638 and not w15639;
w15641 <= not w12558 and not w12561;
w15642 <= not w12559 and w12562;
w15643 <= not w15641 and not w15642;
w15644 <= w10 and not w15643;
w15645 <= w2955 and w12475;
w15646 <= w2958 and w12481;
w15647 <= w2963 and w12478;
w15648 <= not w15646 and not w15647;
w15649 <= not w15645 and w15648;
w15650 <= not w15644 and w15649;
w15651 <= not w15640 and not w15650;
w15652 <= not w15640 and not w15651;
w15653 <= not w15650 and not w15651;
w15654 <= not w15652 and not w15653;
w15655 <= not w15302 and not w15305;
w15656 <= not w15303 and w15306;
w15657 <= not w15655 and not w15656;
w15658 <= w12554 and not w12556;
w15659 <= not w12557 and not w15658;
w15660 <= w10 and w15659;
w15661 <= w2955 and w12478;
w15662 <= w2958 and w12484;
w15663 <= w2963 and w12481;
w15664 <= not w15662 and not w15663;
w15665 <= not w15661 and w15664;
w15666 <= not w15660 and w15665;
w15667 <= not w15657 and not w15666;
w15668 <= not w15657 and not w15667;
w15669 <= not w15666 and not w15667;
w15670 <= not w15668 and not w15669;
w15671 <= not w15298 and not w15301;
w15672 <= not w15299 and w15302;
w15673 <= not w15671 and not w15672;
w15674 <= not w224 and w12765;
w15675 <= not w330 and w15674;
w15676 <= not w108 and w15675;
w15677 <= not w241 and w15676;
w15678 <= not w205 and w15677;
w15679 <= w2719 and w3097;
w15680 <= w2742 and w15679;
w15681 <= w2197 and w15680;
w15682 <= w2026 and w15681;
w15683 <= w623 and w15682;
w15684 <= w4750 and w15683;
w15685 <= w14321 and w15684;
w15686 <= w15678 and w15685;
w15687 <= w223 and w15686;
w15688 <= w291 and w15687;
w15689 <= w51 and w15688;
w15690 <= not w84 and w15689;
w15691 <= not w331 and w15690;
w15692 <= not w102 and w15691;
w15693 <= not w34 and w15692;
w15694 <= not w172 and w15693;
w15695 <= w2955 and w12484;
w15696 <= w2963 and w12487;
w15697 <= w2958 and w12490;
w15698 <= w12546 and not w12548;
w15699 <= not w12549 and not w15698;
w15700 <= w10 and w15699;
w15701 <= not w15697 and not w15700;
w15702 <= not w15696 and w15701;
w15703 <= not w15695 and w15702;
w15704 <= not w15694 and not w15703;
w15705 <= w1008 and w2977;
w15706 <= w2639 and w15705;
w15707 <= w2743 and w15706;
w15708 <= w2357 and w15707;
w15709 <= w13156 and w15708;
w15710 <= w5961 and w15709;
w15711 <= w974 and w15710;
w15712 <= w491 and w15711;
w15713 <= w165 and w15712;
w15714 <= w389 and w15713;
w15715 <= not w236 and w15714;
w15716 <= not w1036 and w15715;
w15717 <= not w651 and w15716;
w15718 <= not w34 and w15717;
w15719 <= not w21 and w15718;
w15720 <= not w364 and w15719;
w15721 <= w2955 and w12487;
w15722 <= w2963 and w12490;
w15723 <= w2958 and w12493;
w15724 <= not w12542 and not w12545;
w15725 <= not w12543 and w12546;
w15726 <= not w15724 and not w15725;
w15727 <= w10 and not w15726;
w15728 <= not w15723 and not w15727;
w15729 <= not w15722 and w15728;
w15730 <= not w15721 and w15729;
w15731 <= not w15720 and not w15730;
w15732 <= w2542 and w3922;
w15733 <= w1539 and w15732;
w15734 <= w1689 and w15733;
w15735 <= w2490 and w15734;
w15736 <= w15265 and w15735;
w15737 <= w809 and w15736;
w15738 <= w1410 and w15737;
w15739 <= w4230 and w15738;
w15740 <= w975 and w15739;
w15741 <= not w216 and w15740;
w15742 <= not w576 and w15741;
w15743 <= not w105 and w15742;
w15744 <= not w592 and w15743;
w15745 <= not w706 and w15744;
w15746 <= w2955 and w12490;
w15747 <= w2963 and w12493;
w15748 <= w2958 and w12496;
w15749 <= not w12538 and not w12541;
w15750 <= not w12539 and w12542;
w15751 <= not w15749 and not w15750;
w15752 <= w10 and not w15751;
w15753 <= not w15748 and not w15752;
w15754 <= not w15747 and w15753;
w15755 <= not w15746 and w15754;
w15756 <= not w15745 and not w15755;
w15757 <= w137 and w812;
w15758 <= not w299 and w15757;
w15759 <= not w274 and w15758;
w15760 <= not w428 and w15759;
w15761 <= not w160 and w15760;
w15762 <= w1207 and w1521;
w15763 <= w12363 and w15762;
w15764 <= w3154 and w15763;
w15765 <= w3350 and w15764;
w15766 <= w6704 and w15765;
w15767 <= w6642 and w15766;
w15768 <= w1851 and w15767;
w15769 <= w1410 and w15768;
w15770 <= w1466 and w15769;
w15771 <= w15761 and w15770;
w15772 <= not w444 and w15771;
w15773 <= not w287 and w15772;
w15774 <= not w396 and w15773;
w15775 <= not w624 and w15774;
w15776 <= not w34 and w15775;
w15777 <= not w212 and w15776;
w15778 <= w2955 and w12493;
w15779 <= w2963 and w12496;
w15780 <= w2958 and w12499;
w15781 <= w12534 and not w12536;
w15782 <= not w12537 and not w15781;
w15783 <= w10 and w15782;
w15784 <= not w15780 and not w15783;
w15785 <= not w15779 and w15784;
w15786 <= not w15778 and w15785;
w15787 <= not w15777 and not w15786;
w15788 <= not w309 and not w440;
w15789 <= not w1138 and w15788;
w15790 <= w1326 and w15789;
w15791 <= w625 and w15790;
w15792 <= w4036 and w15791;
w15793 <= w3094 and w15792;
w15794 <= w6539 and w15793;
w15795 <= w1457 and w15794;
w15796 <= not w537 and w15795;
w15797 <= not w174 and w15796;
w15798 <= not w650 and w15797;
w15799 <= not w102 and w15798;
w15800 <= not w273 and w15799;
w15801 <= not w230 and w15800;
w15802 <= not w184 and w15801;
w15803 <= w2144 and w14453;
w15804 <= w3946 and w15803;
w15805 <= w5125 and w15804;
w15806 <= w6642 and w15805;
w15807 <= w3925 and w15806;
w15808 <= w2508 and w15807;
w15809 <= w872 and w15808;
w15810 <= w128 and w15809;
w15811 <= w505 and w15810;
w15812 <= not w453 and w15811;
w15813 <= not w608 and w15812;
w15814 <= not w62 and w15813;
w15815 <= not w293 and w15814;
w15816 <= not w712 and w12646;
w15817 <= not w16 and w15816;
w15818 <= w1209 and w2677;
w15819 <= w15817 and w15818;
w15820 <= w6452 and w15819;
w15821 <= w14145 and w15820;
w15822 <= w2638 and w15821;
w15823 <= w15815 and w15822;
w15824 <= w1850 and w15823;
w15825 <= w1064 and w15824;
w15826 <= w2518 and w15825;
w15827 <= w137 and w15826;
w15828 <= w15802 and w15827;
w15829 <= not w288 and w15828;
w15830 <= not w86 and w15829;
w15831 <= not w430 and w15830;
w15832 <= not w310 and w15831;
w15833 <= not w1039 and w15832;
w15834 <= not w306 and w15833;
w15835 <= w2955 and w12496;
w15836 <= w2963 and w12499;
w15837 <= w2958 and w12502;
w15838 <= not w12530 and not w12533;
w15839 <= not w12531 and w12534;
w15840 <= not w15838 and not w15839;
w15841 <= w10 and not w15840;
w15842 <= not w15837 and not w15841;
w15843 <= not w15836 and w15842;
w15844 <= not w15835 and w15843;
w15845 <= not w15834 and not w15844;
w15846 <= w12747 and w13184;
w15847 <= w14507 and w15846;
w15848 <= w182 and w15847;
w15849 <= w557 and w15848;
w15850 <= w1199 and w15849;
w15851 <= w1118 and w15850;
w15852 <= w998 and w15851;
w15853 <= w1716 and w15852;
w15854 <= w2402 and w15853;
w15855 <= w569 and w15854;
w15856 <= not w290 and w15855;
w15857 <= not w624 and w15856;
w15858 <= not w726 and w15857;
w15859 <= not w329 and w15858;
w15860 <= w1733 and w2377;
w15861 <= w1957 and w15860;
w15862 <= w12740 and w15861;
w15863 <= w12976 and w15862;
w15864 <= w15859 and w15863;
w15865 <= w666 and w15864;
w15866 <= w913 and w15865;
w15867 <= not w171 and w15866;
w15868 <= not w1181 and w15867;
w15869 <= not w537 and w15868;
w15870 <= not w335 and w15869;
w15871 <= not w127 and w15870;
w15872 <= not w472 and w15871;
w15873 <= not w105 and w15872;
w15874 <= w2955 and w12499;
w15875 <= w2963 and w12502;
w15876 <= w2958 and w12506;
w15877 <= not w12527 and not w12529;
w15878 <= not w12504 and w12530;
w15879 <= not w15877 and not w15878;
w15880 <= w10 and not w15879;
w15881 <= not w15876 and not w15880;
w15882 <= not w15875 and w15881;
w15883 <= not w15874 and w15882;
w15884 <= not w15873 and not w15883;
w15885 <= w3095 and w3326;
w15886 <= not w946 and w15885;
w15887 <= not w103 and w15886;
w15888 <= not w427 and w15887;
w15889 <= not w56 and w13606;
w15890 <= not w760 and w15889;
w15891 <= not w108 and w15890;
w15892 <= w14411 and w15891;
w15893 <= w15888 and w15892;
w15894 <= w406 and w15893;
w15895 <= w944 and w15894;
w15896 <= w2378 and w15895;
w15897 <= w762 and w15896;
w15898 <= not w681 and w15897;
w15899 <= not w89 and w15898;
w15900 <= not w572 and w15899;
w15901 <= not w237 and w15900;
w15902 <= not w209 and w15901;
w15903 <= not w401 and w15902;
w15904 <= not w558 and w15903;
w15905 <= not w298 and w15904;
w15906 <= w1323 and w2127;
w15907 <= w1628 and w15906;
w15908 <= w4754 and w15907;
w15909 <= w394 and w15908;
w15910 <= w1484 and w15909;
w15911 <= w2295 and w15910;
w15912 <= w1066 and w15911;
w15913 <= w15905 and w15912;
w15914 <= w1188 and w15913;
w15915 <= not w70 and w15914;
w15916 <= not w576 and w15915;
w15917 <= not w352 and w15916;
w15918 <= not w431 and w15917;
w15919 <= not w649 and w15918;
w15920 <= w2955 and w12502;
w15921 <= w2963 and w12506;
w15922 <= w2958 and w12509;
w15923 <= w12523 and not w12525;
w15924 <= not w12526 and not w15923;
w15925 <= w10 and w15924;
w15926 <= not w15922 and not w15925;
w15927 <= not w15921 and w15926;
w15928 <= not w15920 and w15927;
w15929 <= not w15919 and not w15928;
w15930 <= w2560 and w3083;
w15931 <= w530 and w15930;
w15932 <= w6500 and w15931;
w15933 <= w5239 and w15932;
w15934 <= w3140 and w15933;
w15935 <= w13145 and w15934;
w15936 <= w13070 and w15935;
w15937 <= w3847 and w15936;
w15938 <= w1851 and w15937;
w15939 <= w2008 and w15938;
w15940 <= not w85 and w15939;
w15941 <= not w498 and w15940;
w15942 <= not w651 and w15941;
w15943 <= not w403 and w15942;
w15944 <= w2955 and w12506;
w15945 <= w2963 and w12509;
w15946 <= w2958 and w12512;
w15947 <= w12519 and not w12521;
w15948 <= not w12522 and not w15947;
w15949 <= w10 and w15948;
w15950 <= not w15946 and not w15949;
w15951 <= not w15945 and w15950;
w15952 <= not w15944 and w15951;
w15953 <= not w15943 and not w15952;
w15954 <= not w85 and not w648;
w15955 <= not w524 and w15954;
w15956 <= w1344 and w15955;
w15957 <= w1038 and w15956;
w15958 <= w812 and w15957;
w15959 <= w743 and w15958;
w15960 <= w1415 and w15959;
w15961 <= w666 and w15960;
w15962 <= not w46 and w15961;
w15963 <= not w262 and w15962;
w15964 <= not w365 and w15963;
w15965 <= not w228 and w15964;
w15966 <= not w364 and w15965;
w15967 <= w2927 and w12720;
w15968 <= w593 and w15967;
w15969 <= w3344 and w15968;
w15970 <= w15966 and w15969;
w15971 <= w14433 and w15970;
w15972 <= w15272 and w15971;
w15973 <= w5020 and w15972;
w15974 <= w1182 and w15973;
w15975 <= w353 and w15974;
w15976 <= not w263 and w15975;
w15977 <= not w446 and w15976;
w15978 <= not w82 and w15977;
w15979 <= not w227 and w15978;
w15980 <= not w448 and w15979;
w15981 <= not w330 and w15980;
w15982 <= not w651 and w15981;
w15983 <= not w371 and w15982;
w15984 <= not w157 and w15983;
w15985 <= w1095 and w2126;
w15986 <= not w687 and w15985;
w15987 <= not w174 and w15986;
w15988 <= not w81 and w15987;
w15989 <= not w387 and w15988;
w15990 <= not w96 and w15989;
w15991 <= w1942 and w3063;
w15992 <= w13203 and w15991;
w15993 <= w3840 and w15992;
w15994 <= w725 and w15993;
w15995 <= w15761 and w15994;
w15996 <= w15990 and w15995;
w15997 <= w217 and w15996;
w15998 <= w762 and w15997;
w15999 <= not w42 and w15998;
w16000 <= not w261 and w15999;
w16001 <= not w16 and w16000;
w16002 <= not w166 and w16001;
w16003 <= w1344 and w1579;
w16004 <= w2376 and w16003;
w16005 <= w2107 and w16004;
w16006 <= w3706 and w16005;
w16007 <= w2007 and w16006;
w16008 <= w6597 and w16007;
w16009 <= w2047 and w16008;
w16010 <= w2281 and w16009;
w16011 <= w16002 and w16010;
w16012 <= not w681 and w16011;
w16013 <= not w227 and w16012;
w16014 <= not w127 and w16013;
w16015 <= not w108 and w16014;
w16016 <= not w371 and w16015;
w16017 <= w2955 and w12512;
w16018 <= w12512 and w12516;
w16019 <= not w12512 and not w12516;
w16020 <= not w16018 and not w16019;
w16021 <= w10 and not w16020;
w16022 <= w2963 and not w12516;
w16023 <= not w16021 and not w16022;
w16024 <= not w16017 and w16023;
w16025 <= not w16016 and not w16024;
w16026 <= not w15984 and w16025;
w16027 <= not w12509 and w16018;
w16028 <= w12509 and not w16018;
w16029 <= not w16027 and not w16028;
w16030 <= w10 and not w16029;
w16031 <= w2955 and w12509;
w16032 <= w2958 and not w12516;
w16033 <= w2963 and w12512;
w16034 <= not w16032 and not w16033;
w16035 <= not w16031 and w16034;
w16036 <= not w16030 and w16035;
w16037 <= w15984 and not w16025;
w16038 <= not w16026 and not w16037;
w16039 <= not w16036 and w16038;
w16040 <= not w16026 and not w16039;
w16041 <= not w15943 and not w15953;
w16042 <= not w15952 and not w15953;
w16043 <= not w16041 and not w16042;
w16044 <= not w16040 and not w16043;
w16045 <= not w15953 and not w16044;
w16046 <= not w15919 and not w15929;
w16047 <= not w15928 and not w15929;
w16048 <= not w16046 and not w16047;
w16049 <= not w16045 and not w16048;
w16050 <= not w15929 and not w16049;
w16051 <= not w15873 and not w15884;
w16052 <= not w15883 and not w15884;
w16053 <= not w16051 and not w16052;
w16054 <= not w16050 and not w16053;
w16055 <= not w15884 and not w16054;
w16056 <= not w15834 and not w15845;
w16057 <= not w15844 and not w15845;
w16058 <= not w16056 and not w16057;
w16059 <= not w16055 and not w16058;
w16060 <= not w15845 and not w16059;
w16061 <= not w15777 and not w15787;
w16062 <= not w15786 and not w15787;
w16063 <= not w16061 and not w16062;
w16064 <= not w16060 and not w16063;
w16065 <= not w15787 and not w16064;
w16066 <= not w15745 and not w15756;
w16067 <= not w15755 and not w15756;
w16068 <= not w16066 and not w16067;
w16069 <= not w16065 and not w16068;
w16070 <= not w15756 and not w16069;
w16071 <= not w15720 and not w15731;
w16072 <= not w15730 and not w15731;
w16073 <= not w16071 and not w16072;
w16074 <= not w16070 and not w16073;
w16075 <= not w15731 and not w16074;
w16076 <= not w15694 and not w15704;
w16077 <= not w15703 and not w15704;
w16078 <= not w16076 and not w16077;
w16079 <= not w16075 and not w16078;
w16080 <= not w15704 and not w16079;
w16081 <= not w15673 and not w16080;
w16082 <= w15673 and w16080;
w16083 <= not w16081 and not w16082;
w16084 <= w3392 and w12472;
w16085 <= w3477 and w12478;
w16086 <= w3541 and w12475;
w16087 <= not w16085 and not w16086;
w16088 <= not w16084 and w16087;
w16089 <= not w3303 and w16088;
w16090 <= w15320 and w16088;
w16091 <= not w16089 and not w16090;
w16092 <= a(29) and not w16091;
w16093 <= not a(29) and w16091;
w16094 <= not w16092 and not w16093;
w16095 <= w16083 and not w16094;
w16096 <= not w16081 and not w16095;
w16097 <= not w15670 and not w16096;
w16098 <= not w15667 and not w16097;
w16099 <= not w15654 and not w16098;
w16100 <= not w15651 and not w16099;
w16101 <= w15317 and w15327;
w16102 <= not w15328 and not w16101;
w16103 <= not w16100 and w16102;
w16104 <= w16100 and not w16102;
w16105 <= not w16103 and not w16104;
w16106 <= w3392 and w12463;
w16107 <= w3477 and w12469;
w16108 <= w3541 and w12466;
w16109 <= not w16107 and not w16108;
w16110 <= not w16106 and w16109;
w16111 <= w3303 and not w14938;
w16112 <= w16110 and not w16111;
w16113 <= a(29) and not w16112;
w16114 <= a(29) and not w16113;
w16115 <= not w16112 and not w16113;
w16116 <= not w16114 and not w16115;
w16117 <= w16105 and not w16116;
w16118 <= not w16103 and not w16117;
w16119 <= not w15335 and w15346;
w16120 <= not w15347 and not w16119;
w16121 <= not w16118 and w16120;
w16122 <= w16118 and not w16120;
w16123 <= not w16121 and not w16122;
w16124 <= w3819 and w12451;
w16125 <= w3902 and w12457;
w16126 <= w3981 and w12454;
w16127 <= not w16125 and not w16126;
w16128 <= not w16124 and w16127;
w16129 <= w3985 and not w14378;
w16130 <= w16128 and not w16129;
w16131 <= a(26) and not w16130;
w16132 <= a(26) and not w16131;
w16133 <= not w16130 and not w16131;
w16134 <= not w16132 and not w16133;
w16135 <= w16123 and not w16134;
w16136 <= not w16121 and not w16135;
w16137 <= not w15637 and not w16136;
w16138 <= w15637 and w16136;
w16139 <= not w16137 and not w16138;
w16140 <= w4629 and w12440;
w16141 <= w4468 and w12448;
w16142 <= w4539 and w12443;
w16143 <= not w16141 and not w16142;
w16144 <= not w16140 and w16143;
w16145 <= w4471 and not w13986;
w16146 <= w16144 and not w16145;
w16147 <= a(23) and not w16146;
w16148 <= a(23) and not w16147;
w16149 <= not w16146 and not w16147;
w16150 <= not w16148 and not w16149;
w16151 <= w16139 and not w16150;
w16152 <= not w16137 and not w16151;
w16153 <= not w15634 and not w16152;
w16154 <= not w15631 and not w16153;
w16155 <= not w15617 and not w16154;
w16156 <= w15617 and w16154;
w16157 <= not w16155 and not w16156;
w16158 <= w5431 and w13426;
w16159 <= w4870 and w12704;
w16160 <= w5342 and w12824;
w16161 <= not w16159 and not w16160;
w16162 <= not w16158 and w16161;
w16163 <= w4873 and not w13438;
w16164 <= w16162 and not w16163;
w16165 <= a(20) and not w16164;
w16166 <= a(20) and not w16165;
w16167 <= not w16164 and not w16165;
w16168 <= not w16166 and not w16167;
w16169 <= w16157 and not w16168;
w16170 <= not w16155 and not w16169;
w16171 <= not w15614 and not w16170;
w16172 <= w15614 and w16170;
w16173 <= not w16171 and not w16172;
w16174 <= w6168 and w13532;
w16175 <= w5598 and w13456;
w16176 <= w5874 and w13450;
w16177 <= not w16175 and not w16176;
w16178 <= not w16174 and w16177;
w16179 <= w5601 and not w13547;
w16180 <= w16178 and not w16179;
w16181 <= a(17) and not w16180;
w16182 <= a(17) and not w16181;
w16183 <= not w16180 and not w16181;
w16184 <= not w16182 and not w16183;
w16185 <= w16173 and not w16184;
w16186 <= not w16171 and not w16185;
w16187 <= not w15611 and not w16186;
w16188 <= not w15608 and not w16187;
w16189 <= not w15594 and not w16188;
w16190 <= w15594 and w16188;
w16191 <= not w16189 and not w16190;
w16192 <= w7036 and not w13373;
w16193 <= w6337 and not w13562;
w16194 <= w6886 and w13876;
w16195 <= not w16193 and not w16194;
w16196 <= not w16192 and w16195;
w16197 <= w6332 and w13963;
w16198 <= w16196 and not w16197;
w16199 <= a(14) and not w16198;
w16200 <= a(14) and not w16199;
w16201 <= not w16198 and not w16199;
w16202 <= not w16200 and not w16201;
w16203 <= w16191 and not w16202;
w16204 <= not w16189 and not w16203;
w16205 <= not w15591 and not w16204;
w16206 <= w15591 and w16204;
w16207 <= not w16205 and not w16206;
w16208 <= w16191 and not w16203;
w16209 <= not w16202 and not w16203;
w16210 <= not w16208 and not w16209;
w16211 <= w16173 and not w16185;
w16212 <= not w16184 and not w16185;
w16213 <= not w16211 and not w16212;
w16214 <= w16157 and not w16169;
w16215 <= not w16168 and not w16169;
w16216 <= not w16214 and not w16215;
w16217 <= w15634 and w16152;
w16218 <= not w16153 and not w16217;
w16219 <= w5431 and w12824;
w16220 <= w4870 and w12437;
w16221 <= w5342 and w12704;
w16222 <= not w16220 and not w16221;
w16223 <= not w16219 and w16222;
w16224 <= w4873 and w12830;
w16225 <= w16223 and not w16224;
w16226 <= a(20) and not w16225;
w16227 <= a(20) and not w16226;
w16228 <= not w16225 and not w16226;
w16229 <= not w16227 and not w16228;
w16230 <= w16218 and not w16229;
w16231 <= w16218 and not w16230;
w16232 <= not w16229 and not w16230;
w16233 <= not w16231 and not w16232;
w16234 <= w16139 and not w16151;
w16235 <= not w16150 and not w16151;
w16236 <= not w16234 and not w16235;
w16237 <= w16123 and not w16135;
w16238 <= not w16134 and not w16135;
w16239 <= not w16237 and not w16238;
w16240 <= w16105 and not w16117;
w16241 <= not w16116 and not w16117;
w16242 <= not w16240 and not w16241;
w16243 <= w3819 and w12454;
w16244 <= w3902 and w12460;
w16245 <= w3981 and w12457;
w16246 <= not w16244 and not w16245;
w16247 <= not w16243 and w16246;
w16248 <= w3985 and w14389;
w16249 <= w16247 and not w16248;
w16250 <= a(26) and not w16249;
w16251 <= a(26) and not w16250;
w16252 <= not w16249 and not w16250;
w16253 <= not w16251 and not w16252;
w16254 <= not w16242 and not w16253;
w16255 <= not w16242 and not w16254;
w16256 <= not w16253 and not w16254;
w16257 <= not w16255 and not w16256;
w16258 <= w15654 and w16098;
w16259 <= not w16099 and not w16258;
w16260 <= w3392 and w12466;
w16261 <= w3477 and w12472;
w16262 <= w3541 and w12469;
w16263 <= not w16261 and not w16262;
w16264 <= not w16260 and w16263;
w16265 <= w3303 and w15190;
w16266 <= w16264 and not w16265;
w16267 <= a(29) and not w16266;
w16268 <= a(29) and not w16267;
w16269 <= not w16266 and not w16267;
w16270 <= not w16268 and not w16269;
w16271 <= w16259 and not w16270;
w16272 <= w16259 and not w16271;
w16273 <= not w16270 and not w16271;
w16274 <= not w16272 and not w16273;
w16275 <= w3902 and w12463;
w16276 <= w3981 and w12460;
w16277 <= w3819 and w12457;
w16278 <= not w16276 and not w16277;
w16279 <= not w16275 and w16278;
w16280 <= w3985 and w14772;
w16281 <= w16279 and not w16280;
w16282 <= a(26) and not w16281;
w16283 <= a(26) and not w16282;
w16284 <= not w16281 and not w16282;
w16285 <= not w16283 and not w16284;
w16286 <= not w16274 and not w16285;
w16287 <= not w16271 and not w16286;
w16288 <= not w16257 and not w16287;
w16289 <= not w16254 and not w16288;
w16290 <= not w16239 and not w16289;
w16291 <= w16239 and w16289;
w16292 <= not w16290 and not w16291;
w16293 <= w4629 and w12443;
w16294 <= w4468 and w12446;
w16295 <= w4539 and w12448;
w16296 <= not w16294 and not w16295;
w16297 <= not w16293 and w16296;
w16298 <= w4471 and w13798;
w16299 <= w16297 and not w16298;
w16300 <= a(23) and not w16299;
w16301 <= a(23) and not w16300;
w16302 <= not w16299 and not w16300;
w16303 <= not w16301 and not w16302;
w16304 <= w16292 and not w16303;
w16305 <= not w16290 and not w16304;
w16306 <= not w16236 and not w16305;
w16307 <= w16236 and w16305;
w16308 <= not w16306 and not w16307;
w16309 <= w5431 and w12704;
w16310 <= w4870 and w12305;
w16311 <= w5342 and w12437;
w16312 <= not w16310 and not w16311;
w16313 <= not w16309 and w16312;
w16314 <= w4873 and w12934;
w16315 <= w16313 and not w16314;
w16316 <= a(20) and not w16315;
w16317 <= a(20) and not w16316;
w16318 <= not w16315 and not w16316;
w16319 <= not w16317 and not w16318;
w16320 <= w16308 and not w16319;
w16321 <= not w16306 and not w16320;
w16322 <= not w16233 and not w16321;
w16323 <= not w16230 and not w16322;
w16324 <= not w16216 and not w16323;
w16325 <= w16216 and w16323;
w16326 <= not w16324 and not w16325;
w16327 <= w6168 and w13450;
w16328 <= w5598 and w13453;
w16329 <= w5874 and w13456;
w16330 <= not w16328 and not w16329;
w16331 <= not w16327 and w16330;
w16332 <= w5601 and w13476;
w16333 <= w16331 and not w16332;
w16334 <= a(17) and not w16333;
w16335 <= a(17) and not w16334;
w16336 <= not w16333 and not w16334;
w16337 <= not w16335 and not w16336;
w16338 <= w16326 and not w16337;
w16339 <= not w16324 and not w16338;
w16340 <= not w16213 and not w16339;
w16341 <= w16213 and w16339;
w16342 <= not w16340 and not w16341;
w16343 <= w7036 and not w13562;
w16344 <= w6337 and w13565;
w16345 <= w6886 and w13568;
w16346 <= not w16344 and not w16345;
w16347 <= not w16343 and w16346;
w16348 <= w6332 and not w13589;
w16349 <= w16347 and not w16348;
w16350 <= a(14) and not w16349;
w16351 <= a(14) and not w16350;
w16352 <= not w16349 and not w16350;
w16353 <= not w16351 and not w16352;
w16354 <= w16342 and not w16353;
w16355 <= not w16340 and not w16354;
w16356 <= w7036 and w13876;
w16357 <= w6337 and w13568;
w16358 <= w6886 and not w13562;
w16359 <= not w16357 and not w16358;
w16360 <= not w16356 and w16359;
w16361 <= w6332 and w14071;
w16362 <= w16360 and not w16361;
w16363 <= a(14) and not w16362;
w16364 <= a(14) and not w16363;
w16365 <= not w16362 and not w16363;
w16366 <= not w16364 and not w16365;
w16367 <= not w16355 and not w16366;
w16368 <= w15611 and w16186;
w16369 <= not w16187 and not w16368;
w16370 <= not w16355 and not w16367;
w16371 <= not w16366 and not w16367;
w16372 <= not w16370 and not w16371;
w16373 <= w16369 and not w16372;
w16374 <= not w16367 and not w16373;
w16375 <= not w16210 and not w16374;
w16376 <= not w16210 and not w16375;
w16377 <= not w16374 and not w16375;
w16378 <= not w16376 and not w16377;
w16379 <= w16326 and not w16338;
w16380 <= not w16337 and not w16338;
w16381 <= not w16379 and not w16380;
w16382 <= w16233 and w16321;
w16383 <= not w16322 and not w16382;
w16384 <= w6168 and w13456;
w16385 <= w5598 and w13426;
w16386 <= w5874 and w13453;
w16387 <= not w16385 and not w16386;
w16388 <= not w16384 and w16387;
w16389 <= w5601 and not w13844;
w16390 <= w16388 and not w16389;
w16391 <= a(17) and not w16390;
w16392 <= a(17) and not w16391;
w16393 <= not w16390 and not w16391;
w16394 <= not w16392 and not w16393;
w16395 <= w16383 and not w16394;
w16396 <= w16383 and not w16395;
w16397 <= not w16394 and not w16395;
w16398 <= not w16396 and not w16397;
w16399 <= w16308 and not w16320;
w16400 <= not w16319 and not w16320;
w16401 <= not w16399 and not w16400;
w16402 <= w16292 and not w16304;
w16403 <= not w16303 and not w16304;
w16404 <= not w16402 and not w16403;
w16405 <= w16257 and w16287;
w16406 <= not w16288 and not w16405;
w16407 <= w4629 and w12448;
w16408 <= w4468 and w12451;
w16409 <= w4539 and w12446;
w16410 <= not w16408 and not w16409;
w16411 <= not w16407 and w16410;
w16412 <= w4471 and w14112;
w16413 <= w16411 and not w16412;
w16414 <= a(23) and not w16413;
w16415 <= a(23) and not w16414;
w16416 <= not w16413 and not w16414;
w16417 <= not w16415 and not w16416;
w16418 <= w16406 and not w16417;
w16419 <= w16406 and not w16418;
w16420 <= not w16417 and not w16418;
w16421 <= not w16419 and not w16420;
w16422 <= not w16274 and not w16286;
w16423 <= not w16285 and not w16286;
w16424 <= not w16422 and not w16423;
w16425 <= w15670 and w16096;
w16426 <= not w16097 and not w16425;
w16427 <= w3392 and w12469;
w16428 <= w3477 and w12475;
w16429 <= w3541 and w12472;
w16430 <= not w16428 and not w16429;
w16431 <= not w16427 and w16430;
w16432 <= w3303 and not w15031;
w16433 <= w16431 and not w16432;
w16434 <= a(29) and not w16433;
w16435 <= a(29) and not w16434;
w16436 <= not w16433 and not w16434;
w16437 <= not w16435 and not w16436;
w16438 <= w16426 and not w16437;
w16439 <= w16426 and not w16438;
w16440 <= not w16437 and not w16438;
w16441 <= not w16439 and not w16440;
w16442 <= w3981 and w12463;
w16443 <= w3819 and w12460;
w16444 <= w3902 and w12466;
w16445 <= not w16443 and not w16444;
w16446 <= not w16442 and w16445;
w16447 <= w3985 and w14543;
w16448 <= w16446 and not w16447;
w16449 <= a(26) and not w16448;
w16450 <= a(26) and not w16449;
w16451 <= not w16448 and not w16449;
w16452 <= not w16450 and not w16451;
w16453 <= not w16441 and not w16452;
w16454 <= not w16438 and not w16453;
w16455 <= not w16424 and not w16454;
w16456 <= w16424 and w16454;
w16457 <= not w16455 and not w16456;
w16458 <= w4629 and w12446;
w16459 <= w4468 and w12454;
w16460 <= w4539 and w12451;
w16461 <= not w16459 and not w16460;
w16462 <= not w16458 and w16461;
w16463 <= w4471 and not w14168;
w16464 <= w16462 and not w16463;
w16465 <= a(23) and not w16464;
w16466 <= a(23) and not w16465;
w16467 <= not w16464 and not w16465;
w16468 <= not w16466 and not w16467;
w16469 <= w16457 and not w16468;
w16470 <= not w16455 and not w16469;
w16471 <= not w16421 and not w16470;
w16472 <= not w16418 and not w16471;
w16473 <= not w16404 and not w16472;
w16474 <= w16404 and w16472;
w16475 <= not w16473 and not w16474;
w16476 <= w5431 and w12437;
w16477 <= w4870 and w12440;
w16478 <= w5342 and w12305;
w16479 <= not w16477 and not w16478;
w16480 <= not w16476 and w16479;
w16481 <= w4873 and not w13671;
w16482 <= w16480 and not w16481;
w16483 <= a(20) and not w16482;
w16484 <= a(20) and not w16483;
w16485 <= not w16482 and not w16483;
w16486 <= not w16484 and not w16485;
w16487 <= w16475 and not w16486;
w16488 <= not w16473 and not w16487;
w16489 <= not w16401 and not w16488;
w16490 <= w16401 and w16488;
w16491 <= not w16489 and not w16490;
w16492 <= w6168 and w13453;
w16493 <= w5598 and w12824;
w16494 <= w5874 and w13426;
w16495 <= not w16493 and not w16494;
w16496 <= not w16492 and w16495;
w16497 <= w5601 and w13519;
w16498 <= w16496 and not w16497;
w16499 <= a(17) and not w16498;
w16500 <= a(17) and not w16499;
w16501 <= not w16498 and not w16499;
w16502 <= not w16500 and not w16501;
w16503 <= w16491 and not w16502;
w16504 <= not w16489 and not w16503;
w16505 <= not w16398 and not w16504;
w16506 <= not w16395 and not w16505;
w16507 <= not w16381 and not w16506;
w16508 <= w16381 and w16506;
w16509 <= not w16507 and not w16508;
w16510 <= w7036 and w13568;
w16511 <= w6337 and w13532;
w16512 <= w6886 and w13565;
w16513 <= not w16511 and not w16512;
w16514 <= not w16510 and w16513;
w16515 <= w6332 and w13864;
w16516 <= w16514 and not w16515;
w16517 <= a(14) and not w16516;
w16518 <= a(14) and not w16517;
w16519 <= not w16516 and not w16517;
w16520 <= not w16518 and not w16519;
w16521 <= w16509 and not w16520;
w16522 <= not w16507 and not w16521;
w16523 <= not w13373 and not w14359;
w16524 <= w7226 and w13876;
w16525 <= not w16523 and not w16524;
w16526 <= not w7229 and w16525;
w16527 <= w13886 and w16525;
w16528 <= not w16526 and not w16527;
w16529 <= a(11) and not w16528;
w16530 <= not a(11) and w16528;
w16531 <= not w16529 and not w16530;
w16532 <= not w16522 and not w16531;
w16533 <= w16342 and not w16354;
w16534 <= not w16353 and not w16354;
w16535 <= not w16533 and not w16534;
w16536 <= w16522 and w16531;
w16537 <= not w16532 and not w16536;
w16538 <= not w16535 and w16537;
w16539 <= not w16532 and not w16538;
w16540 <= not w16369 and w16372;
w16541 <= not w16373 and not w16540;
w16542 <= not w16539 and w16541;
w16543 <= not w16535 and not w16538;
w16544 <= w16537 and not w16538;
w16545 <= not w16543 and not w16544;
w16546 <= w16509 and not w16521;
w16547 <= not w16520 and not w16521;
w16548 <= not w16546 and not w16547;
w16549 <= w16398 and w16504;
w16550 <= not w16505 and not w16549;
w16551 <= w7036 and w13565;
w16552 <= w6337 and w13450;
w16553 <= w6886 and w13532;
w16554 <= not w16552 and not w16553;
w16555 <= not w16551 and w16554;
w16556 <= w6332 and w13911;
w16557 <= w16555 and not w16556;
w16558 <= a(14) and not w16557;
w16559 <= a(14) and not w16558;
w16560 <= not w16557 and not w16558;
w16561 <= not w16559 and not w16560;
w16562 <= w16550 and not w16561;
w16563 <= w16550 and not w16562;
w16564 <= not w16561 and not w16562;
w16565 <= not w16563 and not w16564;
w16566 <= w16491 and not w16503;
w16567 <= not w16502 and not w16503;
w16568 <= not w16566 and not w16567;
w16569 <= w16475 and not w16487;
w16570 <= not w16486 and not w16487;
w16571 <= not w16569 and not w16570;
w16572 <= w16421 and w16470;
w16573 <= not w16471 and not w16572;
w16574 <= w5431 and w12305;
w16575 <= w4870 and w12443;
w16576 <= w5342 and w12440;
w16577 <= not w16575 and not w16576;
w16578 <= not w16574 and w16577;
w16579 <= w4873 and not w13683;
w16580 <= w16578 and not w16579;
w16581 <= a(20) and not w16580;
w16582 <= a(20) and not w16581;
w16583 <= not w16580 and not w16581;
w16584 <= not w16582 and not w16583;
w16585 <= w16573 and not w16584;
w16586 <= w16573 and not w16585;
w16587 <= not w16584 and not w16585;
w16588 <= not w16586 and not w16587;
w16589 <= w16457 and not w16469;
w16590 <= not w16468 and not w16469;
w16591 <= not w16589 and not w16590;
w16592 <= not w16441 and not w16453;
w16593 <= not w16452 and not w16453;
w16594 <= not w16592 and not w16593;
w16595 <= not w16075 and not w16079;
w16596 <= not w16078 and not w16079;
w16597 <= not w16595 and not w16596;
w16598 <= w3392 and w12475;
w16599 <= w3477 and w12481;
w16600 <= w3541 and w12478;
w16601 <= not w16599 and not w16600;
w16602 <= not w16598 and w16601;
w16603 <= not w3303 and w16602;
w16604 <= w15643 and w16602;
w16605 <= not w16603 and not w16604;
w16606 <= a(29) and not w16605;
w16607 <= not a(29) and w16605;
w16608 <= not w16606 and not w16607;
w16609 <= not w16597 and not w16608;
w16610 <= not w16070 and not w16074;
w16611 <= not w16073 and not w16074;
w16612 <= not w16610 and not w16611;
w16613 <= w3392 and w12478;
w16614 <= w3477 and w12484;
w16615 <= w3541 and w12481;
w16616 <= not w16614 and not w16615;
w16617 <= not w16613 and w16616;
w16618 <= not w3303 and w16617;
w16619 <= not w15659 and w16617;
w16620 <= not w16618 and not w16619;
w16621 <= a(29) and not w16620;
w16622 <= not a(29) and w16620;
w16623 <= not w16621 and not w16622;
w16624 <= not w16612 and not w16623;
w16625 <= not w16065 and not w16069;
w16626 <= not w16068 and not w16069;
w16627 <= not w16625 and not w16626;
w16628 <= w3392 and w12481;
w16629 <= w3477 and w12487;
w16630 <= w3541 and w12484;
w16631 <= not w16629 and not w16630;
w16632 <= not w16628 and w16631;
w16633 <= not w3303 and w16632;
w16634 <= w15291 and w16632;
w16635 <= not w16633 and not w16634;
w16636 <= a(29) and not w16635;
w16637 <= not a(29) and w16635;
w16638 <= not w16636 and not w16637;
w16639 <= not w16627 and not w16638;
w16640 <= not w16060 and not w16064;
w16641 <= not w16063 and not w16064;
w16642 <= not w16640 and not w16641;
w16643 <= w3392 and w12484;
w16644 <= w3477 and w12490;
w16645 <= w3541 and w12487;
w16646 <= not w16644 and not w16645;
w16647 <= not w16643 and w16646;
w16648 <= not w3303 and w16647;
w16649 <= not w15699 and w16647;
w16650 <= not w16648 and not w16649;
w16651 <= a(29) and not w16650;
w16652 <= not a(29) and w16650;
w16653 <= not w16651 and not w16652;
w16654 <= not w16642 and not w16653;
w16655 <= not w16055 and not w16059;
w16656 <= not w16058 and not w16059;
w16657 <= not w16655 and not w16656;
w16658 <= w3392 and w12487;
w16659 <= w3477 and w12493;
w16660 <= w3541 and w12490;
w16661 <= not w16659 and not w16660;
w16662 <= not w16658 and w16661;
w16663 <= not w3303 and w16662;
w16664 <= w15726 and w16662;
w16665 <= not w16663 and not w16664;
w16666 <= a(29) and not w16665;
w16667 <= not a(29) and w16665;
w16668 <= not w16666 and not w16667;
w16669 <= not w16657 and not w16668;
w16670 <= w3392 and w12490;
w16671 <= w3477 and w12496;
w16672 <= w3541 and w12493;
w16673 <= not w16671 and not w16672;
w16674 <= not w16670 and w16673;
w16675 <= w3303 and not w15751;
w16676 <= w16674 and not w16675;
w16677 <= a(29) and not w16676;
w16678 <= not w16676 and not w16677;
w16679 <= a(29) and not w16677;
w16680 <= not w16678 and not w16679;
w16681 <= not w16050 and not w16054;
w16682 <= not w16053 and not w16054;
w16683 <= not w16681 and not w16682;
w16684 <= not w16680 and not w16683;
w16685 <= not w16680 and not w16684;
w16686 <= not w16683 and not w16684;
w16687 <= not w16685 and not w16686;
w16688 <= w3392 and w12493;
w16689 <= w3477 and w12499;
w16690 <= w3541 and w12496;
w16691 <= not w16689 and not w16690;
w16692 <= not w16688 and w16691;
w16693 <= w3303 and w15782;
w16694 <= w16692 and not w16693;
w16695 <= a(29) and not w16694;
w16696 <= not w16694 and not w16695;
w16697 <= a(29) and not w16695;
w16698 <= not w16696 and not w16697;
w16699 <= not w16045 and not w16049;
w16700 <= not w16048 and not w16049;
w16701 <= not w16699 and not w16700;
w16702 <= not w16698 and not w16701;
w16703 <= not w16698 and not w16702;
w16704 <= not w16701 and not w16702;
w16705 <= not w16703 and not w16704;
w16706 <= w3392 and w12496;
w16707 <= w3477 and w12502;
w16708 <= w3541 and w12499;
w16709 <= not w16707 and not w16708;
w16710 <= not w16706 and w16709;
w16711 <= w3303 and not w15840;
w16712 <= w16710 and not w16711;
w16713 <= a(29) and not w16712;
w16714 <= not w16712 and not w16713;
w16715 <= a(29) and not w16713;
w16716 <= not w16714 and not w16715;
w16717 <= not w16040 and not w16044;
w16718 <= not w16043 and not w16044;
w16719 <= not w16717 and not w16718;
w16720 <= not w16716 and not w16719;
w16721 <= not w16716 and not w16720;
w16722 <= not w16719 and not w16720;
w16723 <= not w16721 and not w16722;
w16724 <= w3392 and w12499;
w16725 <= w3477 and w12506;
w16726 <= w3541 and w12502;
w16727 <= not w16725 and not w16726;
w16728 <= not w16724 and w16727;
w16729 <= w3303 and not w15879;
w16730 <= w16728 and not w16729;
w16731 <= a(29) and not w16730;
w16732 <= not w16730 and not w16731;
w16733 <= a(29) and not w16731;
w16734 <= not w16732 and not w16733;
w16735 <= not w16036 and not w16039;
w16736 <= w16038 and not w16039;
w16737 <= not w16735 and not w16736;
w16738 <= not w16734 and not w16737;
w16739 <= not w16734 and not w16738;
w16740 <= not w16737 and not w16738;
w16741 <= not w16739 and not w16740;
w16742 <= w3392 and w12502;
w16743 <= w3477 and w12509;
w16744 <= w3541 and w12506;
w16745 <= not w16743 and not w16744;
w16746 <= not w16742 and w16745;
w16747 <= w3303 and w15924;
w16748 <= w16746 and not w16747;
w16749 <= a(29) and not w16748;
w16750 <= not w16748 and not w16749;
w16751 <= a(29) and not w16749;
w16752 <= not w16750 and not w16751;
w16753 <= not w16016 and not w16025;
w16754 <= not w16024 and not w16025;
w16755 <= not w16753 and not w16754;
w16756 <= not w16752 and not w16755;
w16757 <= not w16752 and not w16756;
w16758 <= not w16755 and not w16756;
w16759 <= not w16757 and not w16758;
w16760 <= not w7414 and not w12516;
w16761 <= w3541 and not w12516;
w16762 <= w3392 and w12512;
w16763 <= not w16761 and not w16762;
w16764 <= w3303 and not w16020;
w16765 <= w16763 and not w16764;
w16766 <= a(29) and not w16765;
w16767 <= a(29) and not w16766;
w16768 <= not w16765 and not w16766;
w16769 <= not w16767 and not w16768;
w16770 <= not w3302 and not w12516;
w16771 <= a(29) and not w16770;
w16772 <= not w16769 and w16771;
w16773 <= w3392 and w12509;
w16774 <= w3477 and not w12516;
w16775 <= w3541 and w12512;
w16776 <= not w16774 and not w16775;
w16777 <= not w16773 and w16776;
w16778 <= not w3303 and w16777;
w16779 <= w16029 and w16777;
w16780 <= not w16778 and not w16779;
w16781 <= a(29) and not w16780;
w16782 <= not a(29) and w16780;
w16783 <= not w16781 and not w16782;
w16784 <= w16772 and not w16783;
w16785 <= w16760 and w16784;
w16786 <= w3392 and w12506;
w16787 <= w3477 and w12512;
w16788 <= w3541 and w12509;
w16789 <= not w16787 and not w16788;
w16790 <= not w16786 and w16789;
w16791 <= w3303 and w15948;
w16792 <= w16790 and not w16791;
w16793 <= a(29) and not w16792;
w16794 <= not w16792 and not w16793;
w16795 <= a(29) and not w16793;
w16796 <= not w16794 and not w16795;
w16797 <= not w16760 and w16784;
w16798 <= w16760 and not w16784;
w16799 <= not w16797 and not w16798;
w16800 <= not w16796 and not w16799;
w16801 <= not w16785 and not w16800;
w16802 <= not w16759 and not w16801;
w16803 <= not w16756 and not w16802;
w16804 <= not w16741 and not w16803;
w16805 <= not w16738 and not w16804;
w16806 <= not w16723 and not w16805;
w16807 <= not w16720 and not w16806;
w16808 <= not w16705 and not w16807;
w16809 <= not w16702 and not w16808;
w16810 <= not w16687 and not w16809;
w16811 <= not w16684 and not w16810;
w16812 <= w16657 and w16668;
w16813 <= not w16669 and not w16812;
w16814 <= not w16811 and w16813;
w16815 <= not w16669 and not w16814;
w16816 <= w16642 and w16653;
w16817 <= not w16654 and not w16816;
w16818 <= not w16815 and w16817;
w16819 <= not w16654 and not w16818;
w16820 <= w16627 and w16638;
w16821 <= not w16639 and not w16820;
w16822 <= not w16819 and w16821;
w16823 <= not w16639 and not w16822;
w16824 <= w16612 and w16623;
w16825 <= not w16624 and not w16824;
w16826 <= not w16823 and w16825;
w16827 <= not w16624 and not w16826;
w16828 <= w16597 and w16608;
w16829 <= not w16609 and not w16828;
w16830 <= not w16827 and w16829;
w16831 <= not w16609 and not w16830;
w16832 <= not w16083 and w16094;
w16833 <= not w16095 and not w16832;
w16834 <= not w16831 and w16833;
w16835 <= w16831 and not w16833;
w16836 <= not w16834 and not w16835;
w16837 <= w3819 and w12463;
w16838 <= w3902 and w12469;
w16839 <= w3981 and w12466;
w16840 <= not w16838 and not w16839;
w16841 <= not w16837 and w16840;
w16842 <= w3985 and not w14938;
w16843 <= w16841 and not w16842;
w16844 <= a(26) and not w16843;
w16845 <= a(26) and not w16844;
w16846 <= not w16843 and not w16844;
w16847 <= not w16845 and not w16846;
w16848 <= w16836 and not w16847;
w16849 <= not w16834 and not w16848;
w16850 <= not w16594 and not w16849;
w16851 <= w16594 and w16849;
w16852 <= not w16850 and not w16851;
w16853 <= w4629 and w12451;
w16854 <= w4468 and w12457;
w16855 <= w4539 and w12454;
w16856 <= not w16854 and not w16855;
w16857 <= not w16853 and w16856;
w16858 <= w4471 and not w14378;
w16859 <= w16857 and not w16858;
w16860 <= a(23) and not w16859;
w16861 <= a(23) and not w16860;
w16862 <= not w16859 and not w16860;
w16863 <= not w16861 and not w16862;
w16864 <= w16852 and not w16863;
w16865 <= not w16850 and not w16864;
w16866 <= not w16591 and not w16865;
w16867 <= w16591 and w16865;
w16868 <= not w16866 and not w16867;
w16869 <= w5431 and w12440;
w16870 <= w4870 and w12448;
w16871 <= w5342 and w12443;
w16872 <= not w16870 and not w16871;
w16873 <= not w16869 and w16872;
w16874 <= w4873 and not w13986;
w16875 <= w16873 and not w16874;
w16876 <= a(20) and not w16875;
w16877 <= a(20) and not w16876;
w16878 <= not w16875 and not w16876;
w16879 <= not w16877 and not w16878;
w16880 <= w16868 and not w16879;
w16881 <= not w16866 and not w16880;
w16882 <= not w16588 and not w16881;
w16883 <= not w16585 and not w16882;
w16884 <= not w16571 and not w16883;
w16885 <= w16571 and w16883;
w16886 <= not w16884 and not w16885;
w16887 <= w6168 and w13426;
w16888 <= w5598 and w12704;
w16889 <= w5874 and w12824;
w16890 <= not w16888 and not w16889;
w16891 <= not w16887 and w16890;
w16892 <= w5601 and not w13438;
w16893 <= w16891 and not w16892;
w16894 <= a(17) and not w16893;
w16895 <= a(17) and not w16894;
w16896 <= not w16893 and not w16894;
w16897 <= not w16895 and not w16896;
w16898 <= w16886 and not w16897;
w16899 <= not w16884 and not w16898;
w16900 <= not w16568 and not w16899;
w16901 <= w16568 and w16899;
w16902 <= not w16900 and not w16901;
w16903 <= w7036 and w13532;
w16904 <= w6337 and w13456;
w16905 <= w6886 and w13450;
w16906 <= not w16904 and not w16905;
w16907 <= not w16903 and w16906;
w16908 <= w6332 and not w13547;
w16909 <= w16907 and not w16908;
w16910 <= a(14) and not w16909;
w16911 <= a(14) and not w16910;
w16912 <= not w16909 and not w16910;
w16913 <= not w16911 and not w16912;
w16914 <= w16902 and not w16913;
w16915 <= not w16900 and not w16914;
w16916 <= not w16565 and not w16915;
w16917 <= not w16562 and not w16916;
w16918 <= not w16548 and not w16917;
w16919 <= w16548 and w16917;
w16920 <= not w16918 and not w16919;
w16921 <= w7918 and not w13373;
w16922 <= w7226 and not w13562;
w16923 <= w7567 and w13876;
w16924 <= not w16922 and not w16923;
w16925 <= not w16921 and w16924;
w16926 <= w7229 and w13963;
w16927 <= w16925 and not w16926;
w16928 <= a(11) and not w16927;
w16929 <= a(11) and not w16928;
w16930 <= not w16927 and not w16928;
w16931 <= not w16929 and not w16930;
w16932 <= w16920 and not w16931;
w16933 <= not w16918 and not w16932;
w16934 <= not w16545 and not w16933;
w16935 <= w16545 and w16933;
w16936 <= not w16934 and not w16935;
w16937 <= w16920 and not w16932;
w16938 <= not w16931 and not w16932;
w16939 <= not w16937 and not w16938;
w16940 <= w16902 and not w16914;
w16941 <= not w16913 and not w16914;
w16942 <= not w16940 and not w16941;
w16943 <= w16886 and not w16898;
w16944 <= not w16897 and not w16898;
w16945 <= not w16943 and not w16944;
w16946 <= w16588 and w16881;
w16947 <= not w16882 and not w16946;
w16948 <= w6168 and w12824;
w16949 <= w5598 and w12437;
w16950 <= w5874 and w12704;
w16951 <= not w16949 and not w16950;
w16952 <= not w16948 and w16951;
w16953 <= w5601 and w12830;
w16954 <= w16952 and not w16953;
w16955 <= a(17) and not w16954;
w16956 <= a(17) and not w16955;
w16957 <= not w16954 and not w16955;
w16958 <= not w16956 and not w16957;
w16959 <= w16947 and not w16958;
w16960 <= w16947 and not w16959;
w16961 <= not w16958 and not w16959;
w16962 <= not w16960 and not w16961;
w16963 <= w16868 and not w16880;
w16964 <= not w16879 and not w16880;
w16965 <= not w16963 and not w16964;
w16966 <= w16852 and not w16864;
w16967 <= not w16863 and not w16864;
w16968 <= not w16966 and not w16967;
w16969 <= w16836 and not w16848;
w16970 <= not w16847 and not w16848;
w16971 <= not w16969 and not w16970;
w16972 <= w16827 and not w16829;
w16973 <= not w16830 and not w16972;
w16974 <= w3819 and w12466;
w16975 <= w3902 and w12472;
w16976 <= w3981 and w12469;
w16977 <= not w16975 and not w16976;
w16978 <= not w16974 and w16977;
w16979 <= not w3985 and w16978;
w16980 <= not w15190 and w16978;
w16981 <= not w16979 and not w16980;
w16982 <= a(26) and not w16981;
w16983 <= not a(26) and w16981;
w16984 <= not w16982 and not w16983;
w16985 <= w16973 and not w16984;
w16986 <= w16823 and not w16825;
w16987 <= not w16826 and not w16986;
w16988 <= w3819 and w12469;
w16989 <= w3902 and w12475;
w16990 <= w3981 and w12472;
w16991 <= not w16989 and not w16990;
w16992 <= not w16988 and w16991;
w16993 <= not w3985 and w16992;
w16994 <= w15031 and w16992;
w16995 <= not w16993 and not w16994;
w16996 <= a(26) and not w16995;
w16997 <= not a(26) and w16995;
w16998 <= not w16996 and not w16997;
w16999 <= w16987 and not w16998;
w17000 <= w16819 and not w16821;
w17001 <= not w16822 and not w17000;
w17002 <= w3819 and w12472;
w17003 <= w3902 and w12478;
w17004 <= w3981 and w12475;
w17005 <= not w17003 and not w17004;
w17006 <= not w17002 and w17005;
w17007 <= not w3985 and w17006;
w17008 <= w15320 and w17006;
w17009 <= not w17007 and not w17008;
w17010 <= a(26) and not w17009;
w17011 <= not a(26) and w17009;
w17012 <= not w17010 and not w17011;
w17013 <= w17001 and not w17012;
w17014 <= w16815 and not w16817;
w17015 <= not w16818 and not w17014;
w17016 <= w3819 and w12475;
w17017 <= w3902 and w12481;
w17018 <= w3981 and w12478;
w17019 <= not w17017 and not w17018;
w17020 <= not w17016 and w17019;
w17021 <= not w3985 and w17020;
w17022 <= w15643 and w17020;
w17023 <= not w17021 and not w17022;
w17024 <= a(26) and not w17023;
w17025 <= not a(26) and w17023;
w17026 <= not w17024 and not w17025;
w17027 <= w17015 and not w17026;
w17028 <= w16811 and not w16813;
w17029 <= not w16814 and not w17028;
w17030 <= w3819 and w12478;
w17031 <= w3902 and w12484;
w17032 <= w3981 and w12481;
w17033 <= not w17031 and not w17032;
w17034 <= not w17030 and w17033;
w17035 <= not w3985 and w17034;
w17036 <= not w15659 and w17034;
w17037 <= not w17035 and not w17036;
w17038 <= a(26) and not w17037;
w17039 <= not a(26) and w17037;
w17040 <= not w17038 and not w17039;
w17041 <= w17029 and not w17040;
w17042 <= w16687 and w16809;
w17043 <= not w16810 and not w17042;
w17044 <= w3819 and w12481;
w17045 <= w3902 and w12487;
w17046 <= w3981 and w12484;
w17047 <= not w17045 and not w17046;
w17048 <= not w17044 and w17047;
w17049 <= not w3985 and w17048;
w17050 <= w15291 and w17048;
w17051 <= not w17049 and not w17050;
w17052 <= a(26) and not w17051;
w17053 <= not a(26) and w17051;
w17054 <= not w17052 and not w17053;
w17055 <= w17043 and not w17054;
w17056 <= w16705 and w16807;
w17057 <= not w16808 and not w17056;
w17058 <= w3902 and w12490;
w17059 <= w3981 and w12487;
w17060 <= w3819 and w12484;
w17061 <= not w17059 and not w17060;
w17062 <= not w17058 and w17061;
w17063 <= not w3985 and w17062;
w17064 <= not w15699 and w17062;
w17065 <= not w17063 and not w17064;
w17066 <= a(26) and not w17065;
w17067 <= not a(26) and w17065;
w17068 <= not w17066 and not w17067;
w17069 <= w17057 and not w17068;
w17070 <= w16723 and w16805;
w17071 <= not w16806 and not w17070;
w17072 <= w3902 and w12493;
w17073 <= w3819 and w12487;
w17074 <= w3981 and w12490;
w17075 <= not w17073 and not w17074;
w17076 <= not w17072 and w17075;
w17077 <= not w3985 and w17076;
w17078 <= w15726 and w17076;
w17079 <= not w17077 and not w17078;
w17080 <= a(26) and not w17079;
w17081 <= not a(26) and w17079;
w17082 <= not w17080 and not w17081;
w17083 <= w17071 and not w17082;
w17084 <= w16741 and w16803;
w17085 <= not w16804 and not w17084;
w17086 <= w3981 and w12493;
w17087 <= w3819 and w12490;
w17088 <= w3902 and w12496;
w17089 <= not w17087 and not w17088;
w17090 <= not w17086 and w17089;
w17091 <= not w3985 and w17090;
w17092 <= w15751 and w17090;
w17093 <= not w17091 and not w17092;
w17094 <= a(26) and not w17093;
w17095 <= not a(26) and w17093;
w17096 <= not w17094 and not w17095;
w17097 <= w17085 and not w17096;
w17098 <= not w16759 and not w16802;
w17099 <= not w16801 and not w16802;
w17100 <= not w17098 and not w17099;
w17101 <= w3902 and w12499;
w17102 <= w3981 and w12496;
w17103 <= w3819 and w12493;
w17104 <= not w17102 and not w17103;
w17105 <= not w17101 and w17104;
w17106 <= not w3985 and w17105;
w17107 <= not w15782 and w17105;
w17108 <= not w17106 and not w17107;
w17109 <= a(26) and not w17108;
w17110 <= not a(26) and w17108;
w17111 <= not w17109 and not w17110;
w17112 <= not w17100 and not w17111;
w17113 <= w3981 and w12499;
w17114 <= w3819 and w12496;
w17115 <= w3902 and w12502;
w17116 <= not w17114 and not w17115;
w17117 <= not w17113 and w17116;
w17118 <= w3985 and not w15840;
w17119 <= w17117 and not w17118;
w17120 <= a(26) and not w17119;
w17121 <= not w17119 and not w17120;
w17122 <= a(26) and not w17120;
w17123 <= not w17121 and not w17122;
w17124 <= w16796 and w16799;
w17125 <= not w16800 and not w17124;
w17126 <= not w17123 and w17125;
w17127 <= not w17123 and not w17126;
w17128 <= w17125 and not w17126;
w17129 <= not w17127 and not w17128;
w17130 <= w3902 and w12506;
w17131 <= w3981 and w12502;
w17132 <= w3819 and w12499;
w17133 <= not w17131 and not w17132;
w17134 <= not w17130 and w17133;
w17135 <= w3985 and not w15879;
w17136 <= w17134 and not w17135;
w17137 <= a(26) and not w17136;
w17138 <= not w17136 and not w17137;
w17139 <= a(26) and not w17137;
w17140 <= not w17138 and not w17139;
w17141 <= not w16772 and w16783;
w17142 <= not w16784 and not w17141;
w17143 <= not w17140 and w17142;
w17144 <= not w17140 and not w17143;
w17145 <= w17142 and not w17143;
w17146 <= not w17144 and not w17145;
w17147 <= w16769 and not w16771;
w17148 <= not w16772 and not w17147;
w17149 <= w3902 and w12509;
w17150 <= w3819 and w12502;
w17151 <= w3981 and w12506;
w17152 <= not w17150 and not w17151;
w17153 <= not w17149 and w17152;
w17154 <= not w3985 and w17153;
w17155 <= not w15924 and w17153;
w17156 <= not w17154 and not w17155;
w17157 <= a(26) and not w17156;
w17158 <= not a(26) and w17156;
w17159 <= not w17157 and not w17158;
w17160 <= w17148 and not w17159;
w17161 <= w3819 and w12512;
w17162 <= w3981 and not w12516;
w17163 <= not w17161 and not w17162;
w17164 <= w3985 and not w16020;
w17165 <= w17163 and not w17164;
w17166 <= a(26) and not w17165;
w17167 <= a(26) and not w17166;
w17168 <= not w17165 and not w17166;
w17169 <= not w17167 and not w17168;
w17170 <= not w3815 and not w12516;
w17171 <= a(26) and not w17170;
w17172 <= not w17169 and w17171;
w17173 <= w3902 and not w12516;
w17174 <= w3819 and w12509;
w17175 <= w3981 and w12512;
w17176 <= not w17174 and not w17175;
w17177 <= not w17173 and w17176;
w17178 <= not w3985 and w17177;
w17179 <= w16029 and w17177;
w17180 <= not w17178 and not w17179;
w17181 <= a(26) and not w17180;
w17182 <= not a(26) and w17180;
w17183 <= not w17181 and not w17182;
w17184 <= w17172 and not w17183;
w17185 <= w16770 and w17184;
w17186 <= w17184 and not w17185;
w17187 <= w16770 and not w17185;
w17188 <= not w17186 and not w17187;
w17189 <= w3902 and w12512;
w17190 <= w3819 and w12506;
w17191 <= w3981 and w12509;
w17192 <= not w17190 and not w17191;
w17193 <= not w17189 and w17192;
w17194 <= w3985 and w15948;
w17195 <= w17193 and not w17194;
w17196 <= a(26) and not w17195;
w17197 <= a(26) and not w17196;
w17198 <= not w17195 and not w17196;
w17199 <= not w17197 and not w17198;
w17200 <= not w17188 and not w17199;
w17201 <= not w17185 and not w17200;
w17202 <= not w17148 and w17159;
w17203 <= not w17160 and not w17202;
w17204 <= not w17201 and w17203;
w17205 <= not w17160 and not w17204;
w17206 <= not w17146 and not w17205;
w17207 <= not w17143 and not w17206;
w17208 <= not w17129 and not w17207;
w17209 <= not w17126 and not w17208;
w17210 <= not w17100 and not w17112;
w17211 <= not w17111 and not w17112;
w17212 <= not w17210 and not w17211;
w17213 <= not w17209 and not w17212;
w17214 <= not w17112 and not w17213;
w17215 <= w17085 and not w17097;
w17216 <= not w17096 and not w17097;
w17217 <= not w17215 and not w17216;
w17218 <= not w17214 and not w17217;
w17219 <= not w17097 and not w17218;
w17220 <= w17071 and not w17083;
w17221 <= not w17082 and not w17083;
w17222 <= not w17220 and not w17221;
w17223 <= not w17219 and not w17222;
w17224 <= not w17083 and not w17223;
w17225 <= w17057 and not w17069;
w17226 <= not w17068 and not w17069;
w17227 <= not w17225 and not w17226;
w17228 <= not w17224 and not w17227;
w17229 <= not w17069 and not w17228;
w17230 <= w17043 and not w17055;
w17231 <= not w17054 and not w17055;
w17232 <= not w17230 and not w17231;
w17233 <= not w17229 and not w17232;
w17234 <= not w17055 and not w17233;
w17235 <= w17029 and not w17041;
w17236 <= not w17040 and not w17041;
w17237 <= not w17235 and not w17236;
w17238 <= not w17234 and not w17237;
w17239 <= not w17041 and not w17238;
w17240 <= w17015 and not w17027;
w17241 <= not w17026 and not w17027;
w17242 <= not w17240 and not w17241;
w17243 <= not w17239 and not w17242;
w17244 <= not w17027 and not w17243;
w17245 <= w17001 and not w17013;
w17246 <= not w17012 and not w17013;
w17247 <= not w17245 and not w17246;
w17248 <= not w17244 and not w17247;
w17249 <= not w17013 and not w17248;
w17250 <= w16987 and not w16999;
w17251 <= not w16998 and not w16999;
w17252 <= not w17250 and not w17251;
w17253 <= not w17249 and not w17252;
w17254 <= not w16999 and not w17253;
w17255 <= not w16973 and w16984;
w17256 <= not w16985 and not w17255;
w17257 <= not w17254 and w17256;
w17258 <= not w16985 and not w17257;
w17259 <= not w16971 and not w17258;
w17260 <= w16971 and w17258;
w17261 <= not w17259 and not w17260;
w17262 <= w4629 and w12454;
w17263 <= w4468 and w12460;
w17264 <= w4539 and w12457;
w17265 <= not w17263 and not w17264;
w17266 <= not w17262 and w17265;
w17267 <= w4471 and w14389;
w17268 <= w17266 and not w17267;
w17269 <= a(23) and not w17268;
w17270 <= a(23) and not w17269;
w17271 <= not w17268 and not w17269;
w17272 <= not w17270 and not w17271;
w17273 <= w17261 and not w17272;
w17274 <= not w17259 and not w17273;
w17275 <= not w16968 and not w17274;
w17276 <= w16968 and w17274;
w17277 <= not w17275 and not w17276;
w17278 <= w5431 and w12443;
w17279 <= w4870 and w12446;
w17280 <= w5342 and w12448;
w17281 <= not w17279 and not w17280;
w17282 <= not w17278 and w17281;
w17283 <= w4873 and w13798;
w17284 <= w17282 and not w17283;
w17285 <= a(20) and not w17284;
w17286 <= a(20) and not w17285;
w17287 <= not w17284 and not w17285;
w17288 <= not w17286 and not w17287;
w17289 <= w17277 and not w17288;
w17290 <= not w17275 and not w17289;
w17291 <= not w16965 and not w17290;
w17292 <= w16965 and w17290;
w17293 <= not w17291 and not w17292;
w17294 <= w6168 and w12704;
w17295 <= w5598 and w12305;
w17296 <= w5874 and w12437;
w17297 <= not w17295 and not w17296;
w17298 <= not w17294 and w17297;
w17299 <= w5601 and w12934;
w17300 <= w17298 and not w17299;
w17301 <= a(17) and not w17300;
w17302 <= a(17) and not w17301;
w17303 <= not w17300 and not w17301;
w17304 <= not w17302 and not w17303;
w17305 <= w17293 and not w17304;
w17306 <= not w17291 and not w17305;
w17307 <= not w16962 and not w17306;
w17308 <= not w16959 and not w17307;
w17309 <= not w16945 and not w17308;
w17310 <= w16945 and w17308;
w17311 <= not w17309 and not w17310;
w17312 <= w7036 and w13450;
w17313 <= w6337 and w13453;
w17314 <= w6886 and w13456;
w17315 <= not w17313 and not w17314;
w17316 <= not w17312 and w17315;
w17317 <= w6332 and w13476;
w17318 <= w17316 and not w17317;
w17319 <= a(14) and not w17318;
w17320 <= a(14) and not w17319;
w17321 <= not w17318 and not w17319;
w17322 <= not w17320 and not w17321;
w17323 <= w17311 and not w17322;
w17324 <= not w17309 and not w17323;
w17325 <= not w16942 and not w17324;
w17326 <= w16942 and w17324;
w17327 <= not w17325 and not w17326;
w17328 <= w7918 and not w13562;
w17329 <= w7226 and w13565;
w17330 <= w7567 and w13568;
w17331 <= not w17329 and not w17330;
w17332 <= not w17328 and w17331;
w17333 <= w7229 and not w13589;
w17334 <= w17332 and not w17333;
w17335 <= a(11) and not w17334;
w17336 <= a(11) and not w17335;
w17337 <= not w17334 and not w17335;
w17338 <= not w17336 and not w17337;
w17339 <= w17327 and not w17338;
w17340 <= not w17325 and not w17339;
w17341 <= w7918 and w13876;
w17342 <= w7226 and w13568;
w17343 <= w7567 and not w13562;
w17344 <= not w17342 and not w17343;
w17345 <= not w17341 and w17344;
w17346 <= w7229 and w14071;
w17347 <= w17345 and not w17346;
w17348 <= a(11) and not w17347;
w17349 <= a(11) and not w17348;
w17350 <= not w17347 and not w17348;
w17351 <= not w17349 and not w17350;
w17352 <= not w17340 and not w17351;
w17353 <= w16565 and w16915;
w17354 <= not w16916 and not w17353;
w17355 <= not w17340 and not w17352;
w17356 <= not w17351 and not w17352;
w17357 <= not w17355 and not w17356;
w17358 <= w17354 and not w17357;
w17359 <= not w17352 and not w17358;
w17360 <= not w16939 and not w17359;
w17361 <= not w16939 and not w17360;
w17362 <= not w17359 and not w17360;
w17363 <= not w17361 and not w17362;
w17364 <= w17311 and not w17323;
w17365 <= not w17322 and not w17323;
w17366 <= not w17364 and not w17365;
w17367 <= w16962 and w17306;
w17368 <= not w17307 and not w17367;
w17369 <= w7036 and w13456;
w17370 <= w6337 and w13426;
w17371 <= w6886 and w13453;
w17372 <= not w17370 and not w17371;
w17373 <= not w17369 and w17372;
w17374 <= w6332 and not w13844;
w17375 <= w17373 and not w17374;
w17376 <= a(14) and not w17375;
w17377 <= a(14) and not w17376;
w17378 <= not w17375 and not w17376;
w17379 <= not w17377 and not w17378;
w17380 <= w17368 and not w17379;
w17381 <= w17368 and not w17380;
w17382 <= not w17379 and not w17380;
w17383 <= not w17381 and not w17382;
w17384 <= w17293 and not w17305;
w17385 <= not w17304 and not w17305;
w17386 <= not w17384 and not w17385;
w17387 <= w17277 and not w17289;
w17388 <= not w17288 and not w17289;
w17389 <= not w17387 and not w17388;
w17390 <= w17261 and not w17273;
w17391 <= not w17272 and not w17273;
w17392 <= not w17390 and not w17391;
w17393 <= w4629 and w12457;
w17394 <= w4468 and w12463;
w17395 <= w4539 and w12460;
w17396 <= not w17394 and not w17395;
w17397 <= not w17393 and w17396;
w17398 <= w4471 and w14772;
w17399 <= w17397 and not w17398;
w17400 <= a(23) and not w17399;
w17401 <= not w17399 and not w17400;
w17402 <= a(23) and not w17400;
w17403 <= not w17401 and not w17402;
w17404 <= w17254 and not w17256;
w17405 <= not w17257 and not w17404;
w17406 <= not w17403 and w17405;
w17407 <= not w17403 and not w17406;
w17408 <= w17405 and not w17406;
w17409 <= not w17407 and not w17408;
w17410 <= w4629 and w12460;
w17411 <= w4468 and w12466;
w17412 <= w4539 and w12463;
w17413 <= not w17411 and not w17412;
w17414 <= not w17410 and w17413;
w17415 <= w4471 and w14543;
w17416 <= w17414 and not w17415;
w17417 <= a(23) and not w17416;
w17418 <= not w17416 and not w17417;
w17419 <= a(23) and not w17417;
w17420 <= not w17418 and not w17419;
w17421 <= not w17249 and not w17253;
w17422 <= not w17252 and not w17253;
w17423 <= not w17421 and not w17422;
w17424 <= not w17420 and not w17423;
w17425 <= not w17420 and not w17424;
w17426 <= not w17423 and not w17424;
w17427 <= not w17425 and not w17426;
w17428 <= w4629 and w12463;
w17429 <= w4468 and w12469;
w17430 <= w4539 and w12466;
w17431 <= not w17429 and not w17430;
w17432 <= not w17428 and w17431;
w17433 <= w4471 and not w14938;
w17434 <= w17432 and not w17433;
w17435 <= a(23) and not w17434;
w17436 <= not w17434 and not w17435;
w17437 <= a(23) and not w17435;
w17438 <= not w17436 and not w17437;
w17439 <= not w17244 and not w17248;
w17440 <= not w17247 and not w17248;
w17441 <= not w17439 and not w17440;
w17442 <= not w17438 and not w17441;
w17443 <= not w17438 and not w17442;
w17444 <= not w17441 and not w17442;
w17445 <= not w17443 and not w17444;
w17446 <= w4629 and w12466;
w17447 <= w4468 and w12472;
w17448 <= w4539 and w12469;
w17449 <= not w17447 and not w17448;
w17450 <= not w17446 and w17449;
w17451 <= w4471 and w15190;
w17452 <= w17450 and not w17451;
w17453 <= a(23) and not w17452;
w17454 <= not w17452 and not w17453;
w17455 <= a(23) and not w17453;
w17456 <= not w17454 and not w17455;
w17457 <= not w17239 and not w17243;
w17458 <= not w17242 and not w17243;
w17459 <= not w17457 and not w17458;
w17460 <= not w17456 and not w17459;
w17461 <= not w17456 and not w17460;
w17462 <= not w17459 and not w17460;
w17463 <= not w17461 and not w17462;
w17464 <= w4629 and w12469;
w17465 <= w4468 and w12475;
w17466 <= w4539 and w12472;
w17467 <= not w17465 and not w17466;
w17468 <= not w17464 and w17467;
w17469 <= w4471 and not w15031;
w17470 <= w17468 and not w17469;
w17471 <= a(23) and not w17470;
w17472 <= not w17470 and not w17471;
w17473 <= a(23) and not w17471;
w17474 <= not w17472 and not w17473;
w17475 <= not w17234 and not w17238;
w17476 <= not w17237 and not w17238;
w17477 <= not w17475 and not w17476;
w17478 <= not w17474 and not w17477;
w17479 <= not w17474 and not w17478;
w17480 <= not w17477 and not w17478;
w17481 <= not w17479 and not w17480;
w17482 <= w4629 and w12472;
w17483 <= w4468 and w12478;
w17484 <= w4539 and w12475;
w17485 <= not w17483 and not w17484;
w17486 <= not w17482 and w17485;
w17487 <= w4471 and not w15320;
w17488 <= w17486 and not w17487;
w17489 <= a(23) and not w17488;
w17490 <= not w17488 and not w17489;
w17491 <= a(23) and not w17489;
w17492 <= not w17490 and not w17491;
w17493 <= not w17229 and not w17233;
w17494 <= not w17232 and not w17233;
w17495 <= not w17493 and not w17494;
w17496 <= not w17492 and not w17495;
w17497 <= not w17492 and not w17496;
w17498 <= not w17495 and not w17496;
w17499 <= not w17497 and not w17498;
w17500 <= w4629 and w12475;
w17501 <= w4468 and w12481;
w17502 <= w4539 and w12478;
w17503 <= not w17501 and not w17502;
w17504 <= not w17500 and w17503;
w17505 <= w4471 and not w15643;
w17506 <= w17504 and not w17505;
w17507 <= a(23) and not w17506;
w17508 <= not w17506 and not w17507;
w17509 <= a(23) and not w17507;
w17510 <= not w17508 and not w17509;
w17511 <= not w17224 and not w17228;
w17512 <= not w17227 and not w17228;
w17513 <= not w17511 and not w17512;
w17514 <= not w17510 and not w17513;
w17515 <= not w17510 and not w17514;
w17516 <= not w17513 and not w17514;
w17517 <= not w17515 and not w17516;
w17518 <= w4629 and w12478;
w17519 <= w4468 and w12484;
w17520 <= w4539 and w12481;
w17521 <= not w17519 and not w17520;
w17522 <= not w17518 and w17521;
w17523 <= w4471 and w15659;
w17524 <= w17522 and not w17523;
w17525 <= a(23) and not w17524;
w17526 <= not w17524 and not w17525;
w17527 <= a(23) and not w17525;
w17528 <= not w17526 and not w17527;
w17529 <= not w17219 and not w17223;
w17530 <= not w17222 and not w17223;
w17531 <= not w17529 and not w17530;
w17532 <= not w17528 and not w17531;
w17533 <= not w17528 and not w17532;
w17534 <= not w17531 and not w17532;
w17535 <= not w17533 and not w17534;
w17536 <= w4629 and w12481;
w17537 <= w4468 and w12487;
w17538 <= w4539 and w12484;
w17539 <= not w17537 and not w17538;
w17540 <= not w17536 and w17539;
w17541 <= w4471 and not w15291;
w17542 <= w17540 and not w17541;
w17543 <= a(23) and not w17542;
w17544 <= not w17542 and not w17543;
w17545 <= a(23) and not w17543;
w17546 <= not w17544 and not w17545;
w17547 <= not w17214 and not w17218;
w17548 <= not w17217 and not w17218;
w17549 <= not w17547 and not w17548;
w17550 <= not w17546 and not w17549;
w17551 <= not w17546 and not w17550;
w17552 <= not w17549 and not w17550;
w17553 <= not w17551 and not w17552;
w17554 <= w4629 and w12484;
w17555 <= w4468 and w12490;
w17556 <= w4539 and w12487;
w17557 <= not w17555 and not w17556;
w17558 <= not w17554 and w17557;
w17559 <= w4471 and w15699;
w17560 <= w17558 and not w17559;
w17561 <= a(23) and not w17560;
w17562 <= not w17560 and not w17561;
w17563 <= a(23) and not w17561;
w17564 <= not w17562 and not w17563;
w17565 <= not w17209 and not w17213;
w17566 <= not w17212 and not w17213;
w17567 <= not w17565 and not w17566;
w17568 <= not w17564 and not w17567;
w17569 <= not w17564 and not w17568;
w17570 <= not w17567 and not w17568;
w17571 <= not w17569 and not w17570;
w17572 <= w17129 and w17207;
w17573 <= not w17208 and not w17572;
w17574 <= w4629 and w12487;
w17575 <= w4468 and w12493;
w17576 <= w4539 and w12490;
w17577 <= not w17575 and not w17576;
w17578 <= not w17574 and w17577;
w17579 <= not w4471 and w17578;
w17580 <= w15726 and w17578;
w17581 <= not w17579 and not w17580;
w17582 <= a(23) and not w17581;
w17583 <= not a(23) and w17581;
w17584 <= not w17582 and not w17583;
w17585 <= w17573 and not w17584;
w17586 <= w17146 and w17205;
w17587 <= not w17206 and not w17586;
w17588 <= w4629 and w12490;
w17589 <= w4468 and w12496;
w17590 <= w4539 and w12493;
w17591 <= not w17589 and not w17590;
w17592 <= not w17588 and w17591;
w17593 <= not w4471 and w17592;
w17594 <= w15751 and w17592;
w17595 <= not w17593 and not w17594;
w17596 <= a(23) and not w17595;
w17597 <= not a(23) and w17595;
w17598 <= not w17596 and not w17597;
w17599 <= w17587 and not w17598;
w17600 <= w4629 and w12493;
w17601 <= w4468 and w12499;
w17602 <= w4539 and w12496;
w17603 <= not w17601 and not w17602;
w17604 <= not w17600 and w17603;
w17605 <= w4471 and w15782;
w17606 <= w17604 and not w17605;
w17607 <= a(23) and not w17606;
w17608 <= not w17606 and not w17607;
w17609 <= a(23) and not w17607;
w17610 <= not w17608 and not w17609;
w17611 <= w17201 and not w17203;
w17612 <= not w17204 and not w17611;
w17613 <= not w17610 and w17612;
w17614 <= not w17610 and not w17613;
w17615 <= w17612 and not w17613;
w17616 <= not w17614 and not w17615;
w17617 <= not w17188 and not w17200;
w17618 <= not w17199 and not w17200;
w17619 <= not w17617 and not w17618;
w17620 <= w4629 and w12496;
w17621 <= w4468 and w12502;
w17622 <= w4539 and w12499;
w17623 <= not w17621 and not w17622;
w17624 <= not w17620 and w17623;
w17625 <= not w4471 and w17624;
w17626 <= w15840 and w17624;
w17627 <= not w17625 and not w17626;
w17628 <= a(23) and not w17627;
w17629 <= not a(23) and w17627;
w17630 <= not w17628 and not w17629;
w17631 <= not w17619 and not w17630;
w17632 <= w4629 and w12499;
w17633 <= w4468 and w12506;
w17634 <= w4539 and w12502;
w17635 <= not w17633 and not w17634;
w17636 <= not w17632 and w17635;
w17637 <= w4471 and not w15879;
w17638 <= w17636 and not w17637;
w17639 <= a(23) and not w17638;
w17640 <= not w17638 and not w17639;
w17641 <= a(23) and not w17639;
w17642 <= not w17640 and not w17641;
w17643 <= not w17172 and w17183;
w17644 <= not w17184 and not w17643;
w17645 <= not w17642 and w17644;
w17646 <= not w17642 and not w17645;
w17647 <= w17644 and not w17645;
w17648 <= not w17646 and not w17647;
w17649 <= w17169 and not w17171;
w17650 <= not w17172 and not w17649;
w17651 <= w4629 and w12502;
w17652 <= w4468 and w12509;
w17653 <= w4539 and w12506;
w17654 <= not w17652 and not w17653;
w17655 <= not w17651 and w17654;
w17656 <= not w4471 and w17655;
w17657 <= not w15924 and w17655;
w17658 <= not w17656 and not w17657;
w17659 <= a(23) and not w17658;
w17660 <= not a(23) and w17658;
w17661 <= not w17659 and not w17660;
w17662 <= w17650 and not w17661;
w17663 <= w4539 and not w12516;
w17664 <= w4629 and w12512;
w17665 <= not w17663 and not w17664;
w17666 <= w4471 and not w16020;
w17667 <= w17665 and not w17666;
w17668 <= a(23) and not w17667;
w17669 <= a(23) and not w17668;
w17670 <= not w17667 and not w17668;
w17671 <= not w17669 and not w17670;
w17672 <= not w4463 and not w12516;
w17673 <= a(23) and not w17672;
w17674 <= not w17671 and w17673;
w17675 <= w4629 and w12509;
w17676 <= w4468 and not w12516;
w17677 <= w4539 and w12512;
w17678 <= not w17676 and not w17677;
w17679 <= not w17675 and w17678;
w17680 <= not w4471 and w17679;
w17681 <= w16029 and w17679;
w17682 <= not w17680 and not w17681;
w17683 <= a(23) and not w17682;
w17684 <= not a(23) and w17682;
w17685 <= not w17683 and not w17684;
w17686 <= w17674 and not w17685;
w17687 <= w17170 and w17686;
w17688 <= w17686 and not w17687;
w17689 <= w17170 and not w17687;
w17690 <= not w17688 and not w17689;
w17691 <= w4629 and w12506;
w17692 <= w4468 and w12512;
w17693 <= w4539 and w12509;
w17694 <= not w17692 and not w17693;
w17695 <= not w17691 and w17694;
w17696 <= w4471 and w15948;
w17697 <= w17695 and not w17696;
w17698 <= a(23) and not w17697;
w17699 <= a(23) and not w17698;
w17700 <= not w17697 and not w17698;
w17701 <= not w17699 and not w17700;
w17702 <= not w17690 and not w17701;
w17703 <= not w17687 and not w17702;
w17704 <= not w17650 and w17661;
w17705 <= not w17662 and not w17704;
w17706 <= not w17703 and w17705;
w17707 <= not w17662 and not w17706;
w17708 <= not w17648 and not w17707;
w17709 <= not w17645 and not w17708;
w17710 <= w17619 and w17630;
w17711 <= not w17631 and not w17710;
w17712 <= not w17709 and w17711;
w17713 <= not w17631 and not w17712;
w17714 <= not w17616 and not w17713;
w17715 <= not w17613 and not w17714;
w17716 <= w17587 and not w17599;
w17717 <= not w17598 and not w17599;
w17718 <= not w17716 and not w17717;
w17719 <= not w17715 and not w17718;
w17720 <= not w17599 and not w17719;
w17721 <= not w17573 and w17584;
w17722 <= not w17585 and not w17721;
w17723 <= not w17720 and w17722;
w17724 <= not w17585 and not w17723;
w17725 <= not w17571 and not w17724;
w17726 <= not w17568 and not w17725;
w17727 <= not w17553 and not w17726;
w17728 <= not w17550 and not w17727;
w17729 <= not w17535 and not w17728;
w17730 <= not w17532 and not w17729;
w17731 <= not w17517 and not w17730;
w17732 <= not w17514 and not w17731;
w17733 <= not w17499 and not w17732;
w17734 <= not w17496 and not w17733;
w17735 <= not w17481 and not w17734;
w17736 <= not w17478 and not w17735;
w17737 <= not w17463 and not w17736;
w17738 <= not w17460 and not w17737;
w17739 <= not w17445 and not w17738;
w17740 <= not w17442 and not w17739;
w17741 <= not w17427 and not w17740;
w17742 <= not w17424 and not w17741;
w17743 <= not w17409 and not w17742;
w17744 <= not w17406 and not w17743;
w17745 <= not w17392 and not w17744;
w17746 <= w17392 and w17744;
w17747 <= not w17745 and not w17746;
w17748 <= w5431 and w12448;
w17749 <= w4870 and w12451;
w17750 <= w5342 and w12446;
w17751 <= not w17749 and not w17750;
w17752 <= not w17748 and w17751;
w17753 <= w4873 and w14112;
w17754 <= w17752 and not w17753;
w17755 <= a(20) and not w17754;
w17756 <= a(20) and not w17755;
w17757 <= not w17754 and not w17755;
w17758 <= not w17756 and not w17757;
w17759 <= w17747 and not w17758;
w17760 <= not w17745 and not w17759;
w17761 <= not w17389 and not w17760;
w17762 <= w17389 and w17760;
w17763 <= not w17761 and not w17762;
w17764 <= w6168 and w12437;
w17765 <= w5598 and w12440;
w17766 <= w5874 and w12305;
w17767 <= not w17765 and not w17766;
w17768 <= not w17764 and w17767;
w17769 <= w5601 and not w13671;
w17770 <= w17768 and not w17769;
w17771 <= a(17) and not w17770;
w17772 <= a(17) and not w17771;
w17773 <= not w17770 and not w17771;
w17774 <= not w17772 and not w17773;
w17775 <= w17763 and not w17774;
w17776 <= not w17761 and not w17775;
w17777 <= not w17386 and not w17776;
w17778 <= w17386 and w17776;
w17779 <= not w17777 and not w17778;
w17780 <= w7036 and w13453;
w17781 <= w6337 and w12824;
w17782 <= w6886 and w13426;
w17783 <= not w17781 and not w17782;
w17784 <= not w17780 and w17783;
w17785 <= w6332 and w13519;
w17786 <= w17784 and not w17785;
w17787 <= a(14) and not w17786;
w17788 <= a(14) and not w17787;
w17789 <= not w17786 and not w17787;
w17790 <= not w17788 and not w17789;
w17791 <= w17779 and not w17790;
w17792 <= not w17777 and not w17791;
w17793 <= not w17383 and not w17792;
w17794 <= not w17380 and not w17793;
w17795 <= not w17366 and not w17794;
w17796 <= w17366 and w17794;
w17797 <= not w17795 and not w17796;
w17798 <= w7918 and w13568;
w17799 <= w7226 and w13532;
w17800 <= w7567 and w13565;
w17801 <= not w17799 and not w17800;
w17802 <= not w17798 and w17801;
w17803 <= w7229 and w13864;
w17804 <= w17802 and not w17803;
w17805 <= a(11) and not w17804;
w17806 <= a(11) and not w17805;
w17807 <= not w17804 and not w17805;
w17808 <= not w17806 and not w17807;
w17809 <= w17797 and not w17808;
w17810 <= not w17795 and not w17809;
w17811 <= not w13373 and not w14525;
w17812 <= w8353 and w13876;
w17813 <= not w17811 and not w17812;
w17814 <= not w8356 and w17813;
w17815 <= w13886 and w17813;
w17816 <= not w17814 and not w17815;
w17817 <= a(8) and not w17816;
w17818 <= not a(8) and w17816;
w17819 <= not w17817 and not w17818;
w17820 <= not w17810 and not w17819;
w17821 <= w17327 and not w17339;
w17822 <= not w17338 and not w17339;
w17823 <= not w17821 and not w17822;
w17824 <= w17810 and w17819;
w17825 <= not w17820 and not w17824;
w17826 <= not w17823 and w17825;
w17827 <= not w17820 and not w17826;
w17828 <= not w17354 and w17357;
w17829 <= not w17358 and not w17828;
w17830 <= not w17827 and w17829;
w17831 <= not w17823 and not w17826;
w17832 <= w17825 and not w17826;
w17833 <= not w17831 and not w17832;
w17834 <= w17797 and not w17809;
w17835 <= not w17808 and not w17809;
w17836 <= not w17834 and not w17835;
w17837 <= w17383 and w17792;
w17838 <= not w17793 and not w17837;
w17839 <= w7918 and w13565;
w17840 <= w7226 and w13450;
w17841 <= w7567 and w13532;
w17842 <= not w17840 and not w17841;
w17843 <= not w17839 and w17842;
w17844 <= w7229 and w13911;
w17845 <= w17843 and not w17844;
w17846 <= a(11) and not w17845;
w17847 <= a(11) and not w17846;
w17848 <= not w17845 and not w17846;
w17849 <= not w17847 and not w17848;
w17850 <= w17838 and not w17849;
w17851 <= w17838 and not w17850;
w17852 <= not w17849 and not w17850;
w17853 <= not w17851 and not w17852;
w17854 <= w17779 and not w17791;
w17855 <= not w17790 and not w17791;
w17856 <= not w17854 and not w17855;
w17857 <= w17763 and not w17775;
w17858 <= not w17774 and not w17775;
w17859 <= not w17857 and not w17858;
w17860 <= w17747 and not w17759;
w17861 <= not w17758 and not w17759;
w17862 <= not w17860 and not w17861;
w17863 <= w17409 and w17742;
w17864 <= not w17743 and not w17863;
w17865 <= w5431 and w12446;
w17866 <= w4870 and w12454;
w17867 <= w5342 and w12451;
w17868 <= not w17866 and not w17867;
w17869 <= not w17865 and w17868;
w17870 <= not w4873 and w17869;
w17871 <= w14168 and w17869;
w17872 <= not w17870 and not w17871;
w17873 <= a(20) and not w17872;
w17874 <= not a(20) and w17872;
w17875 <= not w17873 and not w17874;
w17876 <= w17864 and not w17875;
w17877 <= w17427 and w17740;
w17878 <= not w17741 and not w17877;
w17879 <= w5431 and w12451;
w17880 <= w4870 and w12457;
w17881 <= w5342 and w12454;
w17882 <= not w17880 and not w17881;
w17883 <= not w17879 and w17882;
w17884 <= not w4873 and w17883;
w17885 <= w14378 and w17883;
w17886 <= not w17884 and not w17885;
w17887 <= a(20) and not w17886;
w17888 <= not a(20) and w17886;
w17889 <= not w17887 and not w17888;
w17890 <= w17878 and not w17889;
w17891 <= w17445 and w17738;
w17892 <= not w17739 and not w17891;
w17893 <= w5431 and w12454;
w17894 <= w4870 and w12460;
w17895 <= w5342 and w12457;
w17896 <= not w17894 and not w17895;
w17897 <= not w17893 and w17896;
w17898 <= not w4873 and w17897;
w17899 <= not w14389 and w17897;
w17900 <= not w17898 and not w17899;
w17901 <= a(20) and not w17900;
w17902 <= not a(20) and w17900;
w17903 <= not w17901 and not w17902;
w17904 <= w17892 and not w17903;
w17905 <= w17463 and w17736;
w17906 <= not w17737 and not w17905;
w17907 <= w5431 and w12457;
w17908 <= w4870 and w12463;
w17909 <= w5342 and w12460;
w17910 <= not w17908 and not w17909;
w17911 <= not w17907 and w17910;
w17912 <= not w4873 and w17911;
w17913 <= not w14772 and w17911;
w17914 <= not w17912 and not w17913;
w17915 <= a(20) and not w17914;
w17916 <= not a(20) and w17914;
w17917 <= not w17915 and not w17916;
w17918 <= w17906 and not w17917;
w17919 <= w17481 and w17734;
w17920 <= not w17735 and not w17919;
w17921 <= w5431 and w12460;
w17922 <= w4870 and w12466;
w17923 <= w5342 and w12463;
w17924 <= not w17922 and not w17923;
w17925 <= not w17921 and w17924;
w17926 <= not w4873 and w17925;
w17927 <= not w14543 and w17925;
w17928 <= not w17926 and not w17927;
w17929 <= a(20) and not w17928;
w17930 <= not a(20) and w17928;
w17931 <= not w17929 and not w17930;
w17932 <= w17920 and not w17931;
w17933 <= w17499 and w17732;
w17934 <= not w17733 and not w17933;
w17935 <= w5431 and w12463;
w17936 <= w4870 and w12469;
w17937 <= w5342 and w12466;
w17938 <= not w17936 and not w17937;
w17939 <= not w17935 and w17938;
w17940 <= not w4873 and w17939;
w17941 <= w14938 and w17939;
w17942 <= not w17940 and not w17941;
w17943 <= a(20) and not w17942;
w17944 <= not a(20) and w17942;
w17945 <= not w17943 and not w17944;
w17946 <= w17934 and not w17945;
w17947 <= w17517 and w17730;
w17948 <= not w17731 and not w17947;
w17949 <= w5431 and w12466;
w17950 <= w4870 and w12472;
w17951 <= w5342 and w12469;
w17952 <= not w17950 and not w17951;
w17953 <= not w17949 and w17952;
w17954 <= not w4873 and w17953;
w17955 <= not w15190 and w17953;
w17956 <= not w17954 and not w17955;
w17957 <= a(20) and not w17956;
w17958 <= not a(20) and w17956;
w17959 <= not w17957 and not w17958;
w17960 <= w17948 and not w17959;
w17961 <= w17535 and w17728;
w17962 <= not w17729 and not w17961;
w17963 <= w5431 and w12469;
w17964 <= w4870 and w12475;
w17965 <= w5342 and w12472;
w17966 <= not w17964 and not w17965;
w17967 <= not w17963 and w17966;
w17968 <= not w4873 and w17967;
w17969 <= w15031 and w17967;
w17970 <= not w17968 and not w17969;
w17971 <= a(20) and not w17970;
w17972 <= not a(20) and w17970;
w17973 <= not w17971 and not w17972;
w17974 <= w17962 and not w17973;
w17975 <= w17553 and w17726;
w17976 <= not w17727 and not w17975;
w17977 <= w5431 and w12472;
w17978 <= w4870 and w12478;
w17979 <= w5342 and w12475;
w17980 <= not w17978 and not w17979;
w17981 <= not w17977 and w17980;
w17982 <= not w4873 and w17981;
w17983 <= w15320 and w17981;
w17984 <= not w17982 and not w17983;
w17985 <= a(20) and not w17984;
w17986 <= not a(20) and w17984;
w17987 <= not w17985 and not w17986;
w17988 <= w17976 and not w17987;
w17989 <= w17571 and w17724;
w17990 <= not w17725 and not w17989;
w17991 <= w5431 and w12475;
w17992 <= w4870 and w12481;
w17993 <= w5342 and w12478;
w17994 <= not w17992 and not w17993;
w17995 <= not w17991 and w17994;
w17996 <= not w4873 and w17995;
w17997 <= w15643 and w17995;
w17998 <= not w17996 and not w17997;
w17999 <= a(20) and not w17998;
w18000 <= not a(20) and w17998;
w18001 <= not w17999 and not w18000;
w18002 <= w17990 and not w18001;
w18003 <= w5431 and w12478;
w18004 <= w4870 and w12484;
w18005 <= w5342 and w12481;
w18006 <= not w18004 and not w18005;
w18007 <= not w18003 and w18006;
w18008 <= w4873 and w15659;
w18009 <= w18007 and not w18008;
w18010 <= a(20) and not w18009;
w18011 <= not w18009 and not w18010;
w18012 <= a(20) and not w18010;
w18013 <= not w18011 and not w18012;
w18014 <= w17720 and not w17722;
w18015 <= not w17723 and not w18014;
w18016 <= not w18013 and w18015;
w18017 <= not w18013 and not w18016;
w18018 <= w18015 and not w18016;
w18019 <= not w18017 and not w18018;
w18020 <= w5431 and w12481;
w18021 <= w4870 and w12487;
w18022 <= w5342 and w12484;
w18023 <= not w18021 and not w18022;
w18024 <= not w18020 and w18023;
w18025 <= w4873 and not w15291;
w18026 <= w18024 and not w18025;
w18027 <= a(20) and not w18026;
w18028 <= not w18026 and not w18027;
w18029 <= a(20) and not w18027;
w18030 <= not w18028 and not w18029;
w18031 <= not w17715 and not w17719;
w18032 <= not w17718 and not w17719;
w18033 <= not w18031 and not w18032;
w18034 <= not w18030 and not w18033;
w18035 <= not w18030 and not w18034;
w18036 <= not w18033 and not w18034;
w18037 <= not w18035 and not w18036;
w18038 <= w17616 and w17713;
w18039 <= not w17714 and not w18038;
w18040 <= w5431 and w12484;
w18041 <= w4870 and w12490;
w18042 <= w5342 and w12487;
w18043 <= not w18041 and not w18042;
w18044 <= not w18040 and w18043;
w18045 <= not w4873 and w18044;
w18046 <= not w15699 and w18044;
w18047 <= not w18045 and not w18046;
w18048 <= a(20) and not w18047;
w18049 <= not a(20) and w18047;
w18050 <= not w18048 and not w18049;
w18051 <= w18039 and not w18050;
w18052 <= w17709 and not w17711;
w18053 <= not w17712 and not w18052;
w18054 <= w5431 and w12487;
w18055 <= w4870 and w12493;
w18056 <= w5342 and w12490;
w18057 <= not w18055 and not w18056;
w18058 <= not w18054 and w18057;
w18059 <= not w4873 and w18058;
w18060 <= w15726 and w18058;
w18061 <= not w18059 and not w18060;
w18062 <= a(20) and not w18061;
w18063 <= not a(20) and w18061;
w18064 <= not w18062 and not w18063;
w18065 <= w18053 and not w18064;
w18066 <= w17648 and w17707;
w18067 <= not w17708 and not w18066;
w18068 <= w5431 and w12490;
w18069 <= w4870 and w12496;
w18070 <= w5342 and w12493;
w18071 <= not w18069 and not w18070;
w18072 <= not w18068 and w18071;
w18073 <= not w4873 and w18072;
w18074 <= w15751 and w18072;
w18075 <= not w18073 and not w18074;
w18076 <= a(20) and not w18075;
w18077 <= not a(20) and w18075;
w18078 <= not w18076 and not w18077;
w18079 <= w18067 and not w18078;
w18080 <= w5431 and w12493;
w18081 <= w4870 and w12499;
w18082 <= w5342 and w12496;
w18083 <= not w18081 and not w18082;
w18084 <= not w18080 and w18083;
w18085 <= w4873 and w15782;
w18086 <= w18084 and not w18085;
w18087 <= a(20) and not w18086;
w18088 <= not w18086 and not w18087;
w18089 <= a(20) and not w18087;
w18090 <= not w18088 and not w18089;
w18091 <= w17703 and not w17705;
w18092 <= not w17706 and not w18091;
w18093 <= not w18090 and w18092;
w18094 <= not w18090 and not w18093;
w18095 <= w18092 and not w18093;
w18096 <= not w18094 and not w18095;
w18097 <= not w17690 and not w17702;
w18098 <= not w17701 and not w17702;
w18099 <= not w18097 and not w18098;
w18100 <= w5431 and w12496;
w18101 <= w4870 and w12502;
w18102 <= w5342 and w12499;
w18103 <= not w18101 and not w18102;
w18104 <= not w18100 and w18103;
w18105 <= not w4873 and w18104;
w18106 <= w15840 and w18104;
w18107 <= not w18105 and not w18106;
w18108 <= a(20) and not w18107;
w18109 <= not a(20) and w18107;
w18110 <= not w18108 and not w18109;
w18111 <= not w18099 and not w18110;
w18112 <= w5431 and w12499;
w18113 <= w4870 and w12506;
w18114 <= w5342 and w12502;
w18115 <= not w18113 and not w18114;
w18116 <= not w18112 and w18115;
w18117 <= w4873 and not w15879;
w18118 <= w18116 and not w18117;
w18119 <= a(20) and not w18118;
w18120 <= not w18118 and not w18119;
w18121 <= a(20) and not w18119;
w18122 <= not w18120 and not w18121;
w18123 <= not w17674 and w17685;
w18124 <= not w17686 and not w18123;
w18125 <= not w18122 and w18124;
w18126 <= not w18122 and not w18125;
w18127 <= w18124 and not w18125;
w18128 <= not w18126 and not w18127;
w18129 <= w17671 and not w17673;
w18130 <= not w17674 and not w18129;
w18131 <= w5431 and w12502;
w18132 <= w4870 and w12509;
w18133 <= w5342 and w12506;
w18134 <= not w18132 and not w18133;
w18135 <= not w18131 and w18134;
w18136 <= not w4873 and w18135;
w18137 <= not w15924 and w18135;
w18138 <= not w18136 and not w18137;
w18139 <= a(20) and not w18138;
w18140 <= not a(20) and w18138;
w18141 <= not w18139 and not w18140;
w18142 <= w18130 and not w18141;
w18143 <= w5342 and not w12516;
w18144 <= w5431 and w12512;
w18145 <= not w18143 and not w18144;
w18146 <= w4873 and not w16020;
w18147 <= w18145 and not w18146;
w18148 <= a(20) and not w18147;
w18149 <= a(20) and not w18148;
w18150 <= not w18147 and not w18148;
w18151 <= not w18149 and not w18150;
w18152 <= not w4868 and not w12516;
w18153 <= a(20) and not w18152;
w18154 <= not w18151 and w18153;
w18155 <= w5431 and w12509;
w18156 <= w4870 and not w12516;
w18157 <= w5342 and w12512;
w18158 <= not w18156 and not w18157;
w18159 <= not w18155 and w18158;
w18160 <= not w4873 and w18159;
w18161 <= w16029 and w18159;
w18162 <= not w18160 and not w18161;
w18163 <= a(20) and not w18162;
w18164 <= not a(20) and w18162;
w18165 <= not w18163 and not w18164;
w18166 <= w18154 and not w18165;
w18167 <= w17672 and w18166;
w18168 <= w18166 and not w18167;
w18169 <= w17672 and not w18167;
w18170 <= not w18168 and not w18169;
w18171 <= w5431 and w12506;
w18172 <= w4870 and w12512;
w18173 <= w5342 and w12509;
w18174 <= not w18172 and not w18173;
w18175 <= not w18171 and w18174;
w18176 <= w4873 and w15948;
w18177 <= w18175 and not w18176;
w18178 <= a(20) and not w18177;
w18179 <= a(20) and not w18178;
w18180 <= not w18177 and not w18178;
w18181 <= not w18179 and not w18180;
w18182 <= not w18170 and not w18181;
w18183 <= not w18167 and not w18182;
w18184 <= not w18130 and w18141;
w18185 <= not w18142 and not w18184;
w18186 <= not w18183 and w18185;
w18187 <= not w18142 and not w18186;
w18188 <= not w18128 and not w18187;
w18189 <= not w18125 and not w18188;
w18190 <= w18099 and w18110;
w18191 <= not w18111 and not w18190;
w18192 <= not w18189 and w18191;
w18193 <= not w18111 and not w18192;
w18194 <= not w18096 and not w18193;
w18195 <= not w18093 and not w18194;
w18196 <= w18067 and not w18079;
w18197 <= not w18078 and not w18079;
w18198 <= not w18196 and not w18197;
w18199 <= not w18195 and not w18198;
w18200 <= not w18079 and not w18199;
w18201 <= w18053 and not w18065;
w18202 <= not w18064 and not w18065;
w18203 <= not w18201 and not w18202;
w18204 <= not w18200 and not w18203;
w18205 <= not w18065 and not w18204;
w18206 <= not w18039 and w18050;
w18207 <= not w18051 and not w18206;
w18208 <= not w18205 and w18207;
w18209 <= not w18051 and not w18208;
w18210 <= not w18037 and not w18209;
w18211 <= not w18034 and not w18210;
w18212 <= not w18019 and not w18211;
w18213 <= not w18016 and not w18212;
w18214 <= w17990 and not w18002;
w18215 <= not w18001 and not w18002;
w18216 <= not w18214 and not w18215;
w18217 <= not w18213 and not w18216;
w18218 <= not w18002 and not w18217;
w18219 <= w17976 and not w17988;
w18220 <= not w17987 and not w17988;
w18221 <= not w18219 and not w18220;
w18222 <= not w18218 and not w18221;
w18223 <= not w17988 and not w18222;
w18224 <= w17962 and not w17974;
w18225 <= not w17973 and not w17974;
w18226 <= not w18224 and not w18225;
w18227 <= not w18223 and not w18226;
w18228 <= not w17974 and not w18227;
w18229 <= w17948 and not w17960;
w18230 <= not w17959 and not w17960;
w18231 <= not w18229 and not w18230;
w18232 <= not w18228 and not w18231;
w18233 <= not w17960 and not w18232;
w18234 <= w17934 and not w17946;
w18235 <= not w17945 and not w17946;
w18236 <= not w18234 and not w18235;
w18237 <= not w18233 and not w18236;
w18238 <= not w17946 and not w18237;
w18239 <= w17920 and not w17932;
w18240 <= not w17931 and not w17932;
w18241 <= not w18239 and not w18240;
w18242 <= not w18238 and not w18241;
w18243 <= not w17932 and not w18242;
w18244 <= w17906 and not w17918;
w18245 <= not w17917 and not w17918;
w18246 <= not w18244 and not w18245;
w18247 <= not w18243 and not w18246;
w18248 <= not w17918 and not w18247;
w18249 <= w17892 and not w17904;
w18250 <= not w17903 and not w17904;
w18251 <= not w18249 and not w18250;
w18252 <= not w18248 and not w18251;
w18253 <= not w17904 and not w18252;
w18254 <= w17878 and not w17890;
w18255 <= not w17889 and not w17890;
w18256 <= not w18254 and not w18255;
w18257 <= not w18253 and not w18256;
w18258 <= not w17890 and not w18257;
w18259 <= not w17864 and w17875;
w18260 <= not w17876 and not w18259;
w18261 <= not w18258 and w18260;
w18262 <= not w17876 and not w18261;
w18263 <= not w17862 and not w18262;
w18264 <= w17862 and w18262;
w18265 <= not w18263 and not w18264;
w18266 <= w6168 and w12305;
w18267 <= w5598 and w12443;
w18268 <= w5874 and w12440;
w18269 <= not w18267 and not w18268;
w18270 <= not w18266 and w18269;
w18271 <= w5601 and not w13683;
w18272 <= w18270 and not w18271;
w18273 <= a(17) and not w18272;
w18274 <= a(17) and not w18273;
w18275 <= not w18272 and not w18273;
w18276 <= not w18274 and not w18275;
w18277 <= w18265 and not w18276;
w18278 <= not w18263 and not w18277;
w18279 <= not w17859 and not w18278;
w18280 <= w17859 and w18278;
w18281 <= not w18279 and not w18280;
w18282 <= w7036 and w13426;
w18283 <= w6337 and w12704;
w18284 <= w6886 and w12824;
w18285 <= not w18283 and not w18284;
w18286 <= not w18282 and w18285;
w18287 <= w6332 and not w13438;
w18288 <= w18286 and not w18287;
w18289 <= a(14) and not w18288;
w18290 <= a(14) and not w18289;
w18291 <= not w18288 and not w18289;
w18292 <= not w18290 and not w18291;
w18293 <= w18281 and not w18292;
w18294 <= not w18279 and not w18293;
w18295 <= not w17856 and not w18294;
w18296 <= w17856 and w18294;
w18297 <= not w18295 and not w18296;
w18298 <= w7918 and w13532;
w18299 <= w7226 and w13456;
w18300 <= w7567 and w13450;
w18301 <= not w18299 and not w18300;
w18302 <= not w18298 and w18301;
w18303 <= w7229 and not w13547;
w18304 <= w18302 and not w18303;
w18305 <= a(11) and not w18304;
w18306 <= a(11) and not w18305;
w18307 <= not w18304 and not w18305;
w18308 <= not w18306 and not w18307;
w18309 <= w18297 and not w18308;
w18310 <= not w18295 and not w18309;
w18311 <= not w17853 and not w18310;
w18312 <= not w17850 and not w18311;
w18313 <= not w17836 and not w18312;
w18314 <= w17836 and w18312;
w18315 <= not w18313 and not w18314;
w18316 <= w9266 and not w13373;
w18317 <= w8353 and not w13562;
w18318 <= w8795 and w13876;
w18319 <= not w18317 and not w18318;
w18320 <= not w18316 and w18319;
w18321 <= w8356 and w13963;
w18322 <= w18320 and not w18321;
w18323 <= a(8) and not w18322;
w18324 <= a(8) and not w18323;
w18325 <= not w18322 and not w18323;
w18326 <= not w18324 and not w18325;
w18327 <= w18315 and not w18326;
w18328 <= not w18313 and not w18327;
w18329 <= not w17833 and not w18328;
w18330 <= w17833 and w18328;
w18331 <= not w18329 and not w18330;
w18332 <= w18315 and not w18327;
w18333 <= not w18326 and not w18327;
w18334 <= not w18332 and not w18333;
w18335 <= w18297 and not w18309;
w18336 <= not w18308 and not w18309;
w18337 <= not w18335 and not w18336;
w18338 <= w18281 and not w18293;
w18339 <= not w18292 and not w18293;
w18340 <= not w18338 and not w18339;
w18341 <= w18265 and not w18277;
w18342 <= not w18276 and not w18277;
w18343 <= not w18341 and not w18342;
w18344 <= w6168 and w12440;
w18345 <= w5598 and w12448;
w18346 <= w5874 and w12443;
w18347 <= not w18345 and not w18346;
w18348 <= not w18344 and w18347;
w18349 <= w5601 and not w13986;
w18350 <= w18348 and not w18349;
w18351 <= a(17) and not w18350;
w18352 <= not w18350 and not w18351;
w18353 <= a(17) and not w18351;
w18354 <= not w18352 and not w18353;
w18355 <= w18258 and not w18260;
w18356 <= not w18261 and not w18355;
w18357 <= not w18354 and w18356;
w18358 <= not w18354 and not w18357;
w18359 <= w18356 and not w18357;
w18360 <= not w18358 and not w18359;
w18361 <= w6168 and w12443;
w18362 <= w5598 and w12446;
w18363 <= w5874 and w12448;
w18364 <= not w18362 and not w18363;
w18365 <= not w18361 and w18364;
w18366 <= w5601 and w13798;
w18367 <= w18365 and not w18366;
w18368 <= a(17) and not w18367;
w18369 <= not w18367 and not w18368;
w18370 <= a(17) and not w18368;
w18371 <= not w18369 and not w18370;
w18372 <= not w18253 and not w18257;
w18373 <= not w18256 and not w18257;
w18374 <= not w18372 and not w18373;
w18375 <= not w18371 and not w18374;
w18376 <= not w18371 and not w18375;
w18377 <= not w18374 and not w18375;
w18378 <= not w18376 and not w18377;
w18379 <= w6168 and w12448;
w18380 <= w5598 and w12451;
w18381 <= w5874 and w12446;
w18382 <= not w18380 and not w18381;
w18383 <= not w18379 and w18382;
w18384 <= w5601 and w14112;
w18385 <= w18383 and not w18384;
w18386 <= a(17) and not w18385;
w18387 <= not w18385 and not w18386;
w18388 <= a(17) and not w18386;
w18389 <= not w18387 and not w18388;
w18390 <= not w18248 and not w18252;
w18391 <= not w18251 and not w18252;
w18392 <= not w18390 and not w18391;
w18393 <= not w18389 and not w18392;
w18394 <= not w18389 and not w18393;
w18395 <= not w18392 and not w18393;
w18396 <= not w18394 and not w18395;
w18397 <= w6168 and w12446;
w18398 <= w5598 and w12454;
w18399 <= w5874 and w12451;
w18400 <= not w18398 and not w18399;
w18401 <= not w18397 and w18400;
w18402 <= w5601 and not w14168;
w18403 <= w18401 and not w18402;
w18404 <= a(17) and not w18403;
w18405 <= not w18403 and not w18404;
w18406 <= a(17) and not w18404;
w18407 <= not w18405 and not w18406;
w18408 <= not w18243 and not w18247;
w18409 <= not w18246 and not w18247;
w18410 <= not w18408 and not w18409;
w18411 <= not w18407 and not w18410;
w18412 <= not w18407 and not w18411;
w18413 <= not w18410 and not w18411;
w18414 <= not w18412 and not w18413;
w18415 <= w6168 and w12451;
w18416 <= w5598 and w12457;
w18417 <= w5874 and w12454;
w18418 <= not w18416 and not w18417;
w18419 <= not w18415 and w18418;
w18420 <= w5601 and not w14378;
w18421 <= w18419 and not w18420;
w18422 <= a(17) and not w18421;
w18423 <= not w18421 and not w18422;
w18424 <= a(17) and not w18422;
w18425 <= not w18423 and not w18424;
w18426 <= not w18238 and not w18242;
w18427 <= not w18241 and not w18242;
w18428 <= not w18426 and not w18427;
w18429 <= not w18425 and not w18428;
w18430 <= not w18425 and not w18429;
w18431 <= not w18428 and not w18429;
w18432 <= not w18430 and not w18431;
w18433 <= w6168 and w12454;
w18434 <= w5598 and w12460;
w18435 <= w5874 and w12457;
w18436 <= not w18434 and not w18435;
w18437 <= not w18433 and w18436;
w18438 <= w5601 and w14389;
w18439 <= w18437 and not w18438;
w18440 <= a(17) and not w18439;
w18441 <= not w18439 and not w18440;
w18442 <= a(17) and not w18440;
w18443 <= not w18441 and not w18442;
w18444 <= not w18233 and not w18237;
w18445 <= not w18236 and not w18237;
w18446 <= not w18444 and not w18445;
w18447 <= not w18443 and not w18446;
w18448 <= not w18443 and not w18447;
w18449 <= not w18446 and not w18447;
w18450 <= not w18448 and not w18449;
w18451 <= w6168 and w12457;
w18452 <= w5598 and w12463;
w18453 <= w5874 and w12460;
w18454 <= not w18452 and not w18453;
w18455 <= not w18451 and w18454;
w18456 <= w5601 and w14772;
w18457 <= w18455 and not w18456;
w18458 <= a(17) and not w18457;
w18459 <= not w18457 and not w18458;
w18460 <= a(17) and not w18458;
w18461 <= not w18459 and not w18460;
w18462 <= not w18228 and not w18232;
w18463 <= not w18231 and not w18232;
w18464 <= not w18462 and not w18463;
w18465 <= not w18461 and not w18464;
w18466 <= not w18461 and not w18465;
w18467 <= not w18464 and not w18465;
w18468 <= not w18466 and not w18467;
w18469 <= w6168 and w12460;
w18470 <= w5598 and w12466;
w18471 <= w5874 and w12463;
w18472 <= not w18470 and not w18471;
w18473 <= not w18469 and w18472;
w18474 <= w5601 and w14543;
w18475 <= w18473 and not w18474;
w18476 <= a(17) and not w18475;
w18477 <= not w18475 and not w18476;
w18478 <= a(17) and not w18476;
w18479 <= not w18477 and not w18478;
w18480 <= not w18223 and not w18227;
w18481 <= not w18226 and not w18227;
w18482 <= not w18480 and not w18481;
w18483 <= not w18479 and not w18482;
w18484 <= not w18479 and not w18483;
w18485 <= not w18482 and not w18483;
w18486 <= not w18484 and not w18485;
w18487 <= w6168 and w12463;
w18488 <= w5598 and w12469;
w18489 <= w5874 and w12466;
w18490 <= not w18488 and not w18489;
w18491 <= not w18487 and w18490;
w18492 <= w5601 and not w14938;
w18493 <= w18491 and not w18492;
w18494 <= a(17) and not w18493;
w18495 <= not w18493 and not w18494;
w18496 <= a(17) and not w18494;
w18497 <= not w18495 and not w18496;
w18498 <= not w18218 and not w18222;
w18499 <= not w18221 and not w18222;
w18500 <= not w18498 and not w18499;
w18501 <= not w18497 and not w18500;
w18502 <= not w18497 and not w18501;
w18503 <= not w18500 and not w18501;
w18504 <= not w18502 and not w18503;
w18505 <= w6168 and w12466;
w18506 <= w5598 and w12472;
w18507 <= w5874 and w12469;
w18508 <= not w18506 and not w18507;
w18509 <= not w18505 and w18508;
w18510 <= w5601 and w15190;
w18511 <= w18509 and not w18510;
w18512 <= a(17) and not w18511;
w18513 <= not w18511 and not w18512;
w18514 <= a(17) and not w18512;
w18515 <= not w18513 and not w18514;
w18516 <= not w18213 and not w18217;
w18517 <= not w18216 and not w18217;
w18518 <= not w18516 and not w18517;
w18519 <= not w18515 and not w18518;
w18520 <= not w18515 and not w18519;
w18521 <= not w18518 and not w18519;
w18522 <= not w18520 and not w18521;
w18523 <= w18019 and w18211;
w18524 <= not w18212 and not w18523;
w18525 <= w6168 and w12469;
w18526 <= w5598 and w12475;
w18527 <= w5874 and w12472;
w18528 <= not w18526 and not w18527;
w18529 <= not w18525 and w18528;
w18530 <= not w5601 and w18529;
w18531 <= w15031 and w18529;
w18532 <= not w18530 and not w18531;
w18533 <= a(17) and not w18532;
w18534 <= not a(17) and w18532;
w18535 <= not w18533 and not w18534;
w18536 <= w18524 and not w18535;
w18537 <= w18037 and w18209;
w18538 <= not w18210 and not w18537;
w18539 <= w6168 and w12472;
w18540 <= w5598 and w12478;
w18541 <= w5874 and w12475;
w18542 <= not w18540 and not w18541;
w18543 <= not w18539 and w18542;
w18544 <= not w5601 and w18543;
w18545 <= w15320 and w18543;
w18546 <= not w18544 and not w18545;
w18547 <= a(17) and not w18546;
w18548 <= not a(17) and w18546;
w18549 <= not w18547 and not w18548;
w18550 <= w18538 and not w18549;
w18551 <= w6168 and w12475;
w18552 <= w5598 and w12481;
w18553 <= w5874 and w12478;
w18554 <= not w18552 and not w18553;
w18555 <= not w18551 and w18554;
w18556 <= w5601 and not w15643;
w18557 <= w18555 and not w18556;
w18558 <= a(17) and not w18557;
w18559 <= not w18557 and not w18558;
w18560 <= a(17) and not w18558;
w18561 <= not w18559 and not w18560;
w18562 <= w18205 and not w18207;
w18563 <= not w18208 and not w18562;
w18564 <= not w18561 and w18563;
w18565 <= not w18561 and not w18564;
w18566 <= w18563 and not w18564;
w18567 <= not w18565 and not w18566;
w18568 <= w6168 and w12478;
w18569 <= w5598 and w12484;
w18570 <= w5874 and w12481;
w18571 <= not w18569 and not w18570;
w18572 <= not w18568 and w18571;
w18573 <= w5601 and w15659;
w18574 <= w18572 and not w18573;
w18575 <= a(17) and not w18574;
w18576 <= not w18574 and not w18575;
w18577 <= a(17) and not w18575;
w18578 <= not w18576 and not w18577;
w18579 <= not w18200 and not w18204;
w18580 <= not w18203 and not w18204;
w18581 <= not w18579 and not w18580;
w18582 <= not w18578 and not w18581;
w18583 <= not w18578 and not w18582;
w18584 <= not w18581 and not w18582;
w18585 <= not w18583 and not w18584;
w18586 <= w6168 and w12481;
w18587 <= w5598 and w12487;
w18588 <= w5874 and w12484;
w18589 <= not w18587 and not w18588;
w18590 <= not w18586 and w18589;
w18591 <= w5601 and not w15291;
w18592 <= w18590 and not w18591;
w18593 <= a(17) and not w18592;
w18594 <= not w18592 and not w18593;
w18595 <= a(17) and not w18593;
w18596 <= not w18594 and not w18595;
w18597 <= not w18195 and not w18199;
w18598 <= not w18198 and not w18199;
w18599 <= not w18597 and not w18598;
w18600 <= not w18596 and not w18599;
w18601 <= not w18596 and not w18600;
w18602 <= not w18599 and not w18600;
w18603 <= not w18601 and not w18602;
w18604 <= w18096 and w18193;
w18605 <= not w18194 and not w18604;
w18606 <= w6168 and w12484;
w18607 <= w5598 and w12490;
w18608 <= w5874 and w12487;
w18609 <= not w18607 and not w18608;
w18610 <= not w18606 and w18609;
w18611 <= not w5601 and w18610;
w18612 <= not w15699 and w18610;
w18613 <= not w18611 and not w18612;
w18614 <= a(17) and not w18613;
w18615 <= not a(17) and w18613;
w18616 <= not w18614 and not w18615;
w18617 <= w18605 and not w18616;
w18618 <= w18189 and not w18191;
w18619 <= not w18192 and not w18618;
w18620 <= w6168 and w12487;
w18621 <= w5598 and w12493;
w18622 <= w5874 and w12490;
w18623 <= not w18621 and not w18622;
w18624 <= not w18620 and w18623;
w18625 <= not w5601 and w18624;
w18626 <= w15726 and w18624;
w18627 <= not w18625 and not w18626;
w18628 <= a(17) and not w18627;
w18629 <= not a(17) and w18627;
w18630 <= not w18628 and not w18629;
w18631 <= w18619 and not w18630;
w18632 <= w18128 and w18187;
w18633 <= not w18188 and not w18632;
w18634 <= w6168 and w12490;
w18635 <= w5598 and w12496;
w18636 <= w5874 and w12493;
w18637 <= not w18635 and not w18636;
w18638 <= not w18634 and w18637;
w18639 <= not w5601 and w18638;
w18640 <= w15751 and w18638;
w18641 <= not w18639 and not w18640;
w18642 <= a(17) and not w18641;
w18643 <= not a(17) and w18641;
w18644 <= not w18642 and not w18643;
w18645 <= w18633 and not w18644;
w18646 <= w6168 and w12493;
w18647 <= w5598 and w12499;
w18648 <= w5874 and w12496;
w18649 <= not w18647 and not w18648;
w18650 <= not w18646 and w18649;
w18651 <= w5601 and w15782;
w18652 <= w18650 and not w18651;
w18653 <= a(17) and not w18652;
w18654 <= not w18652 and not w18653;
w18655 <= a(17) and not w18653;
w18656 <= not w18654 and not w18655;
w18657 <= w18183 and not w18185;
w18658 <= not w18186 and not w18657;
w18659 <= not w18656 and w18658;
w18660 <= not w18656 and not w18659;
w18661 <= w18658 and not w18659;
w18662 <= not w18660 and not w18661;
w18663 <= not w18170 and not w18182;
w18664 <= not w18181 and not w18182;
w18665 <= not w18663 and not w18664;
w18666 <= w6168 and w12496;
w18667 <= w5598 and w12502;
w18668 <= w5874 and w12499;
w18669 <= not w18667 and not w18668;
w18670 <= not w18666 and w18669;
w18671 <= not w5601 and w18670;
w18672 <= w15840 and w18670;
w18673 <= not w18671 and not w18672;
w18674 <= a(17) and not w18673;
w18675 <= not a(17) and w18673;
w18676 <= not w18674 and not w18675;
w18677 <= not w18665 and not w18676;
w18678 <= w6168 and w12499;
w18679 <= w5598 and w12506;
w18680 <= w5874 and w12502;
w18681 <= not w18679 and not w18680;
w18682 <= not w18678 and w18681;
w18683 <= w5601 and not w15879;
w18684 <= w18682 and not w18683;
w18685 <= a(17) and not w18684;
w18686 <= not w18684 and not w18685;
w18687 <= a(17) and not w18685;
w18688 <= not w18686 and not w18687;
w18689 <= not w18154 and w18165;
w18690 <= not w18166 and not w18689;
w18691 <= not w18688 and w18690;
w18692 <= not w18688 and not w18691;
w18693 <= w18690 and not w18691;
w18694 <= not w18692 and not w18693;
w18695 <= w18151 and not w18153;
w18696 <= not w18154 and not w18695;
w18697 <= w6168 and w12502;
w18698 <= w5598 and w12509;
w18699 <= w5874 and w12506;
w18700 <= not w18698 and not w18699;
w18701 <= not w18697 and w18700;
w18702 <= not w5601 and w18701;
w18703 <= not w15924 and w18701;
w18704 <= not w18702 and not w18703;
w18705 <= a(17) and not w18704;
w18706 <= not a(17) and w18704;
w18707 <= not w18705 and not w18706;
w18708 <= w18696 and not w18707;
w18709 <= w5874 and not w12516;
w18710 <= w6168 and w12512;
w18711 <= not w18709 and not w18710;
w18712 <= w5601 and not w16020;
w18713 <= w18711 and not w18712;
w18714 <= a(17) and not w18713;
w18715 <= a(17) and not w18714;
w18716 <= not w18713 and not w18714;
w18717 <= not w18715 and not w18716;
w18718 <= not w5593 and not w12516;
w18719 <= a(17) and not w18718;
w18720 <= not w18717 and w18719;
w18721 <= w6168 and w12509;
w18722 <= w5598 and not w12516;
w18723 <= w5874 and w12512;
w18724 <= not w18722 and not w18723;
w18725 <= not w18721 and w18724;
w18726 <= not w5601 and w18725;
w18727 <= w16029 and w18725;
w18728 <= not w18726 and not w18727;
w18729 <= a(17) and not w18728;
w18730 <= not a(17) and w18728;
w18731 <= not w18729 and not w18730;
w18732 <= w18720 and not w18731;
w18733 <= w18152 and w18732;
w18734 <= w18732 and not w18733;
w18735 <= w18152 and not w18733;
w18736 <= not w18734 and not w18735;
w18737 <= w6168 and w12506;
w18738 <= w5598 and w12512;
w18739 <= w5874 and w12509;
w18740 <= not w18738 and not w18739;
w18741 <= not w18737 and w18740;
w18742 <= w5601 and w15948;
w18743 <= w18741 and not w18742;
w18744 <= a(17) and not w18743;
w18745 <= a(17) and not w18744;
w18746 <= not w18743 and not w18744;
w18747 <= not w18745 and not w18746;
w18748 <= not w18736 and not w18747;
w18749 <= not w18733 and not w18748;
w18750 <= not w18696 and w18707;
w18751 <= not w18708 and not w18750;
w18752 <= not w18749 and w18751;
w18753 <= not w18708 and not w18752;
w18754 <= not w18694 and not w18753;
w18755 <= not w18691 and not w18754;
w18756 <= w18665 and w18676;
w18757 <= not w18677 and not w18756;
w18758 <= not w18755 and w18757;
w18759 <= not w18677 and not w18758;
w18760 <= not w18662 and not w18759;
w18761 <= not w18659 and not w18760;
w18762 <= w18633 and not w18645;
w18763 <= not w18644 and not w18645;
w18764 <= not w18762 and not w18763;
w18765 <= not w18761 and not w18764;
w18766 <= not w18645 and not w18765;
w18767 <= w18619 and not w18631;
w18768 <= not w18630 and not w18631;
w18769 <= not w18767 and not w18768;
w18770 <= not w18766 and not w18769;
w18771 <= not w18631 and not w18770;
w18772 <= not w18605 and w18616;
w18773 <= not w18617 and not w18772;
w18774 <= not w18771 and w18773;
w18775 <= not w18617 and not w18774;
w18776 <= not w18603 and not w18775;
w18777 <= not w18600 and not w18776;
w18778 <= not w18585 and not w18777;
w18779 <= not w18582 and not w18778;
w18780 <= not w18567 and not w18779;
w18781 <= not w18564 and not w18780;
w18782 <= w18538 and not w18550;
w18783 <= not w18549 and not w18550;
w18784 <= not w18782 and not w18783;
w18785 <= not w18781 and not w18784;
w18786 <= not w18550 and not w18785;
w18787 <= not w18524 and w18535;
w18788 <= not w18536 and not w18787;
w18789 <= not w18786 and w18788;
w18790 <= not w18536 and not w18789;
w18791 <= not w18522 and not w18790;
w18792 <= not w18519 and not w18791;
w18793 <= not w18504 and not w18792;
w18794 <= not w18501 and not w18793;
w18795 <= not w18486 and not w18794;
w18796 <= not w18483 and not w18795;
w18797 <= not w18468 and not w18796;
w18798 <= not w18465 and not w18797;
w18799 <= not w18450 and not w18798;
w18800 <= not w18447 and not w18799;
w18801 <= not w18432 and not w18800;
w18802 <= not w18429 and not w18801;
w18803 <= not w18414 and not w18802;
w18804 <= not w18411 and not w18803;
w18805 <= not w18396 and not w18804;
w18806 <= not w18393 and not w18805;
w18807 <= not w18378 and not w18806;
w18808 <= not w18375 and not w18807;
w18809 <= not w18360 and not w18808;
w18810 <= not w18357 and not w18809;
w18811 <= not w18343 and not w18810;
w18812 <= w18343 and w18810;
w18813 <= not w18811 and not w18812;
w18814 <= w7036 and w12824;
w18815 <= w6337 and w12437;
w18816 <= w6886 and w12704;
w18817 <= not w18815 and not w18816;
w18818 <= not w18814 and w18817;
w18819 <= w6332 and w12830;
w18820 <= w18818 and not w18819;
w18821 <= a(14) and not w18820;
w18822 <= a(14) and not w18821;
w18823 <= not w18820 and not w18821;
w18824 <= not w18822 and not w18823;
w18825 <= w18813 and not w18824;
w18826 <= not w18811 and not w18825;
w18827 <= not w18340 and not w18826;
w18828 <= w18340 and w18826;
w18829 <= not w18827 and not w18828;
w18830 <= w7918 and w13450;
w18831 <= w7226 and w13453;
w18832 <= w7567 and w13456;
w18833 <= not w18831 and not w18832;
w18834 <= not w18830 and w18833;
w18835 <= w7229 and w13476;
w18836 <= w18834 and not w18835;
w18837 <= a(11) and not w18836;
w18838 <= a(11) and not w18837;
w18839 <= not w18836 and not w18837;
w18840 <= not w18838 and not w18839;
w18841 <= w18829 and not w18840;
w18842 <= not w18827 and not w18841;
w18843 <= not w18337 and not w18842;
w18844 <= w18337 and w18842;
w18845 <= not w18843 and not w18844;
w18846 <= w9266 and not w13562;
w18847 <= w8353 and w13565;
w18848 <= w8795 and w13568;
w18849 <= not w18847 and not w18848;
w18850 <= not w18846 and w18849;
w18851 <= w8356 and not w13589;
w18852 <= w18850 and not w18851;
w18853 <= a(8) and not w18852;
w18854 <= a(8) and not w18853;
w18855 <= not w18852 and not w18853;
w18856 <= not w18854 and not w18855;
w18857 <= w18845 and not w18856;
w18858 <= not w18843 and not w18857;
w18859 <= w9266 and w13876;
w18860 <= w8353 and w13568;
w18861 <= w8795 and not w13562;
w18862 <= not w18860 and not w18861;
w18863 <= not w18859 and w18862;
w18864 <= w8356 and w14071;
w18865 <= w18863 and not w18864;
w18866 <= a(8) and not w18865;
w18867 <= a(8) and not w18866;
w18868 <= not w18865 and not w18866;
w18869 <= not w18867 and not w18868;
w18870 <= not w18858 and not w18869;
w18871 <= not w18858 and not w18870;
w18872 <= not w18869 and not w18870;
w18873 <= not w18871 and not w18872;
w18874 <= w17853 and w18310;
w18875 <= not w18311 and not w18874;
w18876 <= not w18873 and w18875;
w18877 <= not w18870 and not w18876;
w18878 <= not w18334 and not w18877;
w18879 <= not w18334 and not w18878;
w18880 <= not w18877 and not w18878;
w18881 <= not w18879 and not w18880;
w18882 <= w18829 and not w18841;
w18883 <= not w18840 and not w18841;
w18884 <= not w18882 and not w18883;
w18885 <= w18813 and not w18825;
w18886 <= not w18824 and not w18825;
w18887 <= not w18885 and not w18886;
w18888 <= w18360 and w18808;
w18889 <= not w18809 and not w18888;
w18890 <= w7036 and w12704;
w18891 <= w6337 and w12305;
w18892 <= w6886 and w12437;
w18893 <= not w18891 and not w18892;
w18894 <= not w18890 and w18893;
w18895 <= not w6332 and w18894;
w18896 <= not w12934 and w18894;
w18897 <= not w18895 and not w18896;
w18898 <= a(14) and not w18897;
w18899 <= not a(14) and w18897;
w18900 <= not w18898 and not w18899;
w18901 <= w18889 and not w18900;
w18902 <= w18378 and w18806;
w18903 <= not w18807 and not w18902;
w18904 <= w7036 and w12437;
w18905 <= w6337 and w12440;
w18906 <= w6886 and w12305;
w18907 <= not w18905 and not w18906;
w18908 <= not w18904 and w18907;
w18909 <= not w6332 and w18908;
w18910 <= w13671 and w18908;
w18911 <= not w18909 and not w18910;
w18912 <= a(14) and not w18911;
w18913 <= not a(14) and w18911;
w18914 <= not w18912 and not w18913;
w18915 <= w18903 and not w18914;
w18916 <= w18396 and w18804;
w18917 <= not w18805 and not w18916;
w18918 <= w7036 and w12305;
w18919 <= w6337 and w12443;
w18920 <= w6886 and w12440;
w18921 <= not w18919 and not w18920;
w18922 <= not w18918 and w18921;
w18923 <= not w6332 and w18922;
w18924 <= w13683 and w18922;
w18925 <= not w18923 and not w18924;
w18926 <= a(14) and not w18925;
w18927 <= not a(14) and w18925;
w18928 <= not w18926 and not w18927;
w18929 <= w18917 and not w18928;
w18930 <= w18414 and w18802;
w18931 <= not w18803 and not w18930;
w18932 <= w7036 and w12440;
w18933 <= w6337 and w12448;
w18934 <= w6886 and w12443;
w18935 <= not w18933 and not w18934;
w18936 <= not w18932 and w18935;
w18937 <= not w6332 and w18936;
w18938 <= w13986 and w18936;
w18939 <= not w18937 and not w18938;
w18940 <= a(14) and not w18939;
w18941 <= not a(14) and w18939;
w18942 <= not w18940 and not w18941;
w18943 <= w18931 and not w18942;
w18944 <= w18432 and w18800;
w18945 <= not w18801 and not w18944;
w18946 <= w7036 and w12443;
w18947 <= w6337 and w12446;
w18948 <= w6886 and w12448;
w18949 <= not w18947 and not w18948;
w18950 <= not w18946 and w18949;
w18951 <= not w6332 and w18950;
w18952 <= not w13798 and w18950;
w18953 <= not w18951 and not w18952;
w18954 <= a(14) and not w18953;
w18955 <= not a(14) and w18953;
w18956 <= not w18954 and not w18955;
w18957 <= w18945 and not w18956;
w18958 <= w18450 and w18798;
w18959 <= not w18799 and not w18958;
w18960 <= w7036 and w12448;
w18961 <= w6337 and w12451;
w18962 <= w6886 and w12446;
w18963 <= not w18961 and not w18962;
w18964 <= not w18960 and w18963;
w18965 <= not w6332 and w18964;
w18966 <= not w14112 and w18964;
w18967 <= not w18965 and not w18966;
w18968 <= a(14) and not w18967;
w18969 <= not a(14) and w18967;
w18970 <= not w18968 and not w18969;
w18971 <= w18959 and not w18970;
w18972 <= w18468 and w18796;
w18973 <= not w18797 and not w18972;
w18974 <= w7036 and w12446;
w18975 <= w6337 and w12454;
w18976 <= w6886 and w12451;
w18977 <= not w18975 and not w18976;
w18978 <= not w18974 and w18977;
w18979 <= not w6332 and w18978;
w18980 <= w14168 and w18978;
w18981 <= not w18979 and not w18980;
w18982 <= a(14) and not w18981;
w18983 <= not a(14) and w18981;
w18984 <= not w18982 and not w18983;
w18985 <= w18973 and not w18984;
w18986 <= w18486 and w18794;
w18987 <= not w18795 and not w18986;
w18988 <= w7036 and w12451;
w18989 <= w6337 and w12457;
w18990 <= w6886 and w12454;
w18991 <= not w18989 and not w18990;
w18992 <= not w18988 and w18991;
w18993 <= not w6332 and w18992;
w18994 <= w14378 and w18992;
w18995 <= not w18993 and not w18994;
w18996 <= a(14) and not w18995;
w18997 <= not a(14) and w18995;
w18998 <= not w18996 and not w18997;
w18999 <= w18987 and not w18998;
w19000 <= w18504 and w18792;
w19001 <= not w18793 and not w19000;
w19002 <= w7036 and w12454;
w19003 <= w6337 and w12460;
w19004 <= w6886 and w12457;
w19005 <= not w19003 and not w19004;
w19006 <= not w19002 and w19005;
w19007 <= not w6332 and w19006;
w19008 <= not w14389 and w19006;
w19009 <= not w19007 and not w19008;
w19010 <= a(14) and not w19009;
w19011 <= not a(14) and w19009;
w19012 <= not w19010 and not w19011;
w19013 <= w19001 and not w19012;
w19014 <= w18522 and w18790;
w19015 <= not w18791 and not w19014;
w19016 <= w7036 and w12457;
w19017 <= w6337 and w12463;
w19018 <= w6886 and w12460;
w19019 <= not w19017 and not w19018;
w19020 <= not w19016 and w19019;
w19021 <= not w6332 and w19020;
w19022 <= not w14772 and w19020;
w19023 <= not w19021 and not w19022;
w19024 <= a(14) and not w19023;
w19025 <= not a(14) and w19023;
w19026 <= not w19024 and not w19025;
w19027 <= w19015 and not w19026;
w19028 <= w7036 and w12460;
w19029 <= w6337 and w12466;
w19030 <= w6886 and w12463;
w19031 <= not w19029 and not w19030;
w19032 <= not w19028 and w19031;
w19033 <= w6332 and w14543;
w19034 <= w19032 and not w19033;
w19035 <= a(14) and not w19034;
w19036 <= not w19034 and not w19035;
w19037 <= a(14) and not w19035;
w19038 <= not w19036 and not w19037;
w19039 <= w18786 and not w18788;
w19040 <= not w18789 and not w19039;
w19041 <= not w19038 and w19040;
w19042 <= not w19038 and not w19041;
w19043 <= w19040 and not w19041;
w19044 <= not w19042 and not w19043;
w19045 <= w7036 and w12463;
w19046 <= w6337 and w12469;
w19047 <= w6886 and w12466;
w19048 <= not w19046 and not w19047;
w19049 <= not w19045 and w19048;
w19050 <= w6332 and not w14938;
w19051 <= w19049 and not w19050;
w19052 <= a(14) and not w19051;
w19053 <= not w19051 and not w19052;
w19054 <= a(14) and not w19052;
w19055 <= not w19053 and not w19054;
w19056 <= not w18781 and not w18785;
w19057 <= not w18784 and not w18785;
w19058 <= not w19056 and not w19057;
w19059 <= not w19055 and not w19058;
w19060 <= not w19055 and not w19059;
w19061 <= not w19058 and not w19059;
w19062 <= not w19060 and not w19061;
w19063 <= w18567 and w18779;
w19064 <= not w18780 and not w19063;
w19065 <= w7036 and w12466;
w19066 <= w6337 and w12472;
w19067 <= w6886 and w12469;
w19068 <= not w19066 and not w19067;
w19069 <= not w19065 and w19068;
w19070 <= not w6332 and w19069;
w19071 <= not w15190 and w19069;
w19072 <= not w19070 and not w19071;
w19073 <= a(14) and not w19072;
w19074 <= not a(14) and w19072;
w19075 <= not w19073 and not w19074;
w19076 <= w19064 and not w19075;
w19077 <= w18585 and w18777;
w19078 <= not w18778 and not w19077;
w19079 <= w7036 and w12469;
w19080 <= w6337 and w12475;
w19081 <= w6886 and w12472;
w19082 <= not w19080 and not w19081;
w19083 <= not w19079 and w19082;
w19084 <= not w6332 and w19083;
w19085 <= w15031 and w19083;
w19086 <= not w19084 and not w19085;
w19087 <= a(14) and not w19086;
w19088 <= not a(14) and w19086;
w19089 <= not w19087 and not w19088;
w19090 <= w19078 and not w19089;
w19091 <= w18603 and w18775;
w19092 <= not w18776 and not w19091;
w19093 <= w7036 and w12472;
w19094 <= w6337 and w12478;
w19095 <= w6886 and w12475;
w19096 <= not w19094 and not w19095;
w19097 <= not w19093 and w19096;
w19098 <= not w6332 and w19097;
w19099 <= w15320 and w19097;
w19100 <= not w19098 and not w19099;
w19101 <= a(14) and not w19100;
w19102 <= not a(14) and w19100;
w19103 <= not w19101 and not w19102;
w19104 <= w19092 and not w19103;
w19105 <= w7036 and w12475;
w19106 <= w6337 and w12481;
w19107 <= w6886 and w12478;
w19108 <= not w19106 and not w19107;
w19109 <= not w19105 and w19108;
w19110 <= w6332 and not w15643;
w19111 <= w19109 and not w19110;
w19112 <= a(14) and not w19111;
w19113 <= not w19111 and not w19112;
w19114 <= a(14) and not w19112;
w19115 <= not w19113 and not w19114;
w19116 <= w18771 and not w18773;
w19117 <= not w18774 and not w19116;
w19118 <= not w19115 and w19117;
w19119 <= not w19115 and not w19118;
w19120 <= w19117 and not w19118;
w19121 <= not w19119 and not w19120;
w19122 <= w7036 and w12478;
w19123 <= w6337 and w12484;
w19124 <= w6886 and w12481;
w19125 <= not w19123 and not w19124;
w19126 <= not w19122 and w19125;
w19127 <= w6332 and w15659;
w19128 <= w19126 and not w19127;
w19129 <= a(14) and not w19128;
w19130 <= not w19128 and not w19129;
w19131 <= a(14) and not w19129;
w19132 <= not w19130 and not w19131;
w19133 <= not w18766 and not w18770;
w19134 <= not w18769 and not w18770;
w19135 <= not w19133 and not w19134;
w19136 <= not w19132 and not w19135;
w19137 <= not w19132 and not w19136;
w19138 <= not w19135 and not w19136;
w19139 <= not w19137 and not w19138;
w19140 <= w7036 and w12481;
w19141 <= w6337 and w12487;
w19142 <= w6886 and w12484;
w19143 <= not w19141 and not w19142;
w19144 <= not w19140 and w19143;
w19145 <= w6332 and not w15291;
w19146 <= w19144 and not w19145;
w19147 <= a(14) and not w19146;
w19148 <= not w19146 and not w19147;
w19149 <= a(14) and not w19147;
w19150 <= not w19148 and not w19149;
w19151 <= not w18761 and not w18765;
w19152 <= not w18764 and not w18765;
w19153 <= not w19151 and not w19152;
w19154 <= not w19150 and not w19153;
w19155 <= not w19150 and not w19154;
w19156 <= not w19153 and not w19154;
w19157 <= not w19155 and not w19156;
w19158 <= w18662 and w18759;
w19159 <= not w18760 and not w19158;
w19160 <= w7036 and w12484;
w19161 <= w6337 and w12490;
w19162 <= w6886 and w12487;
w19163 <= not w19161 and not w19162;
w19164 <= not w19160 and w19163;
w19165 <= not w6332 and w19164;
w19166 <= not w15699 and w19164;
w19167 <= not w19165 and not w19166;
w19168 <= a(14) and not w19167;
w19169 <= not a(14) and w19167;
w19170 <= not w19168 and not w19169;
w19171 <= w19159 and not w19170;
w19172 <= w18755 and not w18757;
w19173 <= not w18758 and not w19172;
w19174 <= w7036 and w12487;
w19175 <= w6337 and w12493;
w19176 <= w6886 and w12490;
w19177 <= not w19175 and not w19176;
w19178 <= not w19174 and w19177;
w19179 <= not w6332 and w19178;
w19180 <= w15726 and w19178;
w19181 <= not w19179 and not w19180;
w19182 <= a(14) and not w19181;
w19183 <= not a(14) and w19181;
w19184 <= not w19182 and not w19183;
w19185 <= w19173 and not w19184;
w19186 <= w18694 and w18753;
w19187 <= not w18754 and not w19186;
w19188 <= w7036 and w12490;
w19189 <= w6337 and w12496;
w19190 <= w6886 and w12493;
w19191 <= not w19189 and not w19190;
w19192 <= not w19188 and w19191;
w19193 <= not w6332 and w19192;
w19194 <= w15751 and w19192;
w19195 <= not w19193 and not w19194;
w19196 <= a(14) and not w19195;
w19197 <= not a(14) and w19195;
w19198 <= not w19196 and not w19197;
w19199 <= w19187 and not w19198;
w19200 <= w7036 and w12493;
w19201 <= w6337 and w12499;
w19202 <= w6886 and w12496;
w19203 <= not w19201 and not w19202;
w19204 <= not w19200 and w19203;
w19205 <= w6332 and w15782;
w19206 <= w19204 and not w19205;
w19207 <= a(14) and not w19206;
w19208 <= not w19206 and not w19207;
w19209 <= a(14) and not w19207;
w19210 <= not w19208 and not w19209;
w19211 <= w18749 and not w18751;
w19212 <= not w18752 and not w19211;
w19213 <= not w19210 and w19212;
w19214 <= not w19210 and not w19213;
w19215 <= w19212 and not w19213;
w19216 <= not w19214 and not w19215;
w19217 <= not w18736 and not w18748;
w19218 <= not w18747 and not w18748;
w19219 <= not w19217 and not w19218;
w19220 <= w7036 and w12496;
w19221 <= w6337 and w12502;
w19222 <= w6886 and w12499;
w19223 <= not w19221 and not w19222;
w19224 <= not w19220 and w19223;
w19225 <= not w6332 and w19224;
w19226 <= w15840 and w19224;
w19227 <= not w19225 and not w19226;
w19228 <= a(14) and not w19227;
w19229 <= not a(14) and w19227;
w19230 <= not w19228 and not w19229;
w19231 <= not w19219 and not w19230;
w19232 <= w7036 and w12499;
w19233 <= w6337 and w12506;
w19234 <= w6886 and w12502;
w19235 <= not w19233 and not w19234;
w19236 <= not w19232 and w19235;
w19237 <= w6332 and not w15879;
w19238 <= w19236 and not w19237;
w19239 <= a(14) and not w19238;
w19240 <= not w19238 and not w19239;
w19241 <= a(14) and not w19239;
w19242 <= not w19240 and not w19241;
w19243 <= not w18720 and w18731;
w19244 <= not w18732 and not w19243;
w19245 <= not w19242 and w19244;
w19246 <= not w19242 and not w19245;
w19247 <= w19244 and not w19245;
w19248 <= not w19246 and not w19247;
w19249 <= w18717 and not w18719;
w19250 <= not w18720 and not w19249;
w19251 <= w7036 and w12502;
w19252 <= w6337 and w12509;
w19253 <= w6886 and w12506;
w19254 <= not w19252 and not w19253;
w19255 <= not w19251 and w19254;
w19256 <= not w6332 and w19255;
w19257 <= not w15924 and w19255;
w19258 <= not w19256 and not w19257;
w19259 <= a(14) and not w19258;
w19260 <= not a(14) and w19258;
w19261 <= not w19259 and not w19260;
w19262 <= w19250 and not w19261;
w19263 <= w6886 and not w12516;
w19264 <= w7036 and w12512;
w19265 <= not w19263 and not w19264;
w19266 <= w6332 and not w16020;
w19267 <= w19265 and not w19266;
w19268 <= a(14) and not w19267;
w19269 <= a(14) and not w19268;
w19270 <= not w19267 and not w19268;
w19271 <= not w19269 and not w19270;
w19272 <= not w6328 and not w12516;
w19273 <= a(14) and not w19272;
w19274 <= not w19271 and w19273;
w19275 <= w7036 and w12509;
w19276 <= w6337 and not w12516;
w19277 <= w6886 and w12512;
w19278 <= not w19276 and not w19277;
w19279 <= not w19275 and w19278;
w19280 <= not w6332 and w19279;
w19281 <= w16029 and w19279;
w19282 <= not w19280 and not w19281;
w19283 <= a(14) and not w19282;
w19284 <= not a(14) and w19282;
w19285 <= not w19283 and not w19284;
w19286 <= w19274 and not w19285;
w19287 <= w18718 and w19286;
w19288 <= w19286 and not w19287;
w19289 <= w18718 and not w19287;
w19290 <= not w19288 and not w19289;
w19291 <= w7036 and w12506;
w19292 <= w6337 and w12512;
w19293 <= w6886 and w12509;
w19294 <= not w19292 and not w19293;
w19295 <= not w19291 and w19294;
w19296 <= w6332 and w15948;
w19297 <= w19295 and not w19296;
w19298 <= a(14) and not w19297;
w19299 <= a(14) and not w19298;
w19300 <= not w19297 and not w19298;
w19301 <= not w19299 and not w19300;
w19302 <= not w19290 and not w19301;
w19303 <= not w19287 and not w19302;
w19304 <= not w19250 and w19261;
w19305 <= not w19262 and not w19304;
w19306 <= not w19303 and w19305;
w19307 <= not w19262 and not w19306;
w19308 <= not w19248 and not w19307;
w19309 <= not w19245 and not w19308;
w19310 <= w19219 and w19230;
w19311 <= not w19231 and not w19310;
w19312 <= not w19309 and w19311;
w19313 <= not w19231 and not w19312;
w19314 <= not w19216 and not w19313;
w19315 <= not w19213 and not w19314;
w19316 <= w19187 and not w19199;
w19317 <= not w19198 and not w19199;
w19318 <= not w19316 and not w19317;
w19319 <= not w19315 and not w19318;
w19320 <= not w19199 and not w19319;
w19321 <= w19173 and not w19185;
w19322 <= not w19184 and not w19185;
w19323 <= not w19321 and not w19322;
w19324 <= not w19320 and not w19323;
w19325 <= not w19185 and not w19324;
w19326 <= not w19159 and w19170;
w19327 <= not w19171 and not w19326;
w19328 <= not w19325 and w19327;
w19329 <= not w19171 and not w19328;
w19330 <= not w19157 and not w19329;
w19331 <= not w19154 and not w19330;
w19332 <= not w19139 and not w19331;
w19333 <= not w19136 and not w19332;
w19334 <= not w19121 and not w19333;
w19335 <= not w19118 and not w19334;
w19336 <= w19092 and not w19104;
w19337 <= not w19103 and not w19104;
w19338 <= not w19336 and not w19337;
w19339 <= not w19335 and not w19338;
w19340 <= not w19104 and not w19339;
w19341 <= w19078 and not w19090;
w19342 <= not w19089 and not w19090;
w19343 <= not w19341 and not w19342;
w19344 <= not w19340 and not w19343;
w19345 <= not w19090 and not w19344;
w19346 <= not w19064 and w19075;
w19347 <= not w19076 and not w19346;
w19348 <= not w19345 and w19347;
w19349 <= not w19076 and not w19348;
w19350 <= not w19062 and not w19349;
w19351 <= not w19059 and not w19350;
w19352 <= not w19044 and not w19351;
w19353 <= not w19041 and not w19352;
w19354 <= w19015 and not w19027;
w19355 <= not w19026 and not w19027;
w19356 <= not w19354 and not w19355;
w19357 <= not w19353 and not w19356;
w19358 <= not w19027 and not w19357;
w19359 <= w19001 and not w19013;
w19360 <= not w19012 and not w19013;
w19361 <= not w19359 and not w19360;
w19362 <= not w19358 and not w19361;
w19363 <= not w19013 and not w19362;
w19364 <= w18987 and not w18999;
w19365 <= not w18998 and not w18999;
w19366 <= not w19364 and not w19365;
w19367 <= not w19363 and not w19366;
w19368 <= not w18999 and not w19367;
w19369 <= w18973 and not w18985;
w19370 <= not w18984 and not w18985;
w19371 <= not w19369 and not w19370;
w19372 <= not w19368 and not w19371;
w19373 <= not w18985 and not w19372;
w19374 <= w18959 and not w18971;
w19375 <= not w18970 and not w18971;
w19376 <= not w19374 and not w19375;
w19377 <= not w19373 and not w19376;
w19378 <= not w18971 and not w19377;
w19379 <= w18945 and not w18957;
w19380 <= not w18956 and not w18957;
w19381 <= not w19379 and not w19380;
w19382 <= not w19378 and not w19381;
w19383 <= not w18957 and not w19382;
w19384 <= w18931 and not w18943;
w19385 <= not w18942 and not w18943;
w19386 <= not w19384 and not w19385;
w19387 <= not w19383 and not w19386;
w19388 <= not w18943 and not w19387;
w19389 <= w18917 and not w18929;
w19390 <= not w18928 and not w18929;
w19391 <= not w19389 and not w19390;
w19392 <= not w19388 and not w19391;
w19393 <= not w18929 and not w19392;
w19394 <= w18903 and not w18915;
w19395 <= not w18914 and not w18915;
w19396 <= not w19394 and not w19395;
w19397 <= not w19393 and not w19396;
w19398 <= not w18915 and not w19397;
w19399 <= not w18889 and w18900;
w19400 <= not w18901 and not w19399;
w19401 <= not w19398 and w19400;
w19402 <= not w18901 and not w19401;
w19403 <= not w18887 and not w19402;
w19404 <= w18887 and w19402;
w19405 <= not w19403 and not w19404;
w19406 <= w7918 and w13456;
w19407 <= w7226 and w13426;
w19408 <= w7567 and w13453;
w19409 <= not w19407 and not w19408;
w19410 <= not w19406 and w19409;
w19411 <= w7229 and not w13844;
w19412 <= w19410 and not w19411;
w19413 <= a(11) and not w19412;
w19414 <= a(11) and not w19413;
w19415 <= not w19412 and not w19413;
w19416 <= not w19414 and not w19415;
w19417 <= w19405 and not w19416;
w19418 <= not w19403 and not w19417;
w19419 <= not w18884 and not w19418;
w19420 <= w18884 and w19418;
w19421 <= not w19419 and not w19420;
w19422 <= w9266 and w13568;
w19423 <= w8353 and w13532;
w19424 <= w8795 and w13565;
w19425 <= not w19423 and not w19424;
w19426 <= not w19422 and w19425;
w19427 <= w8356 and w13864;
w19428 <= w19426 and not w19427;
w19429 <= a(8) and not w19428;
w19430 <= a(8) and not w19429;
w19431 <= not w19428 and not w19429;
w19432 <= not w19430 and not w19431;
w19433 <= w19421 and not w19432;
w19434 <= not w19419 and not w19433;
w19435 <= not w13373 and not w15011;
w19436 <= w9802 and w13876;
w19437 <= not w19435 and not w19436;
w19438 <= not w9805 and w19437;
w19439 <= w13886 and w19437;
w19440 <= not w19438 and not w19439;
w19441 <= a(5) and not w19440;
w19442 <= not a(5) and w19440;
w19443 <= not w19441 and not w19442;
w19444 <= not w19434 and not w19443;
w19445 <= w18845 and not w18857;
w19446 <= not w18856 and not w18857;
w19447 <= not w19445 and not w19446;
w19448 <= w19434 and w19443;
w19449 <= not w19444 and not w19448;
w19450 <= not w19447 and w19449;
w19451 <= not w19444 and not w19450;
w19452 <= w18873 and not w18875;
w19453 <= not w18876 and not w19452;
w19454 <= not w19451 and w19453;
w19455 <= not w19447 and not w19450;
w19456 <= w19449 and not w19450;
w19457 <= not w19455 and not w19456;
w19458 <= w19421 and not w19433;
w19459 <= not w19432 and not w19433;
w19460 <= not w19458 and not w19459;
w19461 <= w19405 and not w19417;
w19462 <= not w19416 and not w19417;
w19463 <= not w19461 and not w19462;
w19464 <= w7918 and w13453;
w19465 <= w7226 and w12824;
w19466 <= w7567 and w13426;
w19467 <= not w19465 and not w19466;
w19468 <= not w19464 and w19467;
w19469 <= w7229 and w13519;
w19470 <= w19468 and not w19469;
w19471 <= a(11) and not w19470;
w19472 <= not w19470 and not w19471;
w19473 <= a(11) and not w19471;
w19474 <= not w19472 and not w19473;
w19475 <= w19398 and not w19400;
w19476 <= not w19401 and not w19475;
w19477 <= not w19474 and w19476;
w19478 <= not w19474 and not w19477;
w19479 <= w19476 and not w19477;
w19480 <= not w19478 and not w19479;
w19481 <= w7918 and w13426;
w19482 <= w7226 and w12704;
w19483 <= w7567 and w12824;
w19484 <= not w19482 and not w19483;
w19485 <= not w19481 and w19484;
w19486 <= w7229 and not w13438;
w19487 <= w19485 and not w19486;
w19488 <= a(11) and not w19487;
w19489 <= not w19487 and not w19488;
w19490 <= a(11) and not w19488;
w19491 <= not w19489 and not w19490;
w19492 <= not w19393 and not w19397;
w19493 <= not w19396 and not w19397;
w19494 <= not w19492 and not w19493;
w19495 <= not w19491 and not w19494;
w19496 <= not w19491 and not w19495;
w19497 <= not w19494 and not w19495;
w19498 <= not w19496 and not w19497;
w19499 <= w7918 and w12824;
w19500 <= w7226 and w12437;
w19501 <= w7567 and w12704;
w19502 <= not w19500 and not w19501;
w19503 <= not w19499 and w19502;
w19504 <= w7229 and w12830;
w19505 <= w19503 and not w19504;
w19506 <= a(11) and not w19505;
w19507 <= not w19505 and not w19506;
w19508 <= a(11) and not w19506;
w19509 <= not w19507 and not w19508;
w19510 <= not w19388 and not w19392;
w19511 <= not w19391 and not w19392;
w19512 <= not w19510 and not w19511;
w19513 <= not w19509 and not w19512;
w19514 <= not w19509 and not w19513;
w19515 <= not w19512 and not w19513;
w19516 <= not w19514 and not w19515;
w19517 <= w7918 and w12704;
w19518 <= w7226 and w12305;
w19519 <= w7567 and w12437;
w19520 <= not w19518 and not w19519;
w19521 <= not w19517 and w19520;
w19522 <= w7229 and w12934;
w19523 <= w19521 and not w19522;
w19524 <= a(11) and not w19523;
w19525 <= not w19523 and not w19524;
w19526 <= a(11) and not w19524;
w19527 <= not w19525 and not w19526;
w19528 <= not w19383 and not w19387;
w19529 <= not w19386 and not w19387;
w19530 <= not w19528 and not w19529;
w19531 <= not w19527 and not w19530;
w19532 <= not w19527 and not w19531;
w19533 <= not w19530 and not w19531;
w19534 <= not w19532 and not w19533;
w19535 <= w7918 and w12437;
w19536 <= w7226 and w12440;
w19537 <= w7567 and w12305;
w19538 <= not w19536 and not w19537;
w19539 <= not w19535 and w19538;
w19540 <= w7229 and not w13671;
w19541 <= w19539 and not w19540;
w19542 <= a(11) and not w19541;
w19543 <= not w19541 and not w19542;
w19544 <= a(11) and not w19542;
w19545 <= not w19543 and not w19544;
w19546 <= not w19378 and not w19382;
w19547 <= not w19381 and not w19382;
w19548 <= not w19546 and not w19547;
w19549 <= not w19545 and not w19548;
w19550 <= not w19545 and not w19549;
w19551 <= not w19548 and not w19549;
w19552 <= not w19550 and not w19551;
w19553 <= w7918 and w12305;
w19554 <= w7226 and w12443;
w19555 <= w7567 and w12440;
w19556 <= not w19554 and not w19555;
w19557 <= not w19553 and w19556;
w19558 <= w7229 and not w13683;
w19559 <= w19557 and not w19558;
w19560 <= a(11) and not w19559;
w19561 <= not w19559 and not w19560;
w19562 <= a(11) and not w19560;
w19563 <= not w19561 and not w19562;
w19564 <= not w19373 and not w19377;
w19565 <= not w19376 and not w19377;
w19566 <= not w19564 and not w19565;
w19567 <= not w19563 and not w19566;
w19568 <= not w19563 and not w19567;
w19569 <= not w19566 and not w19567;
w19570 <= not w19568 and not w19569;
w19571 <= w7918 and w12440;
w19572 <= w7226 and w12448;
w19573 <= w7567 and w12443;
w19574 <= not w19572 and not w19573;
w19575 <= not w19571 and w19574;
w19576 <= w7229 and not w13986;
w19577 <= w19575 and not w19576;
w19578 <= a(11) and not w19577;
w19579 <= not w19577 and not w19578;
w19580 <= a(11) and not w19578;
w19581 <= not w19579 and not w19580;
w19582 <= not w19368 and not w19372;
w19583 <= not w19371 and not w19372;
w19584 <= not w19582 and not w19583;
w19585 <= not w19581 and not w19584;
w19586 <= not w19581 and not w19585;
w19587 <= not w19584 and not w19585;
w19588 <= not w19586 and not w19587;
w19589 <= w7918 and w12443;
w19590 <= w7226 and w12446;
w19591 <= w7567 and w12448;
w19592 <= not w19590 and not w19591;
w19593 <= not w19589 and w19592;
w19594 <= w7229 and w13798;
w19595 <= w19593 and not w19594;
w19596 <= a(11) and not w19595;
w19597 <= not w19595 and not w19596;
w19598 <= a(11) and not w19596;
w19599 <= not w19597 and not w19598;
w19600 <= not w19363 and not w19367;
w19601 <= not w19366 and not w19367;
w19602 <= not w19600 and not w19601;
w19603 <= not w19599 and not w19602;
w19604 <= not w19599 and not w19603;
w19605 <= not w19602 and not w19603;
w19606 <= not w19604 and not w19605;
w19607 <= w7918 and w12448;
w19608 <= w7226 and w12451;
w19609 <= w7567 and w12446;
w19610 <= not w19608 and not w19609;
w19611 <= not w19607 and w19610;
w19612 <= w7229 and w14112;
w19613 <= w19611 and not w19612;
w19614 <= a(11) and not w19613;
w19615 <= not w19613 and not w19614;
w19616 <= a(11) and not w19614;
w19617 <= not w19615 and not w19616;
w19618 <= not w19358 and not w19362;
w19619 <= not w19361 and not w19362;
w19620 <= not w19618 and not w19619;
w19621 <= not w19617 and not w19620;
w19622 <= not w19617 and not w19621;
w19623 <= not w19620 and not w19621;
w19624 <= not w19622 and not w19623;
w19625 <= w7918 and w12446;
w19626 <= w7226 and w12454;
w19627 <= w7567 and w12451;
w19628 <= not w19626 and not w19627;
w19629 <= not w19625 and w19628;
w19630 <= w7229 and not w14168;
w19631 <= w19629 and not w19630;
w19632 <= a(11) and not w19631;
w19633 <= not w19631 and not w19632;
w19634 <= a(11) and not w19632;
w19635 <= not w19633 and not w19634;
w19636 <= not w19353 and not w19357;
w19637 <= not w19356 and not w19357;
w19638 <= not w19636 and not w19637;
w19639 <= not w19635 and not w19638;
w19640 <= not w19635 and not w19639;
w19641 <= not w19638 and not w19639;
w19642 <= not w19640 and not w19641;
w19643 <= w19044 and w19351;
w19644 <= not w19352 and not w19643;
w19645 <= w7918 and w12451;
w19646 <= w7226 and w12457;
w19647 <= w7567 and w12454;
w19648 <= not w19646 and not w19647;
w19649 <= not w19645 and w19648;
w19650 <= not w7229 and w19649;
w19651 <= w14378 and w19649;
w19652 <= not w19650 and not w19651;
w19653 <= a(11) and not w19652;
w19654 <= not a(11) and w19652;
w19655 <= not w19653 and not w19654;
w19656 <= w19644 and not w19655;
w19657 <= w19062 and w19349;
w19658 <= not w19350 and not w19657;
w19659 <= w7918 and w12454;
w19660 <= w7226 and w12460;
w19661 <= w7567 and w12457;
w19662 <= not w19660 and not w19661;
w19663 <= not w19659 and w19662;
w19664 <= not w7229 and w19663;
w19665 <= not w14389 and w19663;
w19666 <= not w19664 and not w19665;
w19667 <= a(11) and not w19666;
w19668 <= not a(11) and w19666;
w19669 <= not w19667 and not w19668;
w19670 <= w19658 and not w19669;
w19671 <= w7918 and w12457;
w19672 <= w7226 and w12463;
w19673 <= w7567 and w12460;
w19674 <= not w19672 and not w19673;
w19675 <= not w19671 and w19674;
w19676 <= w7229 and w14772;
w19677 <= w19675 and not w19676;
w19678 <= a(11) and not w19677;
w19679 <= not w19677 and not w19678;
w19680 <= a(11) and not w19678;
w19681 <= not w19679 and not w19680;
w19682 <= w19345 and not w19347;
w19683 <= not w19348 and not w19682;
w19684 <= not w19681 and w19683;
w19685 <= not w19681 and not w19684;
w19686 <= w19683 and not w19684;
w19687 <= not w19685 and not w19686;
w19688 <= w7918 and w12460;
w19689 <= w7226 and w12466;
w19690 <= w7567 and w12463;
w19691 <= not w19689 and not w19690;
w19692 <= not w19688 and w19691;
w19693 <= w7229 and w14543;
w19694 <= w19692 and not w19693;
w19695 <= a(11) and not w19694;
w19696 <= not w19694 and not w19695;
w19697 <= a(11) and not w19695;
w19698 <= not w19696 and not w19697;
w19699 <= not w19340 and not w19344;
w19700 <= not w19343 and not w19344;
w19701 <= not w19699 and not w19700;
w19702 <= not w19698 and not w19701;
w19703 <= not w19698 and not w19702;
w19704 <= not w19701 and not w19702;
w19705 <= not w19703 and not w19704;
w19706 <= w7918 and w12463;
w19707 <= w7226 and w12469;
w19708 <= w7567 and w12466;
w19709 <= not w19707 and not w19708;
w19710 <= not w19706 and w19709;
w19711 <= w7229 and not w14938;
w19712 <= w19710 and not w19711;
w19713 <= a(11) and not w19712;
w19714 <= not w19712 and not w19713;
w19715 <= a(11) and not w19713;
w19716 <= not w19714 and not w19715;
w19717 <= not w19335 and not w19339;
w19718 <= not w19338 and not w19339;
w19719 <= not w19717 and not w19718;
w19720 <= not w19716 and not w19719;
w19721 <= not w19716 and not w19720;
w19722 <= not w19719 and not w19720;
w19723 <= not w19721 and not w19722;
w19724 <= w19121 and w19333;
w19725 <= not w19334 and not w19724;
w19726 <= w7918 and w12466;
w19727 <= w7226 and w12472;
w19728 <= w7567 and w12469;
w19729 <= not w19727 and not w19728;
w19730 <= not w19726 and w19729;
w19731 <= not w7229 and w19730;
w19732 <= not w15190 and w19730;
w19733 <= not w19731 and not w19732;
w19734 <= a(11) and not w19733;
w19735 <= not a(11) and w19733;
w19736 <= not w19734 and not w19735;
w19737 <= w19725 and not w19736;
w19738 <= w19139 and w19331;
w19739 <= not w19332 and not w19738;
w19740 <= w7918 and w12469;
w19741 <= w7226 and w12475;
w19742 <= w7567 and w12472;
w19743 <= not w19741 and not w19742;
w19744 <= not w19740 and w19743;
w19745 <= not w7229 and w19744;
w19746 <= w15031 and w19744;
w19747 <= not w19745 and not w19746;
w19748 <= a(11) and not w19747;
w19749 <= not a(11) and w19747;
w19750 <= not w19748 and not w19749;
w19751 <= w19739 and not w19750;
w19752 <= w19157 and w19329;
w19753 <= not w19330 and not w19752;
w19754 <= w7918 and w12472;
w19755 <= w7226 and w12478;
w19756 <= w7567 and w12475;
w19757 <= not w19755 and not w19756;
w19758 <= not w19754 and w19757;
w19759 <= not w7229 and w19758;
w19760 <= w15320 and w19758;
w19761 <= not w19759 and not w19760;
w19762 <= a(11) and not w19761;
w19763 <= not a(11) and w19761;
w19764 <= not w19762 and not w19763;
w19765 <= w19753 and not w19764;
w19766 <= w7918 and w12475;
w19767 <= w7226 and w12481;
w19768 <= w7567 and w12478;
w19769 <= not w19767 and not w19768;
w19770 <= not w19766 and w19769;
w19771 <= w7229 and not w15643;
w19772 <= w19770 and not w19771;
w19773 <= a(11) and not w19772;
w19774 <= not w19772 and not w19773;
w19775 <= a(11) and not w19773;
w19776 <= not w19774 and not w19775;
w19777 <= w19325 and not w19327;
w19778 <= not w19328 and not w19777;
w19779 <= not w19776 and w19778;
w19780 <= not w19776 and not w19779;
w19781 <= w19778 and not w19779;
w19782 <= not w19780 and not w19781;
w19783 <= w7918 and w12478;
w19784 <= w7226 and w12484;
w19785 <= w7567 and w12481;
w19786 <= not w19784 and not w19785;
w19787 <= not w19783 and w19786;
w19788 <= w7229 and w15659;
w19789 <= w19787 and not w19788;
w19790 <= a(11) and not w19789;
w19791 <= not w19789 and not w19790;
w19792 <= a(11) and not w19790;
w19793 <= not w19791 and not w19792;
w19794 <= not w19320 and not w19324;
w19795 <= not w19323 and not w19324;
w19796 <= not w19794 and not w19795;
w19797 <= not w19793 and not w19796;
w19798 <= not w19793 and not w19797;
w19799 <= not w19796 and not w19797;
w19800 <= not w19798 and not w19799;
w19801 <= w7918 and w12481;
w19802 <= w7226 and w12487;
w19803 <= w7567 and w12484;
w19804 <= not w19802 and not w19803;
w19805 <= not w19801 and w19804;
w19806 <= w7229 and not w15291;
w19807 <= w19805 and not w19806;
w19808 <= a(11) and not w19807;
w19809 <= not w19807 and not w19808;
w19810 <= a(11) and not w19808;
w19811 <= not w19809 and not w19810;
w19812 <= not w19315 and not w19319;
w19813 <= not w19318 and not w19319;
w19814 <= not w19812 and not w19813;
w19815 <= not w19811 and not w19814;
w19816 <= not w19811 and not w19815;
w19817 <= not w19814 and not w19815;
w19818 <= not w19816 and not w19817;
w19819 <= w19216 and w19313;
w19820 <= not w19314 and not w19819;
w19821 <= w7918 and w12484;
w19822 <= w7226 and w12490;
w19823 <= w7567 and w12487;
w19824 <= not w19822 and not w19823;
w19825 <= not w19821 and w19824;
w19826 <= not w7229 and w19825;
w19827 <= not w15699 and w19825;
w19828 <= not w19826 and not w19827;
w19829 <= a(11) and not w19828;
w19830 <= not a(11) and w19828;
w19831 <= not w19829 and not w19830;
w19832 <= w19820 and not w19831;
w19833 <= w19309 and not w19311;
w19834 <= not w19312 and not w19833;
w19835 <= w7918 and w12487;
w19836 <= w7226 and w12493;
w19837 <= w7567 and w12490;
w19838 <= not w19836 and not w19837;
w19839 <= not w19835 and w19838;
w19840 <= not w7229 and w19839;
w19841 <= w15726 and w19839;
w19842 <= not w19840 and not w19841;
w19843 <= a(11) and not w19842;
w19844 <= not a(11) and w19842;
w19845 <= not w19843 and not w19844;
w19846 <= w19834 and not w19845;
w19847 <= w19248 and w19307;
w19848 <= not w19308 and not w19847;
w19849 <= w7918 and w12490;
w19850 <= w7226 and w12496;
w19851 <= w7567 and w12493;
w19852 <= not w19850 and not w19851;
w19853 <= not w19849 and w19852;
w19854 <= not w7229 and w19853;
w19855 <= w15751 and w19853;
w19856 <= not w19854 and not w19855;
w19857 <= a(11) and not w19856;
w19858 <= not a(11) and w19856;
w19859 <= not w19857 and not w19858;
w19860 <= w19848 and not w19859;
w19861 <= w7918 and w12493;
w19862 <= w7226 and w12499;
w19863 <= w7567 and w12496;
w19864 <= not w19862 and not w19863;
w19865 <= not w19861 and w19864;
w19866 <= w7229 and w15782;
w19867 <= w19865 and not w19866;
w19868 <= a(11) and not w19867;
w19869 <= not w19867 and not w19868;
w19870 <= a(11) and not w19868;
w19871 <= not w19869 and not w19870;
w19872 <= w19303 and not w19305;
w19873 <= not w19306 and not w19872;
w19874 <= not w19871 and w19873;
w19875 <= not w19871 and not w19874;
w19876 <= w19873 and not w19874;
w19877 <= not w19875 and not w19876;
w19878 <= not w19290 and not w19302;
w19879 <= not w19301 and not w19302;
w19880 <= not w19878 and not w19879;
w19881 <= w7918 and w12496;
w19882 <= w7226 and w12502;
w19883 <= w7567 and w12499;
w19884 <= not w19882 and not w19883;
w19885 <= not w19881 and w19884;
w19886 <= not w7229 and w19885;
w19887 <= w15840 and w19885;
w19888 <= not w19886 and not w19887;
w19889 <= a(11) and not w19888;
w19890 <= not a(11) and w19888;
w19891 <= not w19889 and not w19890;
w19892 <= not w19880 and not w19891;
w19893 <= w7918 and w12499;
w19894 <= w7226 and w12506;
w19895 <= w7567 and w12502;
w19896 <= not w19894 and not w19895;
w19897 <= not w19893 and w19896;
w19898 <= w7229 and not w15879;
w19899 <= w19897 and not w19898;
w19900 <= a(11) and not w19899;
w19901 <= not w19899 and not w19900;
w19902 <= a(11) and not w19900;
w19903 <= not w19901 and not w19902;
w19904 <= not w19274 and w19285;
w19905 <= not w19286 and not w19904;
w19906 <= not w19903 and w19905;
w19907 <= not w19903 and not w19906;
w19908 <= w19905 and not w19906;
w19909 <= not w19907 and not w19908;
w19910 <= w19271 and not w19273;
w19911 <= not w19274 and not w19910;
w19912 <= w7918 and w12502;
w19913 <= w7226 and w12509;
w19914 <= w7567 and w12506;
w19915 <= not w19913 and not w19914;
w19916 <= not w19912 and w19915;
w19917 <= not w7229 and w19916;
w19918 <= not w15924 and w19916;
w19919 <= not w19917 and not w19918;
w19920 <= a(11) and not w19919;
w19921 <= not a(11) and w19919;
w19922 <= not w19920 and not w19921;
w19923 <= w19911 and not w19922;
w19924 <= w7567 and not w12516;
w19925 <= w7918 and w12512;
w19926 <= not w19924 and not w19925;
w19927 <= w7229 and not w16020;
w19928 <= w19926 and not w19927;
w19929 <= a(11) and not w19928;
w19930 <= a(11) and not w19929;
w19931 <= not w19928 and not w19929;
w19932 <= not w19930 and not w19931;
w19933 <= not w7224 and not w12516;
w19934 <= a(11) and not w19933;
w19935 <= not w19932 and w19934;
w19936 <= w7918 and w12509;
w19937 <= w7226 and not w12516;
w19938 <= w7567 and w12512;
w19939 <= not w19937 and not w19938;
w19940 <= not w19936 and w19939;
w19941 <= not w7229 and w19940;
w19942 <= w16029 and w19940;
w19943 <= not w19941 and not w19942;
w19944 <= a(11) and not w19943;
w19945 <= not a(11) and w19943;
w19946 <= not w19944 and not w19945;
w19947 <= w19935 and not w19946;
w19948 <= w19272 and w19947;
w19949 <= w19947 and not w19948;
w19950 <= w19272 and not w19948;
w19951 <= not w19949 and not w19950;
w19952 <= w7918 and w12506;
w19953 <= w7226 and w12512;
w19954 <= w7567 and w12509;
w19955 <= not w19953 and not w19954;
w19956 <= not w19952 and w19955;
w19957 <= w7229 and w15948;
w19958 <= w19956 and not w19957;
w19959 <= a(11) and not w19958;
w19960 <= a(11) and not w19959;
w19961 <= not w19958 and not w19959;
w19962 <= not w19960 and not w19961;
w19963 <= not w19951 and not w19962;
w19964 <= not w19948 and not w19963;
w19965 <= not w19911 and w19922;
w19966 <= not w19923 and not w19965;
w19967 <= not w19964 and w19966;
w19968 <= not w19923 and not w19967;
w19969 <= not w19909 and not w19968;
w19970 <= not w19906 and not w19969;
w19971 <= w19880 and w19891;
w19972 <= not w19892 and not w19971;
w19973 <= not w19970 and w19972;
w19974 <= not w19892 and not w19973;
w19975 <= not w19877 and not w19974;
w19976 <= not w19874 and not w19975;
w19977 <= w19848 and not w19860;
w19978 <= not w19859 and not w19860;
w19979 <= not w19977 and not w19978;
w19980 <= not w19976 and not w19979;
w19981 <= not w19860 and not w19980;
w19982 <= w19834 and not w19846;
w19983 <= not w19845 and not w19846;
w19984 <= not w19982 and not w19983;
w19985 <= not w19981 and not w19984;
w19986 <= not w19846 and not w19985;
w19987 <= not w19820 and w19831;
w19988 <= not w19832 and not w19987;
w19989 <= not w19986 and w19988;
w19990 <= not w19832 and not w19989;
w19991 <= not w19818 and not w19990;
w19992 <= not w19815 and not w19991;
w19993 <= not w19800 and not w19992;
w19994 <= not w19797 and not w19993;
w19995 <= not w19782 and not w19994;
w19996 <= not w19779 and not w19995;
w19997 <= w19753 and not w19765;
w19998 <= not w19764 and not w19765;
w19999 <= not w19997 and not w19998;
w20000 <= not w19996 and not w19999;
w20001 <= not w19765 and not w20000;
w20002 <= w19739 and not w19751;
w20003 <= not w19750 and not w19751;
w20004 <= not w20002 and not w20003;
w20005 <= not w20001 and not w20004;
w20006 <= not w19751 and not w20005;
w20007 <= not w19725 and w19736;
w20008 <= not w19737 and not w20007;
w20009 <= not w20006 and w20008;
w20010 <= not w19737 and not w20009;
w20011 <= not w19723 and not w20010;
w20012 <= not w19720 and not w20011;
w20013 <= not w19705 and not w20012;
w20014 <= not w19702 and not w20013;
w20015 <= not w19687 and not w20014;
w20016 <= not w19684 and not w20015;
w20017 <= w19658 and not w19670;
w20018 <= not w19669 and not w19670;
w20019 <= not w20017 and not w20018;
w20020 <= not w20016 and not w20019;
w20021 <= not w19670 and not w20020;
w20022 <= not w19644 and w19655;
w20023 <= not w19656 and not w20022;
w20024 <= not w20021 and w20023;
w20025 <= not w19656 and not w20024;
w20026 <= not w19642 and not w20025;
w20027 <= not w19639 and not w20026;
w20028 <= not w19624 and not w20027;
w20029 <= not w19621 and not w20028;
w20030 <= not w19606 and not w20029;
w20031 <= not w19603 and not w20030;
w20032 <= not w19588 and not w20031;
w20033 <= not w19585 and not w20032;
w20034 <= not w19570 and not w20033;
w20035 <= not w19567 and not w20034;
w20036 <= not w19552 and not w20035;
w20037 <= not w19549 and not w20036;
w20038 <= not w19534 and not w20037;
w20039 <= not w19531 and not w20038;
w20040 <= not w19516 and not w20039;
w20041 <= not w19513 and not w20040;
w20042 <= not w19498 and not w20041;
w20043 <= not w19495 and not w20042;
w20044 <= not w19480 and not w20043;
w20045 <= not w19477 and not w20044;
w20046 <= not w19463 and not w20045;
w20047 <= w19463 and w20045;
w20048 <= not w20046 and not w20047;
w20049 <= w9266 and w13565;
w20050 <= w8353 and w13450;
w20051 <= w8795 and w13532;
w20052 <= not w20050 and not w20051;
w20053 <= not w20049 and w20052;
w20054 <= w8356 and w13911;
w20055 <= w20053 and not w20054;
w20056 <= a(8) and not w20055;
w20057 <= a(8) and not w20056;
w20058 <= not w20055 and not w20056;
w20059 <= not w20057 and not w20058;
w20060 <= w20048 and not w20059;
w20061 <= not w20046 and not w20060;
w20062 <= not w19460 and not w20061;
w20063 <= w19460 and w20061;
w20064 <= not w20062 and not w20063;
w20065 <= w6 and not w13373;
w20066 <= w9802 and not w13562;
w20067 <= w10369 and w13876;
w20068 <= not w20066 and not w20067;
w20069 <= not w20065 and w20068;
w20070 <= w9805 and w13963;
w20071 <= w20069 and not w20070;
w20072 <= a(5) and not w20071;
w20073 <= a(5) and not w20072;
w20074 <= not w20071 and not w20072;
w20075 <= not w20073 and not w20074;
w20076 <= w20064 and not w20075;
w20077 <= not w20062 and not w20076;
w20078 <= not w19457 and not w20077;
w20079 <= w19457 and w20077;
w20080 <= not w20078 and not w20079;
w20081 <= w20064 and not w20076;
w20082 <= not w20075 and not w20076;
w20083 <= not w20081 and not w20082;
w20084 <= w20048 and not w20060;
w20085 <= not w20059 and not w20060;
w20086 <= not w20084 and not w20085;
w20087 <= w19480 and w20043;
w20088 <= not w20044 and not w20087;
w20089 <= w9266 and w13532;
w20090 <= w8353 and w13456;
w20091 <= w8795 and w13450;
w20092 <= not w20090 and not w20091;
w20093 <= not w20089 and w20092;
w20094 <= not w8356 and w20093;
w20095 <= w13547 and w20093;
w20096 <= not w20094 and not w20095;
w20097 <= a(8) and not w20096;
w20098 <= not a(8) and w20096;
w20099 <= not w20097 and not w20098;
w20100 <= w20088 and not w20099;
w20101 <= w19498 and w20041;
w20102 <= not w20042 and not w20101;
w20103 <= w9266 and w13450;
w20104 <= w8353 and w13453;
w20105 <= w8795 and w13456;
w20106 <= not w20104 and not w20105;
w20107 <= not w20103 and w20106;
w20108 <= not w8356 and w20107;
w20109 <= not w13476 and w20107;
w20110 <= not w20108 and not w20109;
w20111 <= a(8) and not w20110;
w20112 <= not a(8) and w20110;
w20113 <= not w20111 and not w20112;
w20114 <= w20102 and not w20113;
w20115 <= w19516 and w20039;
w20116 <= not w20040 and not w20115;
w20117 <= w9266 and w13456;
w20118 <= w8353 and w13426;
w20119 <= w8795 and w13453;
w20120 <= not w20118 and not w20119;
w20121 <= not w20117 and w20120;
w20122 <= not w8356 and w20121;
w20123 <= w13844 and w20121;
w20124 <= not w20122 and not w20123;
w20125 <= a(8) and not w20124;
w20126 <= not a(8) and w20124;
w20127 <= not w20125 and not w20126;
w20128 <= w20116 and not w20127;
w20129 <= w19534 and w20037;
w20130 <= not w20038 and not w20129;
w20131 <= w9266 and w13453;
w20132 <= w8353 and w12824;
w20133 <= w8795 and w13426;
w20134 <= not w20132 and not w20133;
w20135 <= not w20131 and w20134;
w20136 <= not w8356 and w20135;
w20137 <= not w13519 and w20135;
w20138 <= not w20136 and not w20137;
w20139 <= a(8) and not w20138;
w20140 <= not a(8) and w20138;
w20141 <= not w20139 and not w20140;
w20142 <= w20130 and not w20141;
w20143 <= w19552 and w20035;
w20144 <= not w20036 and not w20143;
w20145 <= w9266 and w13426;
w20146 <= w8353 and w12704;
w20147 <= w8795 and w12824;
w20148 <= not w20146 and not w20147;
w20149 <= not w20145 and w20148;
w20150 <= not w8356 and w20149;
w20151 <= w13438 and w20149;
w20152 <= not w20150 and not w20151;
w20153 <= a(8) and not w20152;
w20154 <= not a(8) and w20152;
w20155 <= not w20153 and not w20154;
w20156 <= w20144 and not w20155;
w20157 <= w19570 and w20033;
w20158 <= not w20034 and not w20157;
w20159 <= w9266 and w12824;
w20160 <= w8353 and w12437;
w20161 <= w8795 and w12704;
w20162 <= not w20160 and not w20161;
w20163 <= not w20159 and w20162;
w20164 <= not w8356 and w20163;
w20165 <= not w12830 and w20163;
w20166 <= not w20164 and not w20165;
w20167 <= a(8) and not w20166;
w20168 <= not a(8) and w20166;
w20169 <= not w20167 and not w20168;
w20170 <= w20158 and not w20169;
w20171 <= w19588 and w20031;
w20172 <= not w20032 and not w20171;
w20173 <= w9266 and w12704;
w20174 <= w8353 and w12305;
w20175 <= w8795 and w12437;
w20176 <= not w20174 and not w20175;
w20177 <= not w20173 and w20176;
w20178 <= not w8356 and w20177;
w20179 <= not w12934 and w20177;
w20180 <= not w20178 and not w20179;
w20181 <= a(8) and not w20180;
w20182 <= not a(8) and w20180;
w20183 <= not w20181 and not w20182;
w20184 <= w20172 and not w20183;
w20185 <= w19606 and w20029;
w20186 <= not w20030 and not w20185;
w20187 <= w9266 and w12437;
w20188 <= w8353 and w12440;
w20189 <= w8795 and w12305;
w20190 <= not w20188 and not w20189;
w20191 <= not w20187 and w20190;
w20192 <= not w8356 and w20191;
w20193 <= w13671 and w20191;
w20194 <= not w20192 and not w20193;
w20195 <= a(8) and not w20194;
w20196 <= not a(8) and w20194;
w20197 <= not w20195 and not w20196;
w20198 <= w20186 and not w20197;
w20199 <= w19624 and w20027;
w20200 <= not w20028 and not w20199;
w20201 <= w9266 and w12305;
w20202 <= w8353 and w12443;
w20203 <= w8795 and w12440;
w20204 <= not w20202 and not w20203;
w20205 <= not w20201 and w20204;
w20206 <= not w8356 and w20205;
w20207 <= w13683 and w20205;
w20208 <= not w20206 and not w20207;
w20209 <= a(8) and not w20208;
w20210 <= not a(8) and w20208;
w20211 <= not w20209 and not w20210;
w20212 <= w20200 and not w20211;
w20213 <= w19642 and w20025;
w20214 <= not w20026 and not w20213;
w20215 <= w9266 and w12440;
w20216 <= w8353 and w12448;
w20217 <= w8795 and w12443;
w20218 <= not w20216 and not w20217;
w20219 <= not w20215 and w20218;
w20220 <= not w8356 and w20219;
w20221 <= w13986 and w20219;
w20222 <= not w20220 and not w20221;
w20223 <= a(8) and not w20222;
w20224 <= not a(8) and w20222;
w20225 <= not w20223 and not w20224;
w20226 <= w20214 and not w20225;
w20227 <= w9266 and w12443;
w20228 <= w8353 and w12446;
w20229 <= w8795 and w12448;
w20230 <= not w20228 and not w20229;
w20231 <= not w20227 and w20230;
w20232 <= w8356 and w13798;
w20233 <= w20231 and not w20232;
w20234 <= a(8) and not w20233;
w20235 <= not w20233 and not w20234;
w20236 <= a(8) and not w20234;
w20237 <= not w20235 and not w20236;
w20238 <= w20021 and not w20023;
w20239 <= not w20024 and not w20238;
w20240 <= not w20237 and w20239;
w20241 <= not w20237 and not w20240;
w20242 <= w20239 and not w20240;
w20243 <= not w20241 and not w20242;
w20244 <= w9266 and w12448;
w20245 <= w8353 and w12451;
w20246 <= w8795 and w12446;
w20247 <= not w20245 and not w20246;
w20248 <= not w20244 and w20247;
w20249 <= w8356 and w14112;
w20250 <= w20248 and not w20249;
w20251 <= a(8) and not w20250;
w20252 <= not w20250 and not w20251;
w20253 <= a(8) and not w20251;
w20254 <= not w20252 and not w20253;
w20255 <= not w20016 and not w20020;
w20256 <= not w20019 and not w20020;
w20257 <= not w20255 and not w20256;
w20258 <= not w20254 and not w20257;
w20259 <= not w20254 and not w20258;
w20260 <= not w20257 and not w20258;
w20261 <= not w20259 and not w20260;
w20262 <= w19687 and w20014;
w20263 <= not w20015 and not w20262;
w20264 <= w9266 and w12446;
w20265 <= w8353 and w12454;
w20266 <= w8795 and w12451;
w20267 <= not w20265 and not w20266;
w20268 <= not w20264 and w20267;
w20269 <= not w8356 and w20268;
w20270 <= w14168 and w20268;
w20271 <= not w20269 and not w20270;
w20272 <= a(8) and not w20271;
w20273 <= not a(8) and w20271;
w20274 <= not w20272 and not w20273;
w20275 <= w20263 and not w20274;
w20276 <= w19705 and w20012;
w20277 <= not w20013 and not w20276;
w20278 <= w9266 and w12451;
w20279 <= w8353 and w12457;
w20280 <= w8795 and w12454;
w20281 <= not w20279 and not w20280;
w20282 <= not w20278 and w20281;
w20283 <= not w8356 and w20282;
w20284 <= w14378 and w20282;
w20285 <= not w20283 and not w20284;
w20286 <= a(8) and not w20285;
w20287 <= not a(8) and w20285;
w20288 <= not w20286 and not w20287;
w20289 <= w20277 and not w20288;
w20290 <= w19723 and w20010;
w20291 <= not w20011 and not w20290;
w20292 <= w9266 and w12454;
w20293 <= w8353 and w12460;
w20294 <= w8795 and w12457;
w20295 <= not w20293 and not w20294;
w20296 <= not w20292 and w20295;
w20297 <= not w8356 and w20296;
w20298 <= not w14389 and w20296;
w20299 <= not w20297 and not w20298;
w20300 <= a(8) and not w20299;
w20301 <= not a(8) and w20299;
w20302 <= not w20300 and not w20301;
w20303 <= w20291 and not w20302;
w20304 <= w9266 and w12457;
w20305 <= w8353 and w12463;
w20306 <= w8795 and w12460;
w20307 <= not w20305 and not w20306;
w20308 <= not w20304 and w20307;
w20309 <= w8356 and w14772;
w20310 <= w20308 and not w20309;
w20311 <= a(8) and not w20310;
w20312 <= not w20310 and not w20311;
w20313 <= a(8) and not w20311;
w20314 <= not w20312 and not w20313;
w20315 <= w20006 and not w20008;
w20316 <= not w20009 and not w20315;
w20317 <= not w20314 and w20316;
w20318 <= not w20314 and not w20317;
w20319 <= w20316 and not w20317;
w20320 <= not w20318 and not w20319;
w20321 <= w9266 and w12460;
w20322 <= w8353 and w12466;
w20323 <= w8795 and w12463;
w20324 <= not w20322 and not w20323;
w20325 <= not w20321 and w20324;
w20326 <= w8356 and w14543;
w20327 <= w20325 and not w20326;
w20328 <= a(8) and not w20327;
w20329 <= not w20327 and not w20328;
w20330 <= a(8) and not w20328;
w20331 <= not w20329 and not w20330;
w20332 <= not w20001 and not w20005;
w20333 <= not w20004 and not w20005;
w20334 <= not w20332 and not w20333;
w20335 <= not w20331 and not w20334;
w20336 <= not w20331 and not w20335;
w20337 <= not w20334 and not w20335;
w20338 <= not w20336 and not w20337;
w20339 <= w9266 and w12463;
w20340 <= w8353 and w12469;
w20341 <= w8795 and w12466;
w20342 <= not w20340 and not w20341;
w20343 <= not w20339 and w20342;
w20344 <= w8356 and not w14938;
w20345 <= w20343 and not w20344;
w20346 <= a(8) and not w20345;
w20347 <= not w20345 and not w20346;
w20348 <= a(8) and not w20346;
w20349 <= not w20347 and not w20348;
w20350 <= not w19996 and not w20000;
w20351 <= not w19999 and not w20000;
w20352 <= not w20350 and not w20351;
w20353 <= not w20349 and not w20352;
w20354 <= not w20349 and not w20353;
w20355 <= not w20352 and not w20353;
w20356 <= not w20354 and not w20355;
w20357 <= w19782 and w19994;
w20358 <= not w19995 and not w20357;
w20359 <= w9266 and w12466;
w20360 <= w8353 and w12472;
w20361 <= w8795 and w12469;
w20362 <= not w20360 and not w20361;
w20363 <= not w20359 and w20362;
w20364 <= not w8356 and w20363;
w20365 <= not w15190 and w20363;
w20366 <= not w20364 and not w20365;
w20367 <= a(8) and not w20366;
w20368 <= not a(8) and w20366;
w20369 <= not w20367 and not w20368;
w20370 <= w20358 and not w20369;
w20371 <= w19800 and w19992;
w20372 <= not w19993 and not w20371;
w20373 <= w9266 and w12469;
w20374 <= w8353 and w12475;
w20375 <= w8795 and w12472;
w20376 <= not w20374 and not w20375;
w20377 <= not w20373 and w20376;
w20378 <= not w8356 and w20377;
w20379 <= w15031 and w20377;
w20380 <= not w20378 and not w20379;
w20381 <= a(8) and not w20380;
w20382 <= not a(8) and w20380;
w20383 <= not w20381 and not w20382;
w20384 <= w20372 and not w20383;
w20385 <= w19818 and w19990;
w20386 <= not w19991 and not w20385;
w20387 <= w9266 and w12472;
w20388 <= w8353 and w12478;
w20389 <= w8795 and w12475;
w20390 <= not w20388 and not w20389;
w20391 <= not w20387 and w20390;
w20392 <= not w8356 and w20391;
w20393 <= w15320 and w20391;
w20394 <= not w20392 and not w20393;
w20395 <= a(8) and not w20394;
w20396 <= not a(8) and w20394;
w20397 <= not w20395 and not w20396;
w20398 <= w20386 and not w20397;
w20399 <= w9266 and w12475;
w20400 <= w8353 and w12481;
w20401 <= w8795 and w12478;
w20402 <= not w20400 and not w20401;
w20403 <= not w20399 and w20402;
w20404 <= w8356 and not w15643;
w20405 <= w20403 and not w20404;
w20406 <= a(8) and not w20405;
w20407 <= not w20405 and not w20406;
w20408 <= a(8) and not w20406;
w20409 <= not w20407 and not w20408;
w20410 <= w19986 and not w19988;
w20411 <= not w19989 and not w20410;
w20412 <= not w20409 and w20411;
w20413 <= not w20409 and not w20412;
w20414 <= w20411 and not w20412;
w20415 <= not w20413 and not w20414;
w20416 <= w9266 and w12478;
w20417 <= w8353 and w12484;
w20418 <= w8795 and w12481;
w20419 <= not w20417 and not w20418;
w20420 <= not w20416 and w20419;
w20421 <= w8356 and w15659;
w20422 <= w20420 and not w20421;
w20423 <= a(8) and not w20422;
w20424 <= not w20422 and not w20423;
w20425 <= a(8) and not w20423;
w20426 <= not w20424 and not w20425;
w20427 <= not w19981 and not w19985;
w20428 <= not w19984 and not w19985;
w20429 <= not w20427 and not w20428;
w20430 <= not w20426 and not w20429;
w20431 <= not w20426 and not w20430;
w20432 <= not w20429 and not w20430;
w20433 <= not w20431 and not w20432;
w20434 <= w9266 and w12481;
w20435 <= w8353 and w12487;
w20436 <= w8795 and w12484;
w20437 <= not w20435 and not w20436;
w20438 <= not w20434 and w20437;
w20439 <= w8356 and not w15291;
w20440 <= w20438 and not w20439;
w20441 <= a(8) and not w20440;
w20442 <= not w20440 and not w20441;
w20443 <= a(8) and not w20441;
w20444 <= not w20442 and not w20443;
w20445 <= not w19976 and not w19980;
w20446 <= not w19979 and not w19980;
w20447 <= not w20445 and not w20446;
w20448 <= not w20444 and not w20447;
w20449 <= not w20444 and not w20448;
w20450 <= not w20447 and not w20448;
w20451 <= not w20449 and not w20450;
w20452 <= w19877 and w19974;
w20453 <= not w19975 and not w20452;
w20454 <= w9266 and w12484;
w20455 <= w8353 and w12490;
w20456 <= w8795 and w12487;
w20457 <= not w20455 and not w20456;
w20458 <= not w20454 and w20457;
w20459 <= not w8356 and w20458;
w20460 <= not w15699 and w20458;
w20461 <= not w20459 and not w20460;
w20462 <= a(8) and not w20461;
w20463 <= not a(8) and w20461;
w20464 <= not w20462 and not w20463;
w20465 <= w20453 and not w20464;
w20466 <= w19970 and not w19972;
w20467 <= not w19973 and not w20466;
w20468 <= w9266 and w12487;
w20469 <= w8353 and w12493;
w20470 <= w8795 and w12490;
w20471 <= not w20469 and not w20470;
w20472 <= not w20468 and w20471;
w20473 <= not w8356 and w20472;
w20474 <= w15726 and w20472;
w20475 <= not w20473 and not w20474;
w20476 <= a(8) and not w20475;
w20477 <= not a(8) and w20475;
w20478 <= not w20476 and not w20477;
w20479 <= w20467 and not w20478;
w20480 <= w19909 and w19968;
w20481 <= not w19969 and not w20480;
w20482 <= w9266 and w12490;
w20483 <= w8353 and w12496;
w20484 <= w8795 and w12493;
w20485 <= not w20483 and not w20484;
w20486 <= not w20482 and w20485;
w20487 <= not w8356 and w20486;
w20488 <= w15751 and w20486;
w20489 <= not w20487 and not w20488;
w20490 <= a(8) and not w20489;
w20491 <= not a(8) and w20489;
w20492 <= not w20490 and not w20491;
w20493 <= w20481 and not w20492;
w20494 <= w9266 and w12493;
w20495 <= w8353 and w12499;
w20496 <= w8795 and w12496;
w20497 <= not w20495 and not w20496;
w20498 <= not w20494 and w20497;
w20499 <= w8356 and w15782;
w20500 <= w20498 and not w20499;
w20501 <= a(8) and not w20500;
w20502 <= not w20500 and not w20501;
w20503 <= a(8) and not w20501;
w20504 <= not w20502 and not w20503;
w20505 <= w19964 and not w19966;
w20506 <= not w19967 and not w20505;
w20507 <= not w20504 and w20506;
w20508 <= not w20504 and not w20507;
w20509 <= w20506 and not w20507;
w20510 <= not w20508 and not w20509;
w20511 <= not w19951 and not w19963;
w20512 <= not w19962 and not w19963;
w20513 <= not w20511 and not w20512;
w20514 <= w9266 and w12496;
w20515 <= w8353 and w12502;
w20516 <= w8795 and w12499;
w20517 <= not w20515 and not w20516;
w20518 <= not w20514 and w20517;
w20519 <= not w8356 and w20518;
w20520 <= w15840 and w20518;
w20521 <= not w20519 and not w20520;
w20522 <= a(8) and not w20521;
w20523 <= not a(8) and w20521;
w20524 <= not w20522 and not w20523;
w20525 <= not w20513 and not w20524;
w20526 <= w9266 and w12499;
w20527 <= w8353 and w12506;
w20528 <= w8795 and w12502;
w20529 <= not w20527 and not w20528;
w20530 <= not w20526 and w20529;
w20531 <= w8356 and not w15879;
w20532 <= w20530 and not w20531;
w20533 <= a(8) and not w20532;
w20534 <= not w20532 and not w20533;
w20535 <= a(8) and not w20533;
w20536 <= not w20534 and not w20535;
w20537 <= not w19935 and w19946;
w20538 <= not w19947 and not w20537;
w20539 <= not w20536 and w20538;
w20540 <= not w20536 and not w20539;
w20541 <= w20538 and not w20539;
w20542 <= not w20540 and not w20541;
w20543 <= w19932 and not w19934;
w20544 <= not w19935 and not w20543;
w20545 <= w9266 and w12502;
w20546 <= w8353 and w12509;
w20547 <= w8795 and w12506;
w20548 <= not w20546 and not w20547;
w20549 <= not w20545 and w20548;
w20550 <= not w8356 and w20549;
w20551 <= not w15924 and w20549;
w20552 <= not w20550 and not w20551;
w20553 <= a(8) and not w20552;
w20554 <= not a(8) and w20552;
w20555 <= not w20553 and not w20554;
w20556 <= w20544 and not w20555;
w20557 <= w8795 and not w12516;
w20558 <= w9266 and w12512;
w20559 <= not w20557 and not w20558;
w20560 <= w8356 and not w16020;
w20561 <= w20559 and not w20560;
w20562 <= a(8) and not w20561;
w20563 <= a(8) and not w20562;
w20564 <= not w20561 and not w20562;
w20565 <= not w20563 and not w20564;
w20566 <= not w8351 and not w12516;
w20567 <= a(8) and not w20566;
w20568 <= not w20565 and w20567;
w20569 <= w9266 and w12509;
w20570 <= w8353 and not w12516;
w20571 <= w8795 and w12512;
w20572 <= not w20570 and not w20571;
w20573 <= not w20569 and w20572;
w20574 <= not w8356 and w20573;
w20575 <= w16029 and w20573;
w20576 <= not w20574 and not w20575;
w20577 <= a(8) and not w20576;
w20578 <= not a(8) and w20576;
w20579 <= not w20577 and not w20578;
w20580 <= w20568 and not w20579;
w20581 <= w19933 and w20580;
w20582 <= w20580 and not w20581;
w20583 <= w19933 and not w20581;
w20584 <= not w20582 and not w20583;
w20585 <= w9266 and w12506;
w20586 <= w8353 and w12512;
w20587 <= w8795 and w12509;
w20588 <= not w20586 and not w20587;
w20589 <= not w20585 and w20588;
w20590 <= w8356 and w15948;
w20591 <= w20589 and not w20590;
w20592 <= a(8) and not w20591;
w20593 <= a(8) and not w20592;
w20594 <= not w20591 and not w20592;
w20595 <= not w20593 and not w20594;
w20596 <= not w20584 and not w20595;
w20597 <= not w20581 and not w20596;
w20598 <= not w20544 and w20555;
w20599 <= not w20556 and not w20598;
w20600 <= not w20597 and w20599;
w20601 <= not w20556 and not w20600;
w20602 <= not w20542 and not w20601;
w20603 <= not w20539 and not w20602;
w20604 <= w20513 and w20524;
w20605 <= not w20525 and not w20604;
w20606 <= not w20603 and w20605;
w20607 <= not w20525 and not w20606;
w20608 <= not w20510 and not w20607;
w20609 <= not w20507 and not w20608;
w20610 <= w20481 and not w20493;
w20611 <= not w20492 and not w20493;
w20612 <= not w20610 and not w20611;
w20613 <= not w20609 and not w20612;
w20614 <= not w20493 and not w20613;
w20615 <= w20467 and not w20479;
w20616 <= not w20478 and not w20479;
w20617 <= not w20615 and not w20616;
w20618 <= not w20614 and not w20617;
w20619 <= not w20479 and not w20618;
w20620 <= not w20453 and w20464;
w20621 <= not w20465 and not w20620;
w20622 <= not w20619 and w20621;
w20623 <= not w20465 and not w20622;
w20624 <= not w20451 and not w20623;
w20625 <= not w20448 and not w20624;
w20626 <= not w20433 and not w20625;
w20627 <= not w20430 and not w20626;
w20628 <= not w20415 and not w20627;
w20629 <= not w20412 and not w20628;
w20630 <= w20386 and not w20398;
w20631 <= not w20397 and not w20398;
w20632 <= not w20630 and not w20631;
w20633 <= not w20629 and not w20632;
w20634 <= not w20398 and not w20633;
w20635 <= w20372 and not w20384;
w20636 <= not w20383 and not w20384;
w20637 <= not w20635 and not w20636;
w20638 <= not w20634 and not w20637;
w20639 <= not w20384 and not w20638;
w20640 <= not w20358 and w20369;
w20641 <= not w20370 and not w20640;
w20642 <= not w20639 and w20641;
w20643 <= not w20370 and not w20642;
w20644 <= not w20356 and not w20643;
w20645 <= not w20353 and not w20644;
w20646 <= not w20338 and not w20645;
w20647 <= not w20335 and not w20646;
w20648 <= not w20320 and not w20647;
w20649 <= not w20317 and not w20648;
w20650 <= w20291 and not w20303;
w20651 <= not w20302 and not w20303;
w20652 <= not w20650 and not w20651;
w20653 <= not w20649 and not w20652;
w20654 <= not w20303 and not w20653;
w20655 <= w20277 and not w20289;
w20656 <= not w20288 and not w20289;
w20657 <= not w20655 and not w20656;
w20658 <= not w20654 and not w20657;
w20659 <= not w20289 and not w20658;
w20660 <= not w20263 and w20274;
w20661 <= not w20275 and not w20660;
w20662 <= not w20659 and w20661;
w20663 <= not w20275 and not w20662;
w20664 <= not w20261 and not w20663;
w20665 <= not w20258 and not w20664;
w20666 <= not w20243 and not w20665;
w20667 <= not w20240 and not w20666;
w20668 <= w20214 and not w20226;
w20669 <= not w20225 and not w20226;
w20670 <= not w20668 and not w20669;
w20671 <= not w20667 and not w20670;
w20672 <= not w20226 and not w20671;
w20673 <= w20200 and not w20212;
w20674 <= not w20211 and not w20212;
w20675 <= not w20673 and not w20674;
w20676 <= not w20672 and not w20675;
w20677 <= not w20212 and not w20676;
w20678 <= w20186 and not w20198;
w20679 <= not w20197 and not w20198;
w20680 <= not w20678 and not w20679;
w20681 <= not w20677 and not w20680;
w20682 <= not w20198 and not w20681;
w20683 <= w20172 and not w20184;
w20684 <= not w20183 and not w20184;
w20685 <= not w20683 and not w20684;
w20686 <= not w20682 and not w20685;
w20687 <= not w20184 and not w20686;
w20688 <= w20158 and not w20170;
w20689 <= not w20169 and not w20170;
w20690 <= not w20688 and not w20689;
w20691 <= not w20687 and not w20690;
w20692 <= not w20170 and not w20691;
w20693 <= w20144 and not w20156;
w20694 <= not w20155 and not w20156;
w20695 <= not w20693 and not w20694;
w20696 <= not w20692 and not w20695;
w20697 <= not w20156 and not w20696;
w20698 <= w20130 and not w20142;
w20699 <= not w20141 and not w20142;
w20700 <= not w20698 and not w20699;
w20701 <= not w20697 and not w20700;
w20702 <= not w20142 and not w20701;
w20703 <= w20116 and not w20128;
w20704 <= not w20127 and not w20128;
w20705 <= not w20703 and not w20704;
w20706 <= not w20702 and not w20705;
w20707 <= not w20128 and not w20706;
w20708 <= w20102 and not w20114;
w20709 <= not w20113 and not w20114;
w20710 <= not w20708 and not w20709;
w20711 <= not w20707 and not w20710;
w20712 <= not w20114 and not w20711;
w20713 <= not w20088 and w20099;
w20714 <= not w20100 and not w20713;
w20715 <= not w20712 and w20714;
w20716 <= not w20100 and not w20715;
w20717 <= not w20086 and not w20716;
w20718 <= w20086 and w20716;
w20719 <= not w20717 and not w20718;
w20720 <= w6 and w13876;
w20721 <= w9802 and w13568;
w20722 <= w10369 and not w13562;
w20723 <= not w20721 and not w20722;
w20724 <= not w20720 and w20723;
w20725 <= w9805 and w14071;
w20726 <= w20724 and not w20725;
w20727 <= a(5) and not w20726;
w20728 <= a(5) and not w20727;
w20729 <= not w20726 and not w20727;
w20730 <= not w20728 and not w20729;
w20731 <= w20719 and not w20730;
w20732 <= not w20717 and not w20731;
w20733 <= not w20083 and not w20732;
w20734 <= w20083 and w20732;
w20735 <= not w20733 and not w20734;
w20736 <= w20719 and not w20731;
w20737 <= not w20730 and not w20731;
w20738 <= not w20736 and not w20737;
w20739 <= w6 and not w13562;
w20740 <= w9802 and w13565;
w20741 <= w10369 and w13568;
w20742 <= not w20740 and not w20741;
w20743 <= not w20739 and w20742;
w20744 <= w9805 and not w13589;
w20745 <= w20743 and not w20744;
w20746 <= a(5) and not w20745;
w20747 <= not w20745 and not w20746;
w20748 <= a(5) and not w20746;
w20749 <= not w20747 and not w20748;
w20750 <= w20712 and not w20714;
w20751 <= not w20715 and not w20750;
w20752 <= not w20749 and w20751;
w20753 <= not w20749 and not w20752;
w20754 <= w20751 and not w20752;
w20755 <= not w20753 and not w20754;
w20756 <= not w11650 and not w11662;
w20757 <= not w13373 and not w20756;
w20758 <= w10990 and w13876;
w20759 <= not w20757 and not w20758;
w20760 <= w10992 and not w13886;
w20761 <= w20759 and not w20760;
w20762 <= a(2) and not w20761;
w20763 <= a(2) and not w20762;
w20764 <= not w20761 and not w20762;
w20765 <= not w20763 and not w20764;
w20766 <= not w20755 and not w20765;
w20767 <= not w20752 and not w20766;
w20768 <= not w20738 and not w20767;
w20769 <= w20738 and w20767;
w20770 <= not w20768 and not w20769;
w20771 <= not w20755 and not w20766;
w20772 <= not w20765 and not w20766;
w20773 <= not w20771 and not w20772;
w20774 <= w6 and w13568;
w20775 <= w9802 and w13532;
w20776 <= w10369 and w13565;
w20777 <= not w20775 and not w20776;
w20778 <= not w20774 and w20777;
w20779 <= w9805 and w13864;
w20780 <= w20778 and not w20779;
w20781 <= a(5) and not w20780;
w20782 <= not w20780 and not w20781;
w20783 <= a(5) and not w20781;
w20784 <= not w20782 and not w20783;
w20785 <= not w20707 and not w20711;
w20786 <= not w20710 and not w20711;
w20787 <= not w20785 and not w20786;
w20788 <= not w20784 and not w20787;
w20789 <= not w20784 and not w20788;
w20790 <= not w20787 and not w20788;
w20791 <= not w20789 and not w20790;
w20792 <= w6 and w13565;
w20793 <= w9802 and w13450;
w20794 <= w10369 and w13532;
w20795 <= not w20793 and not w20794;
w20796 <= not w20792 and w20795;
w20797 <= w9805 and w13911;
w20798 <= w20796 and not w20797;
w20799 <= a(5) and not w20798;
w20800 <= not w20798 and not w20799;
w20801 <= a(5) and not w20799;
w20802 <= not w20800 and not w20801;
w20803 <= not w20702 and not w20706;
w20804 <= not w20705 and not w20706;
w20805 <= not w20803 and not w20804;
w20806 <= not w20802 and not w20805;
w20807 <= not w20802 and not w20806;
w20808 <= not w20805 and not w20806;
w20809 <= not w20807 and not w20808;
w20810 <= w6 and w13532;
w20811 <= w9802 and w13456;
w20812 <= w10369 and w13450;
w20813 <= not w20811 and not w20812;
w20814 <= not w20810 and w20813;
w20815 <= w9805 and not w13547;
w20816 <= w20814 and not w20815;
w20817 <= a(5) and not w20816;
w20818 <= not w20816 and not w20817;
w20819 <= a(5) and not w20817;
w20820 <= not w20818 and not w20819;
w20821 <= not w20697 and not w20701;
w20822 <= not w20700 and not w20701;
w20823 <= not w20821 and not w20822;
w20824 <= not w20820 and not w20823;
w20825 <= not w20820 and not w20824;
w20826 <= not w20823 and not w20824;
w20827 <= not w20825 and not w20826;
w20828 <= w6 and w13450;
w20829 <= w9802 and w13453;
w20830 <= w10369 and w13456;
w20831 <= not w20829 and not w20830;
w20832 <= not w20828 and w20831;
w20833 <= w9805 and w13476;
w20834 <= w20832 and not w20833;
w20835 <= a(5) and not w20834;
w20836 <= not w20834 and not w20835;
w20837 <= a(5) and not w20835;
w20838 <= not w20836 and not w20837;
w20839 <= not w20692 and not w20696;
w20840 <= not w20695 and not w20696;
w20841 <= not w20839 and not w20840;
w20842 <= not w20838 and not w20841;
w20843 <= not w20838 and not w20842;
w20844 <= not w20841 and not w20842;
w20845 <= not w20843 and not w20844;
w20846 <= w6 and w13456;
w20847 <= w9802 and w13426;
w20848 <= w10369 and w13453;
w20849 <= not w20847 and not w20848;
w20850 <= not w20846 and w20849;
w20851 <= w9805 and not w13844;
w20852 <= w20850 and not w20851;
w20853 <= a(5) and not w20852;
w20854 <= not w20852 and not w20853;
w20855 <= a(5) and not w20853;
w20856 <= not w20854 and not w20855;
w20857 <= not w20687 and not w20691;
w20858 <= not w20690 and not w20691;
w20859 <= not w20857 and not w20858;
w20860 <= not w20856 and not w20859;
w20861 <= not w20856 and not w20860;
w20862 <= not w20859 and not w20860;
w20863 <= not w20861 and not w20862;
w20864 <= w6 and w13453;
w20865 <= w9802 and w12824;
w20866 <= w10369 and w13426;
w20867 <= not w20865 and not w20866;
w20868 <= not w20864 and w20867;
w20869 <= w9805 and w13519;
w20870 <= w20868 and not w20869;
w20871 <= a(5) and not w20870;
w20872 <= not w20870 and not w20871;
w20873 <= a(5) and not w20871;
w20874 <= not w20872 and not w20873;
w20875 <= not w20682 and not w20686;
w20876 <= not w20685 and not w20686;
w20877 <= not w20875 and not w20876;
w20878 <= not w20874 and not w20877;
w20879 <= not w20874 and not w20878;
w20880 <= not w20877 and not w20878;
w20881 <= not w20879 and not w20880;
w20882 <= w6 and w13426;
w20883 <= w9802 and w12704;
w20884 <= w10369 and w12824;
w20885 <= not w20883 and not w20884;
w20886 <= not w20882 and w20885;
w20887 <= w9805 and not w13438;
w20888 <= w20886 and not w20887;
w20889 <= a(5) and not w20888;
w20890 <= not w20888 and not w20889;
w20891 <= a(5) and not w20889;
w20892 <= not w20890 and not w20891;
w20893 <= not w20677 and not w20681;
w20894 <= not w20680 and not w20681;
w20895 <= not w20893 and not w20894;
w20896 <= not w20892 and not w20895;
w20897 <= not w20892 and not w20896;
w20898 <= not w20895 and not w20896;
w20899 <= not w20897 and not w20898;
w20900 <= w6 and w12824;
w20901 <= w9802 and w12437;
w20902 <= w10369 and w12704;
w20903 <= not w20901 and not w20902;
w20904 <= not w20900 and w20903;
w20905 <= w9805 and w12830;
w20906 <= w20904 and not w20905;
w20907 <= a(5) and not w20906;
w20908 <= not w20906 and not w20907;
w20909 <= a(5) and not w20907;
w20910 <= not w20908 and not w20909;
w20911 <= not w20672 and not w20676;
w20912 <= not w20675 and not w20676;
w20913 <= not w20911 and not w20912;
w20914 <= not w20910 and not w20913;
w20915 <= not w20910 and not w20914;
w20916 <= not w20913 and not w20914;
w20917 <= not w20915 and not w20916;
w20918 <= w6 and w12704;
w20919 <= w9802 and w12305;
w20920 <= w10369 and w12437;
w20921 <= not w20919 and not w20920;
w20922 <= not w20918 and w20921;
w20923 <= w9805 and w12934;
w20924 <= w20922 and not w20923;
w20925 <= a(5) and not w20924;
w20926 <= not w20924 and not w20925;
w20927 <= a(5) and not w20925;
w20928 <= not w20926 and not w20927;
w20929 <= not w20667 and not w20671;
w20930 <= not w20670 and not w20671;
w20931 <= not w20929 and not w20930;
w20932 <= not w20928 and not w20931;
w20933 <= not w20928 and not w20932;
w20934 <= not w20931 and not w20932;
w20935 <= not w20933 and not w20934;
w20936 <= w20243 and w20665;
w20937 <= not w20666 and not w20936;
w20938 <= w6 and w12437;
w20939 <= w9802 and w12440;
w20940 <= w10369 and w12305;
w20941 <= not w20939 and not w20940;
w20942 <= not w20938 and w20941;
w20943 <= not w9805 and w20942;
w20944 <= w13671 and w20942;
w20945 <= not w20943 and not w20944;
w20946 <= a(5) and not w20945;
w20947 <= not a(5) and w20945;
w20948 <= not w20946 and not w20947;
w20949 <= w20937 and not w20948;
w20950 <= w20261 and w20663;
w20951 <= not w20664 and not w20950;
w20952 <= w6 and w12305;
w20953 <= w9802 and w12443;
w20954 <= w10369 and w12440;
w20955 <= not w20953 and not w20954;
w20956 <= not w20952 and w20955;
w20957 <= not w9805 and w20956;
w20958 <= w13683 and w20956;
w20959 <= not w20957 and not w20958;
w20960 <= a(5) and not w20959;
w20961 <= not a(5) and w20959;
w20962 <= not w20960 and not w20961;
w20963 <= w20951 and not w20962;
w20964 <= w6 and w12440;
w20965 <= w9802 and w12448;
w20966 <= w10369 and w12443;
w20967 <= not w20965 and not w20966;
w20968 <= not w20964 and w20967;
w20969 <= w9805 and not w13986;
w20970 <= w20968 and not w20969;
w20971 <= a(5) and not w20970;
w20972 <= not w20970 and not w20971;
w20973 <= a(5) and not w20971;
w20974 <= not w20972 and not w20973;
w20975 <= w20659 and not w20661;
w20976 <= not w20662 and not w20975;
w20977 <= not w20974 and w20976;
w20978 <= not w20974 and not w20977;
w20979 <= w20976 and not w20977;
w20980 <= not w20978 and not w20979;
w20981 <= w6 and w12443;
w20982 <= w9802 and w12446;
w20983 <= w10369 and w12448;
w20984 <= not w20982 and not w20983;
w20985 <= not w20981 and w20984;
w20986 <= w9805 and w13798;
w20987 <= w20985 and not w20986;
w20988 <= a(5) and not w20987;
w20989 <= not w20987 and not w20988;
w20990 <= a(5) and not w20988;
w20991 <= not w20989 and not w20990;
w20992 <= not w20654 and not w20658;
w20993 <= not w20657 and not w20658;
w20994 <= not w20992 and not w20993;
w20995 <= not w20991 and not w20994;
w20996 <= not w20991 and not w20995;
w20997 <= not w20994 and not w20995;
w20998 <= not w20996 and not w20997;
w20999 <= w6 and w12448;
w21000 <= w9802 and w12451;
w21001 <= w10369 and w12446;
w21002 <= not w21000 and not w21001;
w21003 <= not w20999 and w21002;
w21004 <= w9805 and w14112;
w21005 <= w21003 and not w21004;
w21006 <= a(5) and not w21005;
w21007 <= not w21005 and not w21006;
w21008 <= a(5) and not w21006;
w21009 <= not w21007 and not w21008;
w21010 <= not w20649 and not w20653;
w21011 <= not w20652 and not w20653;
w21012 <= not w21010 and not w21011;
w21013 <= not w21009 and not w21012;
w21014 <= not w21009 and not w21013;
w21015 <= not w21012 and not w21013;
w21016 <= not w21014 and not w21015;
w21017 <= w20320 and w20647;
w21018 <= not w20648 and not w21017;
w21019 <= w6 and w12446;
w21020 <= w9802 and w12454;
w21021 <= w10369 and w12451;
w21022 <= not w21020 and not w21021;
w21023 <= not w21019 and w21022;
w21024 <= not w9805 and w21023;
w21025 <= w14168 and w21023;
w21026 <= not w21024 and not w21025;
w21027 <= a(5) and not w21026;
w21028 <= not a(5) and w21026;
w21029 <= not w21027 and not w21028;
w21030 <= w21018 and not w21029;
w21031 <= w20338 and w20645;
w21032 <= not w20646 and not w21031;
w21033 <= w6 and w12451;
w21034 <= w9802 and w12457;
w21035 <= w10369 and w12454;
w21036 <= not w21034 and not w21035;
w21037 <= not w21033 and w21036;
w21038 <= not w9805 and w21037;
w21039 <= w14378 and w21037;
w21040 <= not w21038 and not w21039;
w21041 <= a(5) and not w21040;
w21042 <= not a(5) and w21040;
w21043 <= not w21041 and not w21042;
w21044 <= w21032 and not w21043;
w21045 <= w20356 and w20643;
w21046 <= not w20644 and not w21045;
w21047 <= w6 and w12454;
w21048 <= w9802 and w12460;
w21049 <= w10369 and w12457;
w21050 <= not w21048 and not w21049;
w21051 <= not w21047 and w21050;
w21052 <= not w9805 and w21051;
w21053 <= not w14389 and w21051;
w21054 <= not w21052 and not w21053;
w21055 <= a(5) and not w21054;
w21056 <= not a(5) and w21054;
w21057 <= not w21055 and not w21056;
w21058 <= w21046 and not w21057;
w21059 <= w6 and w12457;
w21060 <= w9802 and w12463;
w21061 <= w10369 and w12460;
w21062 <= not w21060 and not w21061;
w21063 <= not w21059 and w21062;
w21064 <= w9805 and w14772;
w21065 <= w21063 and not w21064;
w21066 <= a(5) and not w21065;
w21067 <= not w21065 and not w21066;
w21068 <= a(5) and not w21066;
w21069 <= not w21067 and not w21068;
w21070 <= w20639 and not w20641;
w21071 <= not w20642 and not w21070;
w21072 <= not w21069 and w21071;
w21073 <= not w21069 and not w21072;
w21074 <= w21071 and not w21072;
w21075 <= not w21073 and not w21074;
w21076 <= w6 and w12460;
w21077 <= w9802 and w12466;
w21078 <= w10369 and w12463;
w21079 <= not w21077 and not w21078;
w21080 <= not w21076 and w21079;
w21081 <= w9805 and w14543;
w21082 <= w21080 and not w21081;
w21083 <= a(5) and not w21082;
w21084 <= not w21082 and not w21083;
w21085 <= a(5) and not w21083;
w21086 <= not w21084 and not w21085;
w21087 <= not w20634 and not w20638;
w21088 <= not w20637 and not w20638;
w21089 <= not w21087 and not w21088;
w21090 <= not w21086 and not w21089;
w21091 <= not w21086 and not w21090;
w21092 <= not w21089 and not w21090;
w21093 <= not w21091 and not w21092;
w21094 <= w6 and w12463;
w21095 <= w9802 and w12469;
w21096 <= w10369 and w12466;
w21097 <= not w21095 and not w21096;
w21098 <= not w21094 and w21097;
w21099 <= w9805 and not w14938;
w21100 <= w21098 and not w21099;
w21101 <= a(5) and not w21100;
w21102 <= not w21100 and not w21101;
w21103 <= a(5) and not w21101;
w21104 <= not w21102 and not w21103;
w21105 <= not w20629 and not w20633;
w21106 <= not w20632 and not w20633;
w21107 <= not w21105 and not w21106;
w21108 <= not w21104 and not w21107;
w21109 <= not w21104 and not w21108;
w21110 <= not w21107 and not w21108;
w21111 <= not w21109 and not w21110;
w21112 <= w20415 and w20627;
w21113 <= not w20628 and not w21112;
w21114 <= w6 and w12466;
w21115 <= w9802 and w12472;
w21116 <= w10369 and w12469;
w21117 <= not w21115 and not w21116;
w21118 <= not w21114 and w21117;
w21119 <= not w9805 and w21118;
w21120 <= not w15190 and w21118;
w21121 <= not w21119 and not w21120;
w21122 <= a(5) and not w21121;
w21123 <= not a(5) and w21121;
w21124 <= not w21122 and not w21123;
w21125 <= w21113 and not w21124;
w21126 <= w20433 and w20625;
w21127 <= not w20626 and not w21126;
w21128 <= w6 and w12469;
w21129 <= w9802 and w12475;
w21130 <= w10369 and w12472;
w21131 <= not w21129 and not w21130;
w21132 <= not w21128 and w21131;
w21133 <= not w9805 and w21132;
w21134 <= w15031 and w21132;
w21135 <= not w21133 and not w21134;
w21136 <= a(5) and not w21135;
w21137 <= not a(5) and w21135;
w21138 <= not w21136 and not w21137;
w21139 <= w21127 and not w21138;
w21140 <= w20451 and w20623;
w21141 <= not w20624 and not w21140;
w21142 <= w6 and w12472;
w21143 <= w9802 and w12478;
w21144 <= w10369 and w12475;
w21145 <= not w21143 and not w21144;
w21146 <= not w21142 and w21145;
w21147 <= not w9805 and w21146;
w21148 <= w15320 and w21146;
w21149 <= not w21147 and not w21148;
w21150 <= a(5) and not w21149;
w21151 <= not a(5) and w21149;
w21152 <= not w21150 and not w21151;
w21153 <= w21141 and not w21152;
w21154 <= w6 and w12475;
w21155 <= w9802 and w12481;
w21156 <= w10369 and w12478;
w21157 <= not w21155 and not w21156;
w21158 <= not w21154 and w21157;
w21159 <= w9805 and not w15643;
w21160 <= w21158 and not w21159;
w21161 <= a(5) and not w21160;
w21162 <= not w21160 and not w21161;
w21163 <= a(5) and not w21161;
w21164 <= not w21162 and not w21163;
w21165 <= w20619 and not w20621;
w21166 <= not w20622 and not w21165;
w21167 <= not w21164 and w21166;
w21168 <= not w21164 and not w21167;
w21169 <= w21166 and not w21167;
w21170 <= not w21168 and not w21169;
w21171 <= w6 and w12478;
w21172 <= w9802 and w12484;
w21173 <= w10369 and w12481;
w21174 <= not w21172 and not w21173;
w21175 <= not w21171 and w21174;
w21176 <= w9805 and w15659;
w21177 <= w21175 and not w21176;
w21178 <= a(5) and not w21177;
w21179 <= not w21177 and not w21178;
w21180 <= a(5) and not w21178;
w21181 <= not w21179 and not w21180;
w21182 <= not w20614 and not w20618;
w21183 <= not w20617 and not w20618;
w21184 <= not w21182 and not w21183;
w21185 <= not w21181 and not w21184;
w21186 <= not w21181 and not w21185;
w21187 <= not w21184 and not w21185;
w21188 <= not w21186 and not w21187;
w21189 <= w6 and w12481;
w21190 <= w9802 and w12487;
w21191 <= w10369 and w12484;
w21192 <= not w21190 and not w21191;
w21193 <= not w21189 and w21192;
w21194 <= w9805 and not w15291;
w21195 <= w21193 and not w21194;
w21196 <= a(5) and not w21195;
w21197 <= not w21195 and not w21196;
w21198 <= a(5) and not w21196;
w21199 <= not w21197 and not w21198;
w21200 <= not w20609 and not w20613;
w21201 <= not w20612 and not w20613;
w21202 <= not w21200 and not w21201;
w21203 <= not w21199 and not w21202;
w21204 <= not w21199 and not w21203;
w21205 <= not w21202 and not w21203;
w21206 <= not w21204 and not w21205;
w21207 <= w20510 and w20607;
w21208 <= not w20608 and not w21207;
w21209 <= w6 and w12484;
w21210 <= w9802 and w12490;
w21211 <= w10369 and w12487;
w21212 <= not w21210 and not w21211;
w21213 <= not w21209 and w21212;
w21214 <= not w9805 and w21213;
w21215 <= not w15699 and w21213;
w21216 <= not w21214 and not w21215;
w21217 <= a(5) and not w21216;
w21218 <= not a(5) and w21216;
w21219 <= not w21217 and not w21218;
w21220 <= w21208 and not w21219;
w21221 <= w20603 and not w20605;
w21222 <= not w20606 and not w21221;
w21223 <= w6 and w12487;
w21224 <= w9802 and w12493;
w21225 <= w10369 and w12490;
w21226 <= not w21224 and not w21225;
w21227 <= not w21223 and w21226;
w21228 <= not w9805 and w21227;
w21229 <= w15726 and w21227;
w21230 <= not w21228 and not w21229;
w21231 <= a(5) and not w21230;
w21232 <= not a(5) and w21230;
w21233 <= not w21231 and not w21232;
w21234 <= w21222 and not w21233;
w21235 <= w20542 and w20601;
w21236 <= not w20602 and not w21235;
w21237 <= w6 and w12490;
w21238 <= w9802 and w12496;
w21239 <= w10369 and w12493;
w21240 <= not w21238 and not w21239;
w21241 <= not w21237 and w21240;
w21242 <= not w9805 and w21241;
w21243 <= w15751 and w21241;
w21244 <= not w21242 and not w21243;
w21245 <= a(5) and not w21244;
w21246 <= not a(5) and w21244;
w21247 <= not w21245 and not w21246;
w21248 <= w21236 and not w21247;
w21249 <= w6 and w12493;
w21250 <= w9802 and w12499;
w21251 <= w10369 and w12496;
w21252 <= not w21250 and not w21251;
w21253 <= not w21249 and w21252;
w21254 <= w9805 and w15782;
w21255 <= w21253 and not w21254;
w21256 <= a(5) and not w21255;
w21257 <= not w21255 and not w21256;
w21258 <= a(5) and not w21256;
w21259 <= not w21257 and not w21258;
w21260 <= w20597 and not w20599;
w21261 <= not w20600 and not w21260;
w21262 <= not w21259 and w21261;
w21263 <= not w21259 and not w21262;
w21264 <= w21261 and not w21262;
w21265 <= not w21263 and not w21264;
w21266 <= not w20584 and not w20596;
w21267 <= not w20595 and not w20596;
w21268 <= not w21266 and not w21267;
w21269 <= w6 and w12496;
w21270 <= w9802 and w12502;
w21271 <= w10369 and w12499;
w21272 <= not w21270 and not w21271;
w21273 <= not w21269 and w21272;
w21274 <= not w9805 and w21273;
w21275 <= w15840 and w21273;
w21276 <= not w21274 and not w21275;
w21277 <= a(5) and not w21276;
w21278 <= not a(5) and w21276;
w21279 <= not w21277 and not w21278;
w21280 <= not w21268 and not w21279;
w21281 <= w6 and w12499;
w21282 <= w9802 and w12506;
w21283 <= w10369 and w12502;
w21284 <= not w21282 and not w21283;
w21285 <= not w21281 and w21284;
w21286 <= w9805 and not w15879;
w21287 <= w21285 and not w21286;
w21288 <= a(5) and not w21287;
w21289 <= not w21287 and not w21288;
w21290 <= a(5) and not w21288;
w21291 <= not w21289 and not w21290;
w21292 <= not w20568 and w20579;
w21293 <= not w20580 and not w21292;
w21294 <= not w21291 and w21293;
w21295 <= not w21291 and not w21294;
w21296 <= w21293 and not w21294;
w21297 <= not w21295 and not w21296;
w21298 <= w20565 and not w20567;
w21299 <= not w20568 and not w21298;
w21300 <= w6 and w12502;
w21301 <= w9802 and w12509;
w21302 <= w10369 and w12506;
w21303 <= not w21301 and not w21302;
w21304 <= not w21300 and w21303;
w21305 <= not w9805 and w21304;
w21306 <= not w15924 and w21304;
w21307 <= not w21305 and not w21306;
w21308 <= a(5) and not w21307;
w21309 <= not a(5) and w21307;
w21310 <= not w21308 and not w21309;
w21311 <= w21299 and not w21310;
w21312 <= w10369 and not w12516;
w21313 <= w6 and w12512;
w21314 <= not w21312 and not w21313;
w21315 <= w9805 and not w16020;
w21316 <= w21314 and not w21315;
w21317 <= a(5) and not w21316;
w21318 <= a(5) and not w21317;
w21319 <= not w21316 and not w21317;
w21320 <= not w21318 and not w21319;
w21321 <= not w5 and not w12516;
w21322 <= a(5) and not w21321;
w21323 <= not w21320 and w21322;
w21324 <= w6 and w12509;
w21325 <= w9802 and not w12516;
w21326 <= w10369 and w12512;
w21327 <= not w21325 and not w21326;
w21328 <= not w21324 and w21327;
w21329 <= not w9805 and w21328;
w21330 <= w16029 and w21328;
w21331 <= not w21329 and not w21330;
w21332 <= a(5) and not w21331;
w21333 <= not a(5) and w21331;
w21334 <= not w21332 and not w21333;
w21335 <= w21323 and not w21334;
w21336 <= w20566 and w21335;
w21337 <= w21335 and not w21336;
w21338 <= w20566 and not w21336;
w21339 <= not w21337 and not w21338;
w21340 <= w6 and w12506;
w21341 <= w9802 and w12512;
w21342 <= w10369 and w12509;
w21343 <= not w21341 and not w21342;
w21344 <= not w21340 and w21343;
w21345 <= w9805 and w15948;
w21346 <= w21344 and not w21345;
w21347 <= a(5) and not w21346;
w21348 <= a(5) and not w21347;
w21349 <= not w21346 and not w21347;
w21350 <= not w21348 and not w21349;
w21351 <= not w21339 and not w21350;
w21352 <= not w21336 and not w21351;
w21353 <= not w21299 and w21310;
w21354 <= not w21311 and not w21353;
w21355 <= not w21352 and w21354;
w21356 <= not w21311 and not w21355;
w21357 <= not w21297 and not w21356;
w21358 <= not w21294 and not w21357;
w21359 <= w21268 and w21279;
w21360 <= not w21280 and not w21359;
w21361 <= not w21358 and w21360;
w21362 <= not w21280 and not w21361;
w21363 <= not w21265 and not w21362;
w21364 <= not w21262 and not w21363;
w21365 <= w21236 and not w21248;
w21366 <= not w21247 and not w21248;
w21367 <= not w21365 and not w21366;
w21368 <= not w21364 and not w21367;
w21369 <= not w21248 and not w21368;
w21370 <= w21222 and not w21234;
w21371 <= not w21233 and not w21234;
w21372 <= not w21370 and not w21371;
w21373 <= not w21369 and not w21372;
w21374 <= not w21234 and not w21373;
w21375 <= not w21208 and w21219;
w21376 <= not w21220 and not w21375;
w21377 <= not w21374 and w21376;
w21378 <= not w21220 and not w21377;
w21379 <= not w21206 and not w21378;
w21380 <= not w21203 and not w21379;
w21381 <= not w21188 and not w21380;
w21382 <= not w21185 and not w21381;
w21383 <= not w21170 and not w21382;
w21384 <= not w21167 and not w21383;
w21385 <= w21141 and not w21153;
w21386 <= not w21152 and not w21153;
w21387 <= not w21385 and not w21386;
w21388 <= not w21384 and not w21387;
w21389 <= not w21153 and not w21388;
w21390 <= w21127 and not w21139;
w21391 <= not w21138 and not w21139;
w21392 <= not w21390 and not w21391;
w21393 <= not w21389 and not w21392;
w21394 <= not w21139 and not w21393;
w21395 <= not w21113 and w21124;
w21396 <= not w21125 and not w21395;
w21397 <= not w21394 and w21396;
w21398 <= not w21125 and not w21397;
w21399 <= not w21111 and not w21398;
w21400 <= not w21108 and not w21399;
w21401 <= not w21093 and not w21400;
w21402 <= not w21090 and not w21401;
w21403 <= not w21075 and not w21402;
w21404 <= not w21072 and not w21403;
w21405 <= w21046 and not w21058;
w21406 <= not w21057 and not w21058;
w21407 <= not w21405 and not w21406;
w21408 <= not w21404 and not w21407;
w21409 <= not w21058 and not w21408;
w21410 <= w21032 and not w21044;
w21411 <= not w21043 and not w21044;
w21412 <= not w21410 and not w21411;
w21413 <= not w21409 and not w21412;
w21414 <= not w21044 and not w21413;
w21415 <= not w21018 and w21029;
w21416 <= not w21030 and not w21415;
w21417 <= not w21414 and w21416;
w21418 <= not w21030 and not w21417;
w21419 <= not w21016 and not w21418;
w21420 <= not w21013 and not w21419;
w21421 <= not w20998 and not w21420;
w21422 <= not w20995 and not w21421;
w21423 <= not w20980 and not w21422;
w21424 <= not w20977 and not w21423;
w21425 <= w20951 and not w20963;
w21426 <= not w20962 and not w20963;
w21427 <= not w21425 and not w21426;
w21428 <= not w21424 and not w21427;
w21429 <= not w20963 and not w21428;
w21430 <= not w20937 and w20948;
w21431 <= not w20949 and not w21430;
w21432 <= not w21429 and w21431;
w21433 <= not w20949 and not w21432;
w21434 <= not w20935 and not w21433;
w21435 <= not w20932 and not w21434;
w21436 <= not w20917 and not w21435;
w21437 <= not w20914 and not w21436;
w21438 <= not w20899 and not w21437;
w21439 <= not w20896 and not w21438;
w21440 <= not w20881 and not w21439;
w21441 <= not w20878 and not w21440;
w21442 <= not w20863 and not w21441;
w21443 <= not w20860 and not w21442;
w21444 <= not w20845 and not w21443;
w21445 <= not w20842 and not w21444;
w21446 <= not w20827 and not w21445;
w21447 <= not w20824 and not w21446;
w21448 <= not w20809 and not w21447;
w21449 <= not w20806 and not w21448;
w21450 <= not w20791 and not w21449;
w21451 <= not w20788 and not w21450;
w21452 <= not w20773 and not w21451;
w21453 <= w20773 and w21451;
w21454 <= not w21452 and not w21453;
w21455 <= w20791 and w21449;
w21456 <= not w21450 and not w21455;
w21457 <= w11662 and not w13373;
w21458 <= w10990 and not w13562;
w21459 <= w11650 and w13876;
w21460 <= not w21458 and not w21459;
w21461 <= not w21457 and w21460;
w21462 <= not w10992 and w21461;
w21463 <= not w13963 and w21461;
w21464 <= not w21462 and not w21463;
w21465 <= a(2) and not w21464;
w21466 <= not a(2) and w21464;
w21467 <= not w21465 and not w21466;
w21468 <= w21456 and not w21467;
w21469 <= w20809 and w21447;
w21470 <= not w21448 and not w21469;
w21471 <= w11662 and w13876;
w21472 <= w10990 and w13568;
w21473 <= w11650 and not w13562;
w21474 <= not w21472 and not w21473;
w21475 <= not w21471 and w21474;
w21476 <= not w10992 and w21475;
w21477 <= not w14071 and w21475;
w21478 <= not w21476 and not w21477;
w21479 <= a(2) and not w21478;
w21480 <= not a(2) and w21478;
w21481 <= not w21479 and not w21480;
w21482 <= w21470 and not w21481;
w21483 <= w20827 and w21445;
w21484 <= not w21446 and not w21483;
w21485 <= w11662 and not w13562;
w21486 <= w10990 and w13565;
w21487 <= w11650 and w13568;
w21488 <= not w21486 and not w21487;
w21489 <= not w21485 and w21488;
w21490 <= not w10992 and w21489;
w21491 <= w13589 and w21489;
w21492 <= not w21490 and not w21491;
w21493 <= a(2) and not w21492;
w21494 <= not a(2) and w21492;
w21495 <= not w21493 and not w21494;
w21496 <= w21484 and not w21495;
w21497 <= w20845 and w21443;
w21498 <= not w21444 and not w21497;
w21499 <= w11662 and w13568;
w21500 <= w10990 and w13532;
w21501 <= w11650 and w13565;
w21502 <= not w21500 and not w21501;
w21503 <= not w21499 and w21502;
w21504 <= not w10992 and w21503;
w21505 <= not w13864 and w21503;
w21506 <= not w21504 and not w21505;
w21507 <= a(2) and not w21506;
w21508 <= not a(2) and w21506;
w21509 <= not w21507 and not w21508;
w21510 <= w21498 and not w21509;
w21511 <= w20863 and w21441;
w21512 <= not w21442 and not w21511;
w21513 <= w11662 and w13565;
w21514 <= w10990 and w13450;
w21515 <= w11650 and w13532;
w21516 <= not w21514 and not w21515;
w21517 <= not w21513 and w21516;
w21518 <= not w10992 and w21517;
w21519 <= not w13911 and w21517;
w21520 <= not w21518 and not w21519;
w21521 <= a(2) and not w21520;
w21522 <= not a(2) and w21520;
w21523 <= not w21521 and not w21522;
w21524 <= w21512 and not w21523;
w21525 <= w20881 and w21439;
w21526 <= not w21440 and not w21525;
w21527 <= w11662 and w13532;
w21528 <= w10990 and w13456;
w21529 <= w11650 and w13450;
w21530 <= not w21528 and not w21529;
w21531 <= not w21527 and w21530;
w21532 <= not w10992 and w21531;
w21533 <= w13547 and w21531;
w21534 <= not w21532 and not w21533;
w21535 <= a(2) and not w21534;
w21536 <= not a(2) and w21534;
w21537 <= not w21535 and not w21536;
w21538 <= w21526 and not w21537;
w21539 <= w20899 and w21437;
w21540 <= not w21438 and not w21539;
w21541 <= w11662 and w13450;
w21542 <= w10990 and w13453;
w21543 <= w11650 and w13456;
w21544 <= not w21542 and not w21543;
w21545 <= not w21541 and w21544;
w21546 <= not w10992 and w21545;
w21547 <= not w13476 and w21545;
w21548 <= not w21546 and not w21547;
w21549 <= a(2) and not w21548;
w21550 <= not a(2) and w21548;
w21551 <= not w21549 and not w21550;
w21552 <= w21540 and not w21551;
w21553 <= w20917 and w21435;
w21554 <= not w21436 and not w21553;
w21555 <= w11662 and w13456;
w21556 <= w10990 and w13426;
w21557 <= w11650 and w13453;
w21558 <= not w21556 and not w21557;
w21559 <= not w21555 and w21558;
w21560 <= not w10992 and w21559;
w21561 <= w13844 and w21559;
w21562 <= not w21560 and not w21561;
w21563 <= a(2) and not w21562;
w21564 <= not a(2) and w21562;
w21565 <= not w21563 and not w21564;
w21566 <= w21554 and not w21565;
w21567 <= w20935 and w21433;
w21568 <= not w21434 and not w21567;
w21569 <= w11662 and w13453;
w21570 <= w10990 and w12824;
w21571 <= w11650 and w13426;
w21572 <= not w21570 and not w21571;
w21573 <= not w21569 and w21572;
w21574 <= not w10992 and w21573;
w21575 <= not w13519 and w21573;
w21576 <= not w21574 and not w21575;
w21577 <= a(2) and not w21576;
w21578 <= not a(2) and w21576;
w21579 <= not w21577 and not w21578;
w21580 <= w21568 and not w21579;
w21581 <= w21429 and not w21431;
w21582 <= not w21432 and not w21581;
w21583 <= w21414 and not w21416;
w21584 <= not w21417 and not w21583;
w21585 <= w21394 and not w21396;
w21586 <= not w21397 and not w21585;
w21587 <= w21374 and not w21376;
w21588 <= not w21377 and not w21587;
w21589 <= w21352 and not w21354;
w21590 <= not w21355 and not w21589;
w21591 <= not w21323 and w21334;
w21592 <= not w21335 and not w21591;
w21593 <= not w11729 and not w12516;
w21594 <= w11731 and not w16029;
w21595 <= w11662 and w12509;
w21596 <= w10990 and not w12516;
w21597 <= w11650 and w12512;
w21598 <= not w21596 and not w21597;
w21599 <= not w21595 and w21598;
w21600 <= a(2) and not w21599;
w21601 <= w11731 and not w16020;
w21602 <= w11740 and not w12516;
w21603 <= w11742 and w12512;
w21604 <= a(2) and not w21603;
w21605 <= not w21602 and w21604;
w21606 <= not w21601 and w21605;
w21607 <= not w21600 and w21606;
w21608 <= not w21594 and w21607;
w21609 <= not w21593 and w21608;
w21610 <= w21321 and w21609;
w21611 <= not w21321 and not w21609;
w21612 <= w11662 and w12506;
w21613 <= w10990 and w12512;
w21614 <= w11650 and w12509;
w21615 <= not w21613 and not w21614;
w21616 <= not w21612 and w21615;
w21617 <= w10992 and w15948;
w21618 <= w21616 and not w21617;
w21619 <= not a(2) and not w21618;
w21620 <= a(2) and w21618;
w21621 <= not w21619 and not w21620;
w21622 <= not w21611 and not w21621;
w21623 <= not w21610 and not w21622;
w21624 <= w11662 and w12502;
w21625 <= w10990 and w12509;
w21626 <= w11650 and w12506;
w21627 <= not w21625 and not w21626;
w21628 <= not w21624 and w21627;
w21629 <= not w10992 and w21628;
w21630 <= not w15924 and w21628;
w21631 <= not w21629 and not w21630;
w21632 <= a(2) and not w21631;
w21633 <= not a(2) and w21631;
w21634 <= not w21632 and not w21633;
w21635 <= w21623 and w21634;
w21636 <= w21320 and not w21322;
w21637 <= not w21323 and not w21636;
w21638 <= not w21635 and w21637;
w21639 <= not w21623 and not w21634;
w21640 <= not w21638 and not w21639;
w21641 <= w21592 and not w21640;
w21642 <= not w21592 and w21640;
w21643 <= w11662 and w12499;
w21644 <= w10990 and w12506;
w21645 <= w11650 and w12502;
w21646 <= not w21644 and not w21645;
w21647 <= not w21643 and w21646;
w21648 <= w10992 and not w15879;
w21649 <= w21647 and not w21648;
w21650 <= not a(2) and not w21649;
w21651 <= a(2) and w21649;
w21652 <= not w21650 and not w21651;
w21653 <= not w21642 and not w21652;
w21654 <= not w21641 and not w21653;
w21655 <= w11662 and w12496;
w21656 <= w10990 and w12502;
w21657 <= w11650 and w12499;
w21658 <= not w21656 and not w21657;
w21659 <= not w21655 and w21658;
w21660 <= not w10992 and w21659;
w21661 <= w15840 and w21659;
w21662 <= not w21660 and not w21661;
w21663 <= a(2) and not w21662;
w21664 <= not a(2) and w21662;
w21665 <= not w21663 and not w21664;
w21666 <= not w21654 and not w21665;
w21667 <= w21654 and w21665;
w21668 <= w21339 and w21350;
w21669 <= not w21351 and not w21668;
w21670 <= not w21667 and w21669;
w21671 <= not w21666 and not w21670;
w21672 <= w21590 and not w21671;
w21673 <= not w21590 and w21671;
w21674 <= w11662 and w12493;
w21675 <= w10990 and w12499;
w21676 <= w11650 and w12496;
w21677 <= not w21675 and not w21676;
w21678 <= not w21674 and w21677;
w21679 <= w10992 and w15782;
w21680 <= w21678 and not w21679;
w21681 <= not a(2) and not w21680;
w21682 <= a(2) and w21680;
w21683 <= not w21681 and not w21682;
w21684 <= not w21673 and not w21683;
w21685 <= not w21672 and not w21684;
w21686 <= w11662 and w12490;
w21687 <= w10990 and w12496;
w21688 <= w11650 and w12493;
w21689 <= not w21687 and not w21688;
w21690 <= not w21686 and w21689;
w21691 <= not w10992 and w21690;
w21692 <= w15751 and w21690;
w21693 <= not w21691 and not w21692;
w21694 <= a(2) and not w21693;
w21695 <= not a(2) and w21693;
w21696 <= not w21694 and not w21695;
w21697 <= w21685 and w21696;
w21698 <= w21297 and w21356;
w21699 <= not w21357 and not w21698;
w21700 <= not w21697 and w21699;
w21701 <= not w21685 and not w21696;
w21702 <= not w21700 and not w21701;
w21703 <= w11662 and w12487;
w21704 <= w10990 and w12493;
w21705 <= w11650 and w12490;
w21706 <= not w21704 and not w21705;
w21707 <= not w21703 and w21706;
w21708 <= not w10992 and w21707;
w21709 <= w15726 and w21707;
w21710 <= not w21708 and not w21709;
w21711 <= a(2) and not w21710;
w21712 <= not a(2) and w21710;
w21713 <= not w21711 and not w21712;
w21714 <= w21702 and w21713;
w21715 <= w21358 and not w21360;
w21716 <= not w21361 and not w21715;
w21717 <= not w21714 and w21716;
w21718 <= not w21702 and not w21713;
w21719 <= not w21717 and not w21718;
w21720 <= w11662 and w12484;
w21721 <= w10990 and w12490;
w21722 <= w11650 and w12487;
w21723 <= not w21721 and not w21722;
w21724 <= not w21720 and w21723;
w21725 <= not w10992 and w21724;
w21726 <= not w15699 and w21724;
w21727 <= not w21725 and not w21726;
w21728 <= a(2) and not w21727;
w21729 <= not a(2) and w21727;
w21730 <= not w21728 and not w21729;
w21731 <= w21719 and w21730;
w21732 <= w21265 and w21362;
w21733 <= not w21363 and not w21732;
w21734 <= not w21731 and w21733;
w21735 <= not w21719 and not w21730;
w21736 <= not w21734 and not w21735;
w21737 <= w21364 and not w21366;
w21738 <= not w21365 and w21737;
w21739 <= not w21368 and not w21738;
w21740 <= not w21736 and w21739;
w21741 <= w21736 and not w21739;
w21742 <= w11662 and w12481;
w21743 <= w10990 and w12487;
w21744 <= w11650 and w12484;
w21745 <= not w21743 and not w21744;
w21746 <= not w21742 and w21745;
w21747 <= w10992 and not w15291;
w21748 <= w21746 and not w21747;
w21749 <= not a(2) and not w21748;
w21750 <= a(2) and w21748;
w21751 <= not w21749 and not w21750;
w21752 <= not w21741 and not w21751;
w21753 <= not w21740 and not w21752;
w21754 <= w21369 and not w21371;
w21755 <= not w21370 and w21754;
w21756 <= not w21373 and not w21755;
w21757 <= not w21753 and w21756;
w21758 <= w21753 and not w21756;
w21759 <= w11662 and w12478;
w21760 <= w10990 and w12484;
w21761 <= w11650 and w12481;
w21762 <= not w21760 and not w21761;
w21763 <= not w21759 and w21762;
w21764 <= w10992 and w15659;
w21765 <= w21763 and not w21764;
w21766 <= not a(2) and not w21765;
w21767 <= a(2) and w21765;
w21768 <= not w21766 and not w21767;
w21769 <= not w21758 and not w21768;
w21770 <= not w21757 and not w21769;
w21771 <= w21588 and not w21770;
w21772 <= not w21588 and w21770;
w21773 <= w11662 and w12475;
w21774 <= w10990 and w12481;
w21775 <= w11650 and w12478;
w21776 <= not w21774 and not w21775;
w21777 <= not w21773 and w21776;
w21778 <= w10992 and not w15643;
w21779 <= w21777 and not w21778;
w21780 <= not a(2) and not w21779;
w21781 <= a(2) and w21779;
w21782 <= not w21780 and not w21781;
w21783 <= not w21772 and not w21782;
w21784 <= not w21771 and not w21783;
w21785 <= w11662 and w12472;
w21786 <= w10990 and w12478;
w21787 <= w11650 and w12475;
w21788 <= not w21786 and not w21787;
w21789 <= not w21785 and w21788;
w21790 <= not w10992 and w21789;
w21791 <= w15320 and w21789;
w21792 <= not w21790 and not w21791;
w21793 <= a(2) and not w21792;
w21794 <= not a(2) and w21792;
w21795 <= not w21793 and not w21794;
w21796 <= w21784 and w21795;
w21797 <= w21206 and w21378;
w21798 <= not w21379 and not w21797;
w21799 <= not w21796 and w21798;
w21800 <= not w21784 and not w21795;
w21801 <= not w21799 and not w21800;
w21802 <= w11662 and w12469;
w21803 <= w10990 and w12475;
w21804 <= w11650 and w12472;
w21805 <= not w21803 and not w21804;
w21806 <= not w21802 and w21805;
w21807 <= not w10992 and w21806;
w21808 <= w15031 and w21806;
w21809 <= not w21807 and not w21808;
w21810 <= a(2) and not w21809;
w21811 <= not a(2) and w21809;
w21812 <= not w21810 and not w21811;
w21813 <= w21801 and w21812;
w21814 <= w21188 and w21380;
w21815 <= not w21381 and not w21814;
w21816 <= not w21813 and w21815;
w21817 <= not w21801 and not w21812;
w21818 <= not w21816 and not w21817;
w21819 <= w11662 and w12466;
w21820 <= w10990 and w12472;
w21821 <= w11650 and w12469;
w21822 <= not w21820 and not w21821;
w21823 <= not w21819 and w21822;
w21824 <= not w10992 and w21823;
w21825 <= not w15190 and w21823;
w21826 <= not w21824 and not w21825;
w21827 <= a(2) and not w21826;
w21828 <= not a(2) and w21826;
w21829 <= not w21827 and not w21828;
w21830 <= w21818 and w21829;
w21831 <= w21170 and w21382;
w21832 <= not w21383 and not w21831;
w21833 <= not w21830 and w21832;
w21834 <= not w21818 and not w21829;
w21835 <= not w21833 and not w21834;
w21836 <= w21384 and not w21386;
w21837 <= not w21385 and w21836;
w21838 <= not w21388 and not w21837;
w21839 <= not w21835 and w21838;
w21840 <= w21835 and not w21838;
w21841 <= w11662 and w12463;
w21842 <= w10990 and w12469;
w21843 <= w11650 and w12466;
w21844 <= not w21842 and not w21843;
w21845 <= not w21841 and w21844;
w21846 <= w10992 and not w14938;
w21847 <= w21845 and not w21846;
w21848 <= not a(2) and not w21847;
w21849 <= a(2) and w21847;
w21850 <= not w21848 and not w21849;
w21851 <= not w21840 and not w21850;
w21852 <= not w21839 and not w21851;
w21853 <= w21389 and not w21391;
w21854 <= not w21390 and w21853;
w21855 <= not w21393 and not w21854;
w21856 <= not w21852 and w21855;
w21857 <= w21852 and not w21855;
w21858 <= w11662 and w12460;
w21859 <= w10990 and w12466;
w21860 <= w11650 and w12463;
w21861 <= not w21859 and not w21860;
w21862 <= not w21858 and w21861;
w21863 <= w10992 and w14543;
w21864 <= w21862 and not w21863;
w21865 <= not a(2) and not w21864;
w21866 <= a(2) and w21864;
w21867 <= not w21865 and not w21866;
w21868 <= not w21857 and not w21867;
w21869 <= not w21856 and not w21868;
w21870 <= w21586 and not w21869;
w21871 <= not w21586 and w21869;
w21872 <= w11662 and w12457;
w21873 <= w10990 and w12463;
w21874 <= w11650 and w12460;
w21875 <= not w21873 and not w21874;
w21876 <= not w21872 and w21875;
w21877 <= w10992 and w14772;
w21878 <= w21876 and not w21877;
w21879 <= not a(2) and not w21878;
w21880 <= a(2) and w21878;
w21881 <= not w21879 and not w21880;
w21882 <= not w21871 and not w21881;
w21883 <= not w21870 and not w21882;
w21884 <= w11662 and w12454;
w21885 <= w10990 and w12460;
w21886 <= w11650 and w12457;
w21887 <= not w21885 and not w21886;
w21888 <= not w21884 and w21887;
w21889 <= not w10992 and w21888;
w21890 <= not w14389 and w21888;
w21891 <= not w21889 and not w21890;
w21892 <= a(2) and not w21891;
w21893 <= not a(2) and w21891;
w21894 <= not w21892 and not w21893;
w21895 <= w21883 and w21894;
w21896 <= w21111 and w21398;
w21897 <= not w21399 and not w21896;
w21898 <= not w21895 and w21897;
w21899 <= not w21883 and not w21894;
w21900 <= not w21898 and not w21899;
w21901 <= w11662 and w12451;
w21902 <= w10990 and w12457;
w21903 <= w11650 and w12454;
w21904 <= not w21902 and not w21903;
w21905 <= not w21901 and w21904;
w21906 <= not w10992 and w21905;
w21907 <= w14378 and w21905;
w21908 <= not w21906 and not w21907;
w21909 <= a(2) and not w21908;
w21910 <= not a(2) and w21908;
w21911 <= not w21909 and not w21910;
w21912 <= w21900 and w21911;
w21913 <= w21093 and w21400;
w21914 <= not w21401 and not w21913;
w21915 <= not w21912 and w21914;
w21916 <= not w21900 and not w21911;
w21917 <= not w21915 and not w21916;
w21918 <= w11662 and w12446;
w21919 <= w10990 and w12454;
w21920 <= w11650 and w12451;
w21921 <= not w21919 and not w21920;
w21922 <= not w21918 and w21921;
w21923 <= not w10992 and w21922;
w21924 <= w14168 and w21922;
w21925 <= not w21923 and not w21924;
w21926 <= a(2) and not w21925;
w21927 <= not a(2) and w21925;
w21928 <= not w21926 and not w21927;
w21929 <= w21917 and w21928;
w21930 <= w21075 and w21402;
w21931 <= not w21403 and not w21930;
w21932 <= not w21929 and w21931;
w21933 <= not w21917 and not w21928;
w21934 <= not w21932 and not w21933;
w21935 <= w21404 and not w21406;
w21936 <= not w21405 and w21935;
w21937 <= not w21408 and not w21936;
w21938 <= not w21934 and w21937;
w21939 <= w21934 and not w21937;
w21940 <= w11662 and w12448;
w21941 <= w10990 and w12451;
w21942 <= w11650 and w12446;
w21943 <= not w21941 and not w21942;
w21944 <= not w21940 and w21943;
w21945 <= w10992 and w14112;
w21946 <= w21944 and not w21945;
w21947 <= not a(2) and not w21946;
w21948 <= a(2) and w21946;
w21949 <= not w21947 and not w21948;
w21950 <= not w21939 and not w21949;
w21951 <= not w21938 and not w21950;
w21952 <= w21409 and not w21411;
w21953 <= not w21410 and w21952;
w21954 <= not w21413 and not w21953;
w21955 <= not w21951 and w21954;
w21956 <= w21951 and not w21954;
w21957 <= w11662 and w12443;
w21958 <= w10990 and w12446;
w21959 <= w11650 and w12448;
w21960 <= not w21958 and not w21959;
w21961 <= not w21957 and w21960;
w21962 <= w10992 and w13798;
w21963 <= w21961 and not w21962;
w21964 <= not a(2) and not w21963;
w21965 <= a(2) and w21963;
w21966 <= not w21964 and not w21965;
w21967 <= not w21956 and not w21966;
w21968 <= not w21955 and not w21967;
w21969 <= w21584 and not w21968;
w21970 <= not w21584 and w21968;
w21971 <= w11662 and w12440;
w21972 <= w10990 and w12448;
w21973 <= w11650 and w12443;
w21974 <= not w21972 and not w21973;
w21975 <= not w21971 and w21974;
w21976 <= w10992 and not w13986;
w21977 <= w21975 and not w21976;
w21978 <= not a(2) and not w21977;
w21979 <= a(2) and w21977;
w21980 <= not w21978 and not w21979;
w21981 <= not w21970 and not w21980;
w21982 <= not w21969 and not w21981;
w21983 <= w11662 and w12305;
w21984 <= w10990 and w12443;
w21985 <= w11650 and w12440;
w21986 <= not w21984 and not w21985;
w21987 <= not w21983 and w21986;
w21988 <= not w10992 and w21987;
w21989 <= w13683 and w21987;
w21990 <= not w21988 and not w21989;
w21991 <= a(2) and not w21990;
w21992 <= not a(2) and w21990;
w21993 <= not w21991 and not w21992;
w21994 <= w21982 and w21993;
w21995 <= w21016 and w21418;
w21996 <= not w21419 and not w21995;
w21997 <= not w21994 and w21996;
w21998 <= not w21982 and not w21993;
w21999 <= not w21997 and not w21998;
w22000 <= w11662 and w12437;
w22001 <= w10990 and w12440;
w22002 <= w11650 and w12305;
w22003 <= not w22001 and not w22002;
w22004 <= not w22000 and w22003;
w22005 <= not w10992 and w22004;
w22006 <= w13671 and w22004;
w22007 <= not w22005 and not w22006;
w22008 <= a(2) and not w22007;
w22009 <= not a(2) and w22007;
w22010 <= not w22008 and not w22009;
w22011 <= w21999 and w22010;
w22012 <= w20998 and w21420;
w22013 <= not w21421 and not w22012;
w22014 <= not w22011 and w22013;
w22015 <= not w21999 and not w22010;
w22016 <= not w22014 and not w22015;
w22017 <= w11662 and w12704;
w22018 <= w10990 and w12305;
w22019 <= w11650 and w12437;
w22020 <= not w22018 and not w22019;
w22021 <= not w22017 and w22020;
w22022 <= not w10992 and w22021;
w22023 <= not w12934 and w22021;
w22024 <= not w22022 and not w22023;
w22025 <= a(2) and not w22024;
w22026 <= not a(2) and w22024;
w22027 <= not w22025 and not w22026;
w22028 <= w22016 and w22027;
w22029 <= w20980 and w21422;
w22030 <= not w21423 and not w22029;
w22031 <= not w22028 and w22030;
w22032 <= not w22016 and not w22027;
w22033 <= not w22031 and not w22032;
w22034 <= w21424 and not w21426;
w22035 <= not w21425 and w22034;
w22036 <= not w21428 and not w22035;
w22037 <= not w22033 and w22036;
w22038 <= w22033 and not w22036;
w22039 <= w11662 and w12824;
w22040 <= w10990 and w12437;
w22041 <= w11650 and w12704;
w22042 <= not w22040 and not w22041;
w22043 <= not w22039 and w22042;
w22044 <= w10992 and w12830;
w22045 <= w22043 and not w22044;
w22046 <= not a(2) and not w22045;
w22047 <= a(2) and w22045;
w22048 <= not w22046 and not w22047;
w22049 <= not w22038 and not w22048;
w22050 <= not w22037 and not w22049;
w22051 <= w21582 and not w22050;
w22052 <= not w21582 and w22050;
w22053 <= w11662 and w13426;
w22054 <= w10990 and w12704;
w22055 <= w11650 and w12824;
w22056 <= not w22054 and not w22055;
w22057 <= not w22053 and w22056;
w22058 <= w10992 and not w13438;
w22059 <= w22057 and not w22058;
w22060 <= not a(2) and not w22059;
w22061 <= a(2) and w22059;
w22062 <= not w22060 and not w22061;
w22063 <= not w22052 and not w22062;
w22064 <= not w22051 and not w22063;
w22065 <= w21568 and not w21580;
w22066 <= not w21579 and not w21580;
w22067 <= not w22065 and not w22066;
w22068 <= not w22064 and not w22067;
w22069 <= not w21580 and not w22068;
w22070 <= not w21554 and w21565;
w22071 <= not w21566 and not w22070;
w22072 <= not w22069 and w22071;
w22073 <= not w21566 and not w22072;
w22074 <= not w21540 and w21551;
w22075 <= not w21552 and not w22074;
w22076 <= not w22073 and w22075;
w22077 <= not w21552 and not w22076;
w22078 <= not w21526 and w21537;
w22079 <= not w21538 and not w22078;
w22080 <= not w22077 and w22079;
w22081 <= not w21538 and not w22080;
w22082 <= not w21512 and w21523;
w22083 <= not w21524 and not w22082;
w22084 <= not w22081 and w22083;
w22085 <= not w21524 and not w22084;
w22086 <= not w21498 and w21509;
w22087 <= not w21510 and not w22086;
w22088 <= not w22085 and w22087;
w22089 <= not w21510 and not w22088;
w22090 <= not w21484 and w21495;
w22091 <= not w21496 and not w22090;
w22092 <= not w22089 and w22091;
w22093 <= not w21496 and not w22092;
w22094 <= not w21470 and w21481;
w22095 <= not w21482 and not w22094;
w22096 <= not w22093 and w22095;
w22097 <= not w21482 and not w22096;
w22098 <= not w21456 and w21467;
w22099 <= not w21468 and not w22098;
w22100 <= not w22097 and w22099;
w22101 <= not w21468 and not w22100;
w22102 <= w21454 and not w22101;
w22103 <= not w21452 and not w22102;
w22104 <= w20770 and not w22103;
w22105 <= not w20768 and not w22104;
w22106 <= w20735 and not w22105;
w22107 <= not w20733 and not w22106;
w22108 <= w20080 and not w22107;
w22109 <= not w20078 and not w22108;
w22110 <= w19451 and not w19453;
w22111 <= not w19454 and not w22110;
w22112 <= not w22109 and w22111;
w22113 <= not w19454 and not w22112;
w22114 <= not w18881 and not w22113;
w22115 <= not w18878 and not w22114;
w22116 <= w18331 and not w22115;
w22117 <= not w18329 and not w22116;
w22118 <= w17827 and not w17829;
w22119 <= not w17830 and not w22118;
w22120 <= not w22117 and w22119;
w22121 <= not w17830 and not w22120;
w22122 <= not w17363 and not w22121;
w22123 <= not w17360 and not w22122;
w22124 <= w16936 and not w22123;
w22125 <= not w16934 and not w22124;
w22126 <= w16539 and not w16541;
w22127 <= not w16542 and not w22126;
w22128 <= not w22125 and w22127;
w22129 <= not w16542 and not w22128;
w22130 <= not w16378 and not w22129;
w22131 <= not w16375 and not w22130;
w22132 <= w16207 and not w22131;
w22133 <= not w16205 and not w22132;
w22134 <= w15585 and not w15587;
w22135 <= not w15588 and not w22134;
w22136 <= not w22133 and w22135;
w22137 <= not w15588 and not w22136;
w22138 <= not w15443 and not w22137;
w22139 <= not w15440 and not w22138;
w22140 <= w15138 and not w22139;
w22141 <= not w15136 and not w22140;
w22142 <= w14885 and not w14887;
w22143 <= not w14888 and not w22142;
w22144 <= not w22141 and w22143;
w22145 <= not w14888 and not w22144;
w22146 <= not w14744 and not w22145;
w22147 <= not w14741 and not w22146;
w22148 <= w14631 and not w22147;
w22149 <= not w14629 and not w22148;
w22150 <= w14256 and not w14258;
w22151 <= not w14259 and not w22150;
w22152 <= not w22149 and w22151;
w22153 <= not w14259 and not w22152;
w22154 <= not w14089 and not w22153;
w22155 <= not w14086 and not w22154;
w22156 <= w13974 and not w22155;
w22157 <= not w13972 and not w22156;
w22158 <= not w13892 and not w13895;
w22159 <= not w13556 and not w13596;
w22160 <= w3819 and w13876;
w22161 <= w3902 and w13568;
w22162 <= w3981 and not w13562;
w22163 <= not w22161 and not w22162;
w22164 <= not w22160 and w22163;
w22165 <= w3985 and w14071;
w22166 <= w22164 and not w22165;
w22167 <= a(26) and not w22166;
w22168 <= a(26) and not w22167;
w22169 <= not w22166 and not w22167;
w22170 <= not w22168 and not w22169;
w22171 <= not w22159 and not w22170;
w22172 <= not w22159 and not w22171;
w22173 <= not w22170 and not w22171;
w22174 <= not w22172 and not w22173;
w22175 <= w10 and not w13844;
w22176 <= w2955 and w13456;
w22177 <= w2958 and w13426;
w22178 <= w2963 and w13453;
w22179 <= not w22177 and not w22178;
w22180 <= not w22176 and w22179;
w22181 <= not w22175 and w22180;
w22182 <= not w4468 and w13873;
w22183 <= not w4471 and w22182;
w22184 <= not w13373 and not w22183;
w22185 <= a(23) and not w22184;
w22186 <= not a(23) and w22184;
w22187 <= not w22185 and not w22186;
w22188 <= w238 and w2977;
w22189 <= w6502 and w22188;
w22190 <= w4762 and w22189;
w22191 <= w15966 and w22190;
w22192 <= w13722 and w22191;
w22193 <= w14469 and w22192;
w22194 <= w709 and w22193;
w22195 <= w406 and w22194;
w22196 <= w3668 and w22195;
w22197 <= w1204 and w22196;
w22198 <= not w782 and w22197;
w22199 <= not w302 and w22198;
w22200 <= not w161 and w22199;
w22201 <= not w241 and w22200;
w22202 <= not w93 and w22201;
w22203 <= not w205 and w22202;
w22204 <= w13509 and w22203;
w22205 <= not w13509 and not w22203;
w22206 <= not w22204 and not w22205;
w22207 <= w22187 and w22206;
w22208 <= not w22187 and not w22206;
w22209 <= not w22207 and not w22208;
w22210 <= not w13515 and w22209;
w22211 <= w13515 and not w22209;
w22212 <= not w22210 and not w22211;
w22213 <= not w22181 and w22212;
w22214 <= w22212 and not w22213;
w22215 <= not w22181 and not w22213;
w22216 <= not w22214 and not w22215;
w22217 <= not w13527 and not w13553;
w22218 <= w22216 and w22217;
w22219 <= not w22216 and not w22217;
w22220 <= not w22218 and not w22219;
w22221 <= w3392 and w13565;
w22222 <= w3477 and w13450;
w22223 <= w3541 and w13532;
w22224 <= not w22222 and not w22223;
w22225 <= not w22221 and w22224;
w22226 <= w3303 and w13911;
w22227 <= w22225 and not w22226;
w22228 <= a(29) and not w22227;
w22229 <= a(29) and not w22228;
w22230 <= not w22227 and not w22228;
w22231 <= not w22229 and not w22230;
w22232 <= w22220 and not w22231;
w22233 <= w22220 and not w22232;
w22234 <= not w22231 and not w22232;
w22235 <= not w22233 and not w22234;
w22236 <= not w22174 and w22235;
w22237 <= w22174 and not w22235;
w22238 <= not w22236 and not w22237;
w22239 <= not w22158 and not w22238;
w22240 <= w22158 and w22238;
w22241 <= not w22239 and not w22240;
w22242 <= not w22157 and w22241;
w22243 <= w22157 and not w22241;
w22244 <= not w22242 and not w22243;
w22245 <= w6 and w22244;
w22246 <= w14089 and w22153;
w22247 <= not w22154 and not w22246;
w22248 <= w9802 and w22247;
w22249 <= not w13974 and w22155;
w22250 <= not w22156 and not w22249;
w22251 <= w10369 and w22250;
w22252 <= not w22248 and not w22251;
w22253 <= not w22245 and w22252;
w22254 <= w22149 and not w22151;
w22255 <= not w22152 and not w22254;
w22256 <= w22247 and w22255;
w22257 <= not w14631 and w22147;
w22258 <= not w22148 and not w22257;
w22259 <= w22255 and w22258;
w22260 <= w14744 and w22145;
w22261 <= not w22146 and not w22260;
w22262 <= w22258 and w22261;
w22263 <= w22141 and not w22143;
w22264 <= not w22144 and not w22263;
w22265 <= w22261 and w22264;
w22266 <= not w15138 and w22139;
w22267 <= not w22140 and not w22266;
w22268 <= w22264 and w22267;
w22269 <= w15443 and w22137;
w22270 <= not w22138 and not w22269;
w22271 <= w22267 and w22270;
w22272 <= w22133 and not w22135;
w22273 <= not w22136 and not w22272;
w22274 <= w22270 and w22273;
w22275 <= not w16207 and w22131;
w22276 <= not w22132 and not w22275;
w22277 <= w22273 and w22276;
w22278 <= w16378 and w22129;
w22279 <= not w22130 and not w22278;
w22280 <= w22276 and w22279;
w22281 <= w22125 and not w22127;
w22282 <= not w22128 and not w22281;
w22283 <= w22279 and w22282;
w22284 <= not w16936 and w22123;
w22285 <= not w22124 and not w22284;
w22286 <= w22282 and w22285;
w22287 <= w17363 and w22121;
w22288 <= not w22122 and not w22287;
w22289 <= w22285 and w22288;
w22290 <= w22117 and not w22119;
w22291 <= not w22120 and not w22290;
w22292 <= w22288 and w22291;
w22293 <= not w18331 and w22115;
w22294 <= not w22116 and not w22293;
w22295 <= w22291 and w22294;
w22296 <= w18881 and w22113;
w22297 <= not w22114 and not w22296;
w22298 <= w22294 and w22297;
w22299 <= w22109 and not w22111;
w22300 <= not w22112 and not w22299;
w22301 <= w22297 and w22300;
w22302 <= not w20080 and w22107;
w22303 <= not w22108 and not w22302;
w22304 <= w22300 and w22303;
w22305 <= not w20735 and w22105;
w22306 <= not w22106 and not w22305;
w22307 <= w22303 and w22306;
w22308 <= not w20770 and w22103;
w22309 <= not w22104 and not w22308;
w22310 <= w22306 and w22309;
w22311 <= not w21454 and w22101;
w22312 <= not w22102 and not w22311;
w22313 <= w22309 and w22312;
w22314 <= w22097 and not w22099;
w22315 <= not w22100 and not w22314;
w22316 <= w22312 and w22315;
w22317 <= not w22312 and not w22315;
w22318 <= w22093 and not w22095;
w22319 <= not w22096 and not w22318;
w22320 <= w22315 and w22319;
w22321 <= w22089 and not w22091;
w22322 <= not w22092 and not w22321;
w22323 <= w22319 and w22322;
w22324 <= w22085 and not w22087;
w22325 <= not w22088 and not w22324;
w22326 <= w22322 and w22325;
w22327 <= w22081 and not w22083;
w22328 <= not w22084 and not w22327;
w22329 <= w22325 and w22328;
w22330 <= w22077 and not w22079;
w22331 <= not w22080 and not w22330;
w22332 <= w22328 and w22331;
w22333 <= w22073 and not w22075;
w22334 <= not w22076 and not w22333;
w22335 <= w22331 and w22334;
w22336 <= w22069 and not w22071;
w22337 <= not w22072 and not w22336;
w22338 <= w22334 and w22337;
w22339 <= not w22064 and not w22068;
w22340 <= not w22067 and not w22068;
w22341 <= not w22339 and not w22340;
w22342 <= w22337 and not w22341;
w22343 <= not w22334 and w22342;
w22344 <= not w22338 and not w22343;
w22345 <= not w22331 and not w22334;
w22346 <= not w22335 and not w22345;
w22347 <= not w22344 and w22346;
w22348 <= not w22335 and not w22347;
w22349 <= not w22328 and not w22331;
w22350 <= not w22332 and not w22349;
w22351 <= not w22348 and w22350;
w22352 <= not w22332 and not w22351;
w22353 <= not w22325 and not w22328;
w22354 <= not w22329 and not w22353;
w22355 <= not w22352 and w22354;
w22356 <= not w22329 and not w22355;
w22357 <= not w22322 and not w22325;
w22358 <= not w22326 and not w22357;
w22359 <= not w22356 and w22358;
w22360 <= not w22326 and not w22359;
w22361 <= not w22319 and not w22322;
w22362 <= not w22323 and not w22361;
w22363 <= not w22360 and w22362;
w22364 <= not w22323 and not w22363;
w22365 <= not w22315 and not w22319;
w22366 <= not w22320 and not w22365;
w22367 <= not w22364 and w22366;
w22368 <= not w22320 and not w22367;
w22369 <= not w22316 and not w22368;
w22370 <= not w22317 and w22369;
w22371 <= not w22316 and not w22370;
w22372 <= not w22309 and not w22312;
w22373 <= not w22313 and not w22372;
w22374 <= not w22371 and w22373;
w22375 <= not w22313 and not w22374;
w22376 <= not w22306 and not w22309;
w22377 <= not w22310 and not w22376;
w22378 <= not w22375 and w22377;
w22379 <= not w22310 and not w22378;
w22380 <= not w22303 and not w22306;
w22381 <= not w22307 and not w22380;
w22382 <= not w22379 and w22381;
w22383 <= not w22307 and not w22382;
w22384 <= not w22300 and not w22303;
w22385 <= not w22383 and not w22384;
w22386 <= not w22304 and w22385;
w22387 <= not w22304 and not w22386;
w22388 <= not w22297 and not w22300;
w22389 <= not w22387 and not w22388;
w22390 <= not w22301 and w22389;
w22391 <= not w22301 and not w22390;
w22392 <= not w22294 and not w22297;
w22393 <= not w22298 and not w22392;
w22394 <= not w22391 and w22393;
w22395 <= not w22298 and not w22394;
w22396 <= not w22291 and not w22294;
w22397 <= not w22395 and not w22396;
w22398 <= not w22295 and w22397;
w22399 <= not w22295 and not w22398;
w22400 <= not w22288 and not w22291;
w22401 <= not w22399 and not w22400;
w22402 <= not w22292 and w22401;
w22403 <= not w22292 and not w22402;
w22404 <= not w22285 and not w22288;
w22405 <= not w22289 and not w22404;
w22406 <= not w22403 and w22405;
w22407 <= not w22289 and not w22406;
w22408 <= not w22282 and not w22285;
w22409 <= not w22407 and not w22408;
w22410 <= not w22286 and w22409;
w22411 <= not w22286 and not w22410;
w22412 <= not w22279 and not w22282;
w22413 <= not w22411 and not w22412;
w22414 <= not w22283 and w22413;
w22415 <= not w22283 and not w22414;
w22416 <= not w22276 and not w22279;
w22417 <= not w22280 and not w22416;
w22418 <= not w22415 and w22417;
w22419 <= not w22280 and not w22418;
w22420 <= not w22273 and not w22276;
w22421 <= not w22419 and not w22420;
w22422 <= not w22277 and w22421;
w22423 <= not w22277 and not w22422;
w22424 <= not w22270 and not w22273;
w22425 <= not w22423 and not w22424;
w22426 <= not w22274 and w22425;
w22427 <= not w22274 and not w22426;
w22428 <= not w22267 and not w22270;
w22429 <= not w22271 and not w22428;
w22430 <= not w22427 and w22429;
w22431 <= not w22271 and not w22430;
w22432 <= not w22264 and not w22267;
w22433 <= not w22431 and not w22432;
w22434 <= not w22268 and w22433;
w22435 <= not w22268 and not w22434;
w22436 <= not w22261 and not w22264;
w22437 <= not w22435 and not w22436;
w22438 <= not w22265 and w22437;
w22439 <= not w22265 and not w22438;
w22440 <= not w22258 and not w22261;
w22441 <= not w22262 and not w22440;
w22442 <= not w22439 and w22441;
w22443 <= not w22262 and not w22442;
w22444 <= not w22255 and not w22258;
w22445 <= not w22443 and not w22444;
w22446 <= not w22259 and w22445;
w22447 <= not w22259 and not w22446;
w22448 <= not w22247 and not w22255;
w22449 <= not w22447 and not w22448;
w22450 <= not w22256 and w22449;
w22451 <= not w22256 and not w22450;
w22452 <= not w22247 and not w22250;
w22453 <= w22247 and w22250;
w22454 <= not w22452 and not w22453;
w22455 <= not w22451 and w22454;
w22456 <= not w22453 and not w22455;
w22457 <= w22244 and w22250;
w22458 <= not w22244 and not w22250;
w22459 <= not w22456 and not w22458;
w22460 <= not w22457 and w22459;
w22461 <= not w22456 and not w22460;
w22462 <= not w22457 and not w22460;
w22463 <= not w22458 and w22462;
w22464 <= not w22461 and not w22463;
w22465 <= w9805 and not w22464;
w22466 <= w22253 and not w22465;
w22467 <= a(5) and not w22466;
w22468 <= not w22466 and not w22467;
w22469 <= a(5) and not w22467;
w22470 <= not w22468 and not w22469;
w22471 <= w7918 and w22267;
w22472 <= w7226 and w22273;
w22473 <= w7567 and w22270;
w22474 <= not w22472 and not w22473;
w22475 <= not w22471 and w22474;
w22476 <= w22427 and not w22429;
w22477 <= not w22430 and not w22476;
w22478 <= w7229 and w22477;
w22479 <= w22475 and not w22478;
w22480 <= a(11) and not w22479;
w22481 <= not w22479 and not w22480;
w22482 <= a(11) and not w22480;
w22483 <= not w22481 and not w22482;
w22484 <= w6168 and w22288;
w22485 <= w5598 and w22294;
w22486 <= w5874 and w22291;
w22487 <= not w22485 and not w22486;
w22488 <= not w22484 and w22487;
w22489 <= not w22399 and not w22402;
w22490 <= not w22400 and w22403;
w22491 <= not w22489 and not w22490;
w22492 <= w5601 and not w22491;
w22493 <= w22488 and not w22492;
w22494 <= a(17) and not w22493;
w22495 <= not w22493 and not w22494;
w22496 <= a(17) and not w22494;
w22497 <= not w22495 and not w22496;
w22498 <= w4629 and w22309;
w22499 <= w4468 and w22315;
w22500 <= w4539 and w22312;
w22501 <= not w22499 and not w22500;
w22502 <= not w22498 and w22501;
w22503 <= w22371 and not w22373;
w22504 <= not w22374 and not w22503;
w22505 <= w4471 and w22504;
w22506 <= w22502 and not w22505;
w22507 <= a(23) and not w22506;
w22508 <= not w22506 and not w22507;
w22509 <= a(23) and not w22507;
w22510 <= not w22508 and not w22509;
w22511 <= w3819 and w22322;
w22512 <= w3902 and w22328;
w22513 <= w3981 and w22325;
w22514 <= not w22512 and not w22513;
w22515 <= not w22511 and w22514;
w22516 <= w22356 and not w22358;
w22517 <= not w22359 and not w22516;
w22518 <= w3985 and w22517;
w22519 <= w22515 and not w22518;
w22520 <= a(26) and not w22519;
w22521 <= not w22519 and not w22520;
w22522 <= a(26) and not w22520;
w22523 <= not w22521 and not w22522;
w22524 <= w3392 and w22331;
w22525 <= w3477 and w22337;
w22526 <= w3541 and w22334;
w22527 <= not w22525 and not w22526;
w22528 <= not w22524 and w22527;
w22529 <= w22344 and not w22346;
w22530 <= not w22347 and not w22529;
w22531 <= w3303 and w22530;
w22532 <= w22528 and not w22531;
w22533 <= a(29) and not w22532;
w22534 <= not w22532 and not w22533;
w22535 <= a(29) and not w22533;
w22536 <= not w22534 and not w22535;
w22537 <= not w3302 and not w22341;
w22538 <= a(29) and not w22537;
w22539 <= w3541 and not w22341;
w22540 <= w3392 and w22337;
w22541 <= not w22539 and not w22540;
w22542 <= w22337 and w22341;
w22543 <= not w22337 and not w22341;
w22544 <= not w22542 and not w22543;
w22545 <= w3303 and not w22544;
w22546 <= w22541 and not w22545;
w22547 <= a(29) and not w22546;
w22548 <= a(29) and not w22547;
w22549 <= not w22546 and not w22547;
w22550 <= not w22548 and not w22549;
w22551 <= w22538 and not w22550;
w22552 <= w3392 and w22334;
w22553 <= w3477 and not w22341;
w22554 <= w3541 and w22337;
w22555 <= not w22553 and not w22554;
w22556 <= not w22552 and w22555;
w22557 <= not w3303 and w22556;
w22558 <= not w22334 and w22542;
w22559 <= w22334 and not w22542;
w22560 <= not w22558 and not w22559;
w22561 <= w22556 and w22560;
w22562 <= not w22557 and not w22561;
w22563 <= a(29) and not w22562;
w22564 <= not a(29) and w22562;
w22565 <= not w22563 and not w22564;
w22566 <= w22551 and not w22565;
w22567 <= not w7414 and not w22341;
w22568 <= w22566 and not w22567;
w22569 <= not w22566 and w22567;
w22570 <= not w22568 and not w22569;
w22571 <= not w22536 and not w22570;
w22572 <= w22536 and w22570;
w22573 <= not w22571 and not w22572;
w22574 <= not w22523 and w22573;
w22575 <= not w22523 and not w22574;
w22576 <= w22573 and not w22574;
w22577 <= not w22575 and not w22576;
w22578 <= w3819 and w22325;
w22579 <= w3902 and w22331;
w22580 <= w3981 and w22328;
w22581 <= not w22579 and not w22580;
w22582 <= not w22578 and w22581;
w22583 <= w22352 and not w22354;
w22584 <= not w22355 and not w22583;
w22585 <= w3985 and w22584;
w22586 <= w22582 and not w22585;
w22587 <= a(26) and not w22586;
w22588 <= not w22586 and not w22587;
w22589 <= a(26) and not w22587;
w22590 <= not w22588 and not w22589;
w22591 <= not w22551 and w22565;
w22592 <= not w22566 and not w22591;
w22593 <= not w22590 and w22592;
w22594 <= not w22590 and not w22593;
w22595 <= w22592 and not w22593;
w22596 <= not w22594 and not w22595;
w22597 <= not w22538 and w22550;
w22598 <= not w22551 and not w22597;
w22599 <= w3819 and w22328;
w22600 <= w3902 and w22334;
w22601 <= w3981 and w22331;
w22602 <= not w22600 and not w22601;
w22603 <= not w22599 and w22602;
w22604 <= not w3985 and w22603;
w22605 <= w22348 and not w22350;
w22606 <= not w22351 and not w22605;
w22607 <= w22603 and not w22606;
w22608 <= not w22604 and not w22607;
w22609 <= a(26) and not w22608;
w22610 <= not a(26) and w22608;
w22611 <= not w22609 and not w22610;
w22612 <= w22598 and not w22611;
w22613 <= not w3815 and not w22341;
w22614 <= a(26) and not w22613;
w22615 <= w3981 and not w22341;
w22616 <= w3819 and w22337;
w22617 <= not w22615 and not w22616;
w22618 <= w3985 and not w22544;
w22619 <= w22617 and not w22618;
w22620 <= a(26) and not w22619;
w22621 <= a(26) and not w22620;
w22622 <= not w22619 and not w22620;
w22623 <= not w22621 and not w22622;
w22624 <= w22614 and not w22623;
w22625 <= w3819 and w22334;
w22626 <= w3902 and not w22341;
w22627 <= w3981 and w22337;
w22628 <= not w22626 and not w22627;
w22629 <= not w22625 and w22628;
w22630 <= not w3985 and w22629;
w22631 <= w22560 and w22629;
w22632 <= not w22630 and not w22631;
w22633 <= a(26) and not w22632;
w22634 <= not a(26) and w22632;
w22635 <= not w22633 and not w22634;
w22636 <= w22624 and not w22635;
w22637 <= w22537 and w22636;
w22638 <= w22636 and not w22637;
w22639 <= w22537 and not w22637;
w22640 <= not w22638 and not w22639;
w22641 <= w3819 and w22331;
w22642 <= w3902 and w22337;
w22643 <= w3981 and w22334;
w22644 <= not w22642 and not w22643;
w22645 <= not w22641 and w22644;
w22646 <= w3985 and w22530;
w22647 <= w22645 and not w22646;
w22648 <= a(26) and not w22647;
w22649 <= a(26) and not w22648;
w22650 <= not w22647 and not w22648;
w22651 <= not w22649 and not w22650;
w22652 <= not w22640 and not w22651;
w22653 <= not w22637 and not w22652;
w22654 <= not w22598 and w22611;
w22655 <= not w22612 and not w22654;
w22656 <= not w22653 and w22655;
w22657 <= not w22612 and not w22656;
w22658 <= not w22596 and not w22657;
w22659 <= not w22593 and not w22658;
w22660 <= not w22577 and not w22659;
w22661 <= not w22574 and not w22660;
w22662 <= w3392 and w22328;
w22663 <= w3477 and w22334;
w22664 <= w3541 and w22331;
w22665 <= not w22663 and not w22664;
w22666 <= not w22662 and w22665;
w22667 <= w3303 and w22606;
w22668 <= w22666 and not w22667;
w22669 <= a(29) and not w22668;
w22670 <= not w22668 and not w22669;
w22671 <= a(29) and not w22669;
w22672 <= not w22670 and not w22671;
w22673 <= w372 and w2026;
w22674 <= w820 and w22673;
w22675 <= w43 and w22674;
w22676 <= w1302 and w22675;
w22677 <= not w397 and w22676;
w22678 <= not w84 and w22677;
w22679 <= not w163 and w22678;
w22680 <= not w351 and w22679;
w22681 <= not w915 and w22680;
w22682 <= not w726 and w22681;
w22683 <= not w647 and w22682;
w22684 <= w3141 and w3793;
w22685 <= w2744 and w22684;
w22686 <= w4039 and w22685;
w22687 <= w14124 and w22686;
w22688 <= w739 and w22687;
w22689 <= w3098 and w22688;
w22690 <= w2211 and w22689;
w22691 <= w569 and w22690;
w22692 <= w353 and w22691;
w22693 <= w473 and w22692;
w22694 <= not w425 and w22693;
w22695 <= not w524 and w22694;
w22696 <= not w98 and w22695;
w22697 <= not w386 and w22696;
w22698 <= w670 and w2010;
w22699 <= w979 and w22698;
w22700 <= w15891 and w22699;
w22701 <= w22697 and w22700;
w22702 <= w22683 and w22701;
w22703 <= w15802 and w22702;
w22704 <= w1096 and w22703;
w22705 <= w1204 and w22704;
w22706 <= w1115 and w22705;
w22707 <= w745 and w22706;
w22708 <= w1063 and w22707;
w22709 <= w276 and w22708;
w22710 <= not w332 and w22709;
w22711 <= not w124 and w22710;
w22712 <= not w266 and w22711;
w22713 <= not w79 and w22712;
w22714 <= not w301 and w22713;
w22715 <= w2955 and w22337;
w22716 <= w10 and not w22544;
w22717 <= w2963 and not w22341;
w22718 <= not w22716 and not w22717;
w22719 <= not w22715 and w22718;
w22720 <= not w22714 and not w22719;
w22721 <= not w22714 and not w22720;
w22722 <= not w22719 and not w22720;
w22723 <= not w22721 and not w22722;
w22724 <= not w22672 and not w22723;
w22725 <= not w22672 and not w22724;
w22726 <= not w22723 and not w22724;
w22727 <= not w22725 and not w22726;
w22728 <= w22566 and w22567;
w22729 <= not w22571 and not w22728;
w22730 <= not w22727 and not w22729;
w22731 <= not w22727 and not w22730;
w22732 <= not w22729 and not w22730;
w22733 <= not w22731 and not w22732;
w22734 <= w3819 and w22319;
w22735 <= w3902 and w22325;
w22736 <= w3981 and w22322;
w22737 <= not w22735 and not w22736;
w22738 <= not w22734 and w22737;
w22739 <= not w3985 and w22738;
w22740 <= w22360 and not w22362;
w22741 <= not w22363 and not w22740;
w22742 <= w22738 and not w22741;
w22743 <= not w22739 and not w22742;
w22744 <= a(26) and not w22743;
w22745 <= not a(26) and w22743;
w22746 <= not w22744 and not w22745;
w22747 <= not w22733 and not w22746;
w22748 <= not w22733 and not w22747;
w22749 <= not w22746 and not w22747;
w22750 <= not w22748 and not w22749;
w22751 <= not w22661 and not w22750;
w22752 <= not w22661 and not w22751;
w22753 <= not w22750 and not w22751;
w22754 <= not w22752 and not w22753;
w22755 <= not w22510 and not w22754;
w22756 <= not w22510 and not w22755;
w22757 <= not w22754 and not w22755;
w22758 <= not w22756 and not w22757;
w22759 <= w22577 and w22659;
w22760 <= not w22660 and not w22759;
w22761 <= w4629 and w22312;
w22762 <= w4468 and w22319;
w22763 <= w4539 and w22315;
w22764 <= not w22762 and not w22763;
w22765 <= not w22761 and w22764;
w22766 <= not w4471 and w22765;
w22767 <= not w22368 and not w22370;
w22768 <= not w22317 and w22371;
w22769 <= not w22767 and not w22768;
w22770 <= w22765 and w22769;
w22771 <= not w22766 and not w22770;
w22772 <= a(23) and not w22771;
w22773 <= not a(23) and w22771;
w22774 <= not w22772 and not w22773;
w22775 <= w22760 and not w22774;
w22776 <= w22596 and w22657;
w22777 <= not w22658 and not w22776;
w22778 <= w4629 and w22315;
w22779 <= w4468 and w22322;
w22780 <= w4539 and w22319;
w22781 <= not w22779 and not w22780;
w22782 <= not w22778 and w22781;
w22783 <= not w4471 and w22782;
w22784 <= w22364 and not w22366;
w22785 <= not w22367 and not w22784;
w22786 <= w22782 and not w22785;
w22787 <= not w22783 and not w22786;
w22788 <= a(23) and not w22787;
w22789 <= not a(23) and w22787;
w22790 <= not w22788 and not w22789;
w22791 <= w22777 and not w22790;
w22792 <= w4629 and w22319;
w22793 <= w4468 and w22325;
w22794 <= w4539 and w22322;
w22795 <= not w22793 and not w22794;
w22796 <= not w22792 and w22795;
w22797 <= w4471 and w22741;
w22798 <= w22796 and not w22797;
w22799 <= a(23) and not w22798;
w22800 <= not w22798 and not w22799;
w22801 <= a(23) and not w22799;
w22802 <= not w22800 and not w22801;
w22803 <= w22653 and not w22655;
w22804 <= not w22656 and not w22803;
w22805 <= not w22802 and w22804;
w22806 <= not w22802 and not w22805;
w22807 <= w22804 and not w22805;
w22808 <= not w22806 and not w22807;
w22809 <= not w22640 and not w22652;
w22810 <= not w22651 and not w22652;
w22811 <= not w22809 and not w22810;
w22812 <= w4629 and w22322;
w22813 <= w4468 and w22328;
w22814 <= w4539 and w22325;
w22815 <= not w22813 and not w22814;
w22816 <= not w22812 and w22815;
w22817 <= not w4471 and w22816;
w22818 <= not w22517 and w22816;
w22819 <= not w22817 and not w22818;
w22820 <= a(23) and not w22819;
w22821 <= not a(23) and w22819;
w22822 <= not w22820 and not w22821;
w22823 <= not w22811 and not w22822;
w22824 <= w4629 and w22325;
w22825 <= w4468 and w22331;
w22826 <= w4539 and w22328;
w22827 <= not w22825 and not w22826;
w22828 <= not w22824 and w22827;
w22829 <= w4471 and w22584;
w22830 <= w22828 and not w22829;
w22831 <= a(23) and not w22830;
w22832 <= not w22830 and not w22831;
w22833 <= a(23) and not w22831;
w22834 <= not w22832 and not w22833;
w22835 <= not w22624 and w22635;
w22836 <= not w22636 and not w22835;
w22837 <= not w22834 and w22836;
w22838 <= not w22834 and not w22837;
w22839 <= w22836 and not w22837;
w22840 <= not w22838 and not w22839;
w22841 <= not w22614 and w22623;
w22842 <= not w22624 and not w22841;
w22843 <= w4629 and w22328;
w22844 <= w4468 and w22334;
w22845 <= w4539 and w22331;
w22846 <= not w22844 and not w22845;
w22847 <= not w22843 and w22846;
w22848 <= not w4471 and w22847;
w22849 <= not w22606 and w22847;
w22850 <= not w22848 and not w22849;
w22851 <= a(23) and not w22850;
w22852 <= not a(23) and w22850;
w22853 <= not w22851 and not w22852;
w22854 <= w22842 and not w22853;
w22855 <= not w4463 and not w22341;
w22856 <= a(23) and not w22855;
w22857 <= w4539 and not w22341;
w22858 <= w4629 and w22337;
w22859 <= not w22857 and not w22858;
w22860 <= w4471 and not w22544;
w22861 <= w22859 and not w22860;
w22862 <= a(23) and not w22861;
w22863 <= a(23) and not w22862;
w22864 <= not w22861 and not w22862;
w22865 <= not w22863 and not w22864;
w22866 <= w22856 and not w22865;
w22867 <= w4629 and w22334;
w22868 <= w4468 and not w22341;
w22869 <= w4539 and w22337;
w22870 <= not w22868 and not w22869;
w22871 <= not w22867 and w22870;
w22872 <= not w4471 and w22871;
w22873 <= w22560 and w22871;
w22874 <= not w22872 and not w22873;
w22875 <= a(23) and not w22874;
w22876 <= not a(23) and w22874;
w22877 <= not w22875 and not w22876;
w22878 <= w22866 and not w22877;
w22879 <= w22613 and w22878;
w22880 <= w22878 and not w22879;
w22881 <= w22613 and not w22879;
w22882 <= not w22880 and not w22881;
w22883 <= w4629 and w22331;
w22884 <= w4468 and w22337;
w22885 <= w4539 and w22334;
w22886 <= not w22884 and not w22885;
w22887 <= not w22883 and w22886;
w22888 <= w4471 and w22530;
w22889 <= w22887 and not w22888;
w22890 <= a(23) and not w22889;
w22891 <= a(23) and not w22890;
w22892 <= not w22889 and not w22890;
w22893 <= not w22891 and not w22892;
w22894 <= not w22882 and not w22893;
w22895 <= not w22879 and not w22894;
w22896 <= not w22842 and w22853;
w22897 <= not w22854 and not w22896;
w22898 <= not w22895 and w22897;
w22899 <= not w22854 and not w22898;
w22900 <= not w22840 and not w22899;
w22901 <= not w22837 and not w22900;
w22902 <= w22811 and w22822;
w22903 <= not w22823 and not w22902;
w22904 <= not w22901 and w22903;
w22905 <= not w22823 and not w22904;
w22906 <= not w22808 and not w22905;
w22907 <= not w22805 and not w22906;
w22908 <= w22777 and not w22791;
w22909 <= not w22790 and not w22791;
w22910 <= not w22908 and not w22909;
w22911 <= not w22907 and not w22910;
w22912 <= not w22791 and not w22911;
w22913 <= not w22760 and w22774;
w22914 <= not w22775 and not w22913;
w22915 <= not w22912 and w22914;
w22916 <= not w22775 and not w22915;
w22917 <= w22758 and w22916;
w22918 <= not w22758 and not w22916;
w22919 <= not w22917 and not w22918;
w22920 <= w5431 and w22300;
w22921 <= w4870 and w22306;
w22922 <= w5342 and w22303;
w22923 <= not w22921 and not w22922;
w22924 <= not w22920 and w22923;
w22925 <= not w4873 and w22924;
w22926 <= not w22383 and not w22386;
w22927 <= not w22384 and w22387;
w22928 <= not w22926 and not w22927;
w22929 <= w22924 and w22928;
w22930 <= not w22925 and not w22929;
w22931 <= a(20) and not w22930;
w22932 <= not a(20) and w22930;
w22933 <= not w22931 and not w22932;
w22934 <= w22919 and not w22933;
w22935 <= w5431 and w22303;
w22936 <= w4870 and w22309;
w22937 <= w5342 and w22306;
w22938 <= not w22936 and not w22937;
w22939 <= not w22935 and w22938;
w22940 <= w22379 and not w22381;
w22941 <= not w22382 and not w22940;
w22942 <= w4873 and w22941;
w22943 <= w22939 and not w22942;
w22944 <= a(20) and not w22943;
w22945 <= not w22943 and not w22944;
w22946 <= a(20) and not w22944;
w22947 <= not w22945 and not w22946;
w22948 <= w22912 and not w22914;
w22949 <= not w22915 and not w22948;
w22950 <= not w22947 and w22949;
w22951 <= not w22947 and not w22950;
w22952 <= w22949 and not w22950;
w22953 <= not w22951 and not w22952;
w22954 <= w5431 and w22306;
w22955 <= w4870 and w22312;
w22956 <= w5342 and w22309;
w22957 <= not w22955 and not w22956;
w22958 <= not w22954 and w22957;
w22959 <= w22375 and not w22377;
w22960 <= not w22378 and not w22959;
w22961 <= w4873 and w22960;
w22962 <= w22958 and not w22961;
w22963 <= a(20) and not w22962;
w22964 <= not w22962 and not w22963;
w22965 <= a(20) and not w22963;
w22966 <= not w22964 and not w22965;
w22967 <= not w22907 and not w22911;
w22968 <= not w22910 and not w22911;
w22969 <= not w22967 and not w22968;
w22970 <= not w22966 and not w22969;
w22971 <= not w22966 and not w22970;
w22972 <= not w22969 and not w22970;
w22973 <= not w22971 and not w22972;
w22974 <= w22808 and w22905;
w22975 <= not w22906 and not w22974;
w22976 <= w5431 and w22309;
w22977 <= w4870 and w22315;
w22978 <= w5342 and w22312;
w22979 <= not w22977 and not w22978;
w22980 <= not w22976 and w22979;
w22981 <= not w4873 and w22980;
w22982 <= not w22504 and w22980;
w22983 <= not w22981 and not w22982;
w22984 <= a(20) and not w22983;
w22985 <= not a(20) and w22983;
w22986 <= not w22984 and not w22985;
w22987 <= w22975 and not w22986;
w22988 <= w22901 and not w22903;
w22989 <= not w22904 and not w22988;
w22990 <= w5431 and w22312;
w22991 <= w4870 and w22319;
w22992 <= w5342 and w22315;
w22993 <= not w22991 and not w22992;
w22994 <= not w22990 and w22993;
w22995 <= not w4873 and w22994;
w22996 <= w22769 and w22994;
w22997 <= not w22995 and not w22996;
w22998 <= a(20) and not w22997;
w22999 <= not a(20) and w22997;
w23000 <= not w22998 and not w22999;
w23001 <= w22989 and not w23000;
w23002 <= w22840 and w22899;
w23003 <= not w22900 and not w23002;
w23004 <= w5431 and w22315;
w23005 <= w4870 and w22322;
w23006 <= w5342 and w22319;
w23007 <= not w23005 and not w23006;
w23008 <= not w23004 and w23007;
w23009 <= not w4873 and w23008;
w23010 <= not w22785 and w23008;
w23011 <= not w23009 and not w23010;
w23012 <= a(20) and not w23011;
w23013 <= not a(20) and w23011;
w23014 <= not w23012 and not w23013;
w23015 <= w23003 and not w23014;
w23016 <= w5431 and w22319;
w23017 <= w4870 and w22325;
w23018 <= w5342 and w22322;
w23019 <= not w23017 and not w23018;
w23020 <= not w23016 and w23019;
w23021 <= w4873 and w22741;
w23022 <= w23020 and not w23021;
w23023 <= a(20) and not w23022;
w23024 <= not w23022 and not w23023;
w23025 <= a(20) and not w23023;
w23026 <= not w23024 and not w23025;
w23027 <= w22895 and not w22897;
w23028 <= not w22898 and not w23027;
w23029 <= not w23026 and w23028;
w23030 <= not w23026 and not w23029;
w23031 <= w23028 and not w23029;
w23032 <= not w23030 and not w23031;
w23033 <= not w22882 and not w22894;
w23034 <= not w22893 and not w22894;
w23035 <= not w23033 and not w23034;
w23036 <= w5431 and w22322;
w23037 <= w4870 and w22328;
w23038 <= w5342 and w22325;
w23039 <= not w23037 and not w23038;
w23040 <= not w23036 and w23039;
w23041 <= not w4873 and w23040;
w23042 <= not w22517 and w23040;
w23043 <= not w23041 and not w23042;
w23044 <= a(20) and not w23043;
w23045 <= not a(20) and w23043;
w23046 <= not w23044 and not w23045;
w23047 <= not w23035 and not w23046;
w23048 <= w5431 and w22325;
w23049 <= w4870 and w22331;
w23050 <= w5342 and w22328;
w23051 <= not w23049 and not w23050;
w23052 <= not w23048 and w23051;
w23053 <= w4873 and w22584;
w23054 <= w23052 and not w23053;
w23055 <= a(20) and not w23054;
w23056 <= not w23054 and not w23055;
w23057 <= a(20) and not w23055;
w23058 <= not w23056 and not w23057;
w23059 <= not w22866 and w22877;
w23060 <= not w22878 and not w23059;
w23061 <= not w23058 and w23060;
w23062 <= not w23058 and not w23061;
w23063 <= w23060 and not w23061;
w23064 <= not w23062 and not w23063;
w23065 <= not w22856 and w22865;
w23066 <= not w22866 and not w23065;
w23067 <= w5431 and w22328;
w23068 <= w4870 and w22334;
w23069 <= w5342 and w22331;
w23070 <= not w23068 and not w23069;
w23071 <= not w23067 and w23070;
w23072 <= not w4873 and w23071;
w23073 <= not w22606 and w23071;
w23074 <= not w23072 and not w23073;
w23075 <= a(20) and not w23074;
w23076 <= not a(20) and w23074;
w23077 <= not w23075 and not w23076;
w23078 <= w23066 and not w23077;
w23079 <= w5342 and not w22341;
w23080 <= w5431 and w22337;
w23081 <= not w23079 and not w23080;
w23082 <= w4873 and not w22544;
w23083 <= w23081 and not w23082;
w23084 <= a(20) and not w23083;
w23085 <= a(20) and not w23084;
w23086 <= not w23083 and not w23084;
w23087 <= not w23085 and not w23086;
w23088 <= not w4868 and not w22341;
w23089 <= a(20) and not w23088;
w23090 <= not w23087 and w23089;
w23091 <= w5431 and w22334;
w23092 <= w4870 and not w22341;
w23093 <= w5342 and w22337;
w23094 <= not w23092 and not w23093;
w23095 <= not w23091 and w23094;
w23096 <= not w4873 and w23095;
w23097 <= w22560 and w23095;
w23098 <= not w23096 and not w23097;
w23099 <= a(20) and not w23098;
w23100 <= not a(20) and w23098;
w23101 <= not w23099 and not w23100;
w23102 <= w23090 and not w23101;
w23103 <= w22855 and w23102;
w23104 <= w23102 and not w23103;
w23105 <= w22855 and not w23103;
w23106 <= not w23104 and not w23105;
w23107 <= w5431 and w22331;
w23108 <= w4870 and w22337;
w23109 <= w5342 and w22334;
w23110 <= not w23108 and not w23109;
w23111 <= not w23107 and w23110;
w23112 <= w4873 and w22530;
w23113 <= w23111 and not w23112;
w23114 <= a(20) and not w23113;
w23115 <= a(20) and not w23114;
w23116 <= not w23113 and not w23114;
w23117 <= not w23115 and not w23116;
w23118 <= not w23106 and not w23117;
w23119 <= not w23103 and not w23118;
w23120 <= not w23066 and w23077;
w23121 <= not w23078 and not w23120;
w23122 <= not w23119 and w23121;
w23123 <= not w23078 and not w23122;
w23124 <= not w23064 and not w23123;
w23125 <= not w23061 and not w23124;
w23126 <= w23035 and w23046;
w23127 <= not w23047 and not w23126;
w23128 <= not w23125 and w23127;
w23129 <= not w23047 and not w23128;
w23130 <= not w23032 and not w23129;
w23131 <= not w23029 and not w23130;
w23132 <= w23003 and not w23015;
w23133 <= not w23014 and not w23015;
w23134 <= not w23132 and not w23133;
w23135 <= not w23131 and not w23134;
w23136 <= not w23015 and not w23135;
w23137 <= w22989 and not w23001;
w23138 <= not w23000 and not w23001;
w23139 <= not w23137 and not w23138;
w23140 <= not w23136 and not w23139;
w23141 <= not w23001 and not w23140;
w23142 <= not w22975 and w22986;
w23143 <= not w22987 and not w23142;
w23144 <= not w23141 and w23143;
w23145 <= not w22987 and not w23144;
w23146 <= not w22973 and not w23145;
w23147 <= not w22970 and not w23146;
w23148 <= not w22953 and not w23147;
w23149 <= not w22950 and not w23148;
w23150 <= w22919 and not w22934;
w23151 <= not w22933 and not w22934;
w23152 <= not w23150 and not w23151;
w23153 <= not w23149 and not w23152;
w23154 <= not w22934 and not w23153;
w23155 <= w4629 and w22306;
w23156 <= w4468 and w22312;
w23157 <= w4539 and w22309;
w23158 <= not w23156 and not w23157;
w23159 <= not w23155 and w23158;
w23160 <= w4471 and w22960;
w23161 <= w23159 and not w23160;
w23162 <= a(23) and not w23161;
w23163 <= not w23161 and not w23162;
w23164 <= a(23) and not w23162;
w23165 <= not w23163 and not w23164;
w23166 <= not w22747 and not w22751;
w23167 <= w3392 and w22325;
w23168 <= w3477 and w22331;
w23169 <= w3541 and w22328;
w23170 <= not w23168 and not w23169;
w23171 <= not w23167 and w23170;
w23172 <= w3303 and w22584;
w23173 <= w23171 and not w23172;
w23174 <= a(29) and not w23173;
w23175 <= not w23173 and not w23174;
w23176 <= a(29) and not w23174;
w23177 <= not w23175 and not w23176;
w23178 <= w10 and not w22560;
w23179 <= w2955 and w22334;
w23180 <= w2958 and not w22341;
w23181 <= w2963 and w22337;
w23182 <= not w23180 and not w23181;
w23183 <= not w23179 and w23182;
w23184 <= not w23178 and w23183;
w23185 <= not w168 and not w267;
w23186 <= not w21 and w23185;
w23187 <= w13709 and w23186;
w23188 <= w2976 and w23187;
w23189 <= w12322 and w23188;
w23190 <= w667 and w23189;
w23191 <= w3196 and w23190;
w23192 <= w6560 and w23191;
w23193 <= w5144 and w23192;
w23194 <= w902 and w23193;
w23195 <= w229 and w23194;
w23196 <= w1064 and w23195;
w23197 <= w666 and w23196;
w23198 <= w15802 and w23197;
w23199 <= not w355 and w23198;
w23200 <= not w215 and w23199;
w23201 <= not w163 and w23200;
w23202 <= not w915 and w23201;
w23203 <= not w608 and w23202;
w23204 <= not w502 and w23203;
w23205 <= w22720 and not w23204;
w23206 <= not w22720 and w23204;
w23207 <= not w23205 and not w23206;
w23208 <= not w23184 and w23207;
w23209 <= not w23184 and not w23208;
w23210 <= w23207 and not w23208;
w23211 <= not w23209 and not w23210;
w23212 <= not w23177 and not w23211;
w23213 <= not w23177 and not w23212;
w23214 <= not w23211 and not w23212;
w23215 <= not w23213 and not w23214;
w23216 <= not w22724 and not w22730;
w23217 <= w23215 and w23216;
w23218 <= not w23215 and not w23216;
w23219 <= not w23217 and not w23218;
w23220 <= w3819 and w22315;
w23221 <= w3902 and w22322;
w23222 <= w3981 and w22319;
w23223 <= not w23221 and not w23222;
w23224 <= not w23220 and w23223;
w23225 <= not w3985 and w23224;
w23226 <= not w22785 and w23224;
w23227 <= not w23225 and not w23226;
w23228 <= a(26) and not w23227;
w23229 <= not a(26) and w23227;
w23230 <= not w23228 and not w23229;
w23231 <= w23219 and not w23230;
w23232 <= w23219 and not w23231;
w23233 <= not w23230 and not w23231;
w23234 <= not w23232 and not w23233;
w23235 <= not w23166 and not w23234;
w23236 <= not w23166 and not w23235;
w23237 <= not w23234 and not w23235;
w23238 <= not w23236 and not w23237;
w23239 <= not w23165 and not w23238;
w23240 <= not w23165 and not w23239;
w23241 <= not w23238 and not w23239;
w23242 <= not w23240 and not w23241;
w23243 <= not w22755 and not w22918;
w23244 <= w23242 and w23243;
w23245 <= not w23242 and not w23243;
w23246 <= not w23244 and not w23245;
w23247 <= w5431 and w22297;
w23248 <= w4870 and w22303;
w23249 <= w5342 and w22300;
w23250 <= not w23248 and not w23249;
w23251 <= not w23247 and w23250;
w23252 <= not w4873 and w23251;
w23253 <= not w22387 and not w22390;
w23254 <= not w22388 and w22391;
w23255 <= not w23253 and not w23254;
w23256 <= w23251 and w23255;
w23257 <= not w23252 and not w23256;
w23258 <= a(20) and not w23257;
w23259 <= not a(20) and w23257;
w23260 <= not w23258 and not w23259;
w23261 <= w23246 and not w23260;
w23262 <= w23246 and not w23261;
w23263 <= not w23260 and not w23261;
w23264 <= not w23262 and not w23263;
w23265 <= not w23154 and not w23264;
w23266 <= not w23154 and not w23265;
w23267 <= not w23264 and not w23265;
w23268 <= not w23266 and not w23267;
w23269 <= not w22497 and not w23268;
w23270 <= not w22497 and not w23269;
w23271 <= not w23268 and not w23269;
w23272 <= not w23270 and not w23271;
w23273 <= w6168 and w22291;
w23274 <= w5598 and w22297;
w23275 <= w5874 and w22294;
w23276 <= not w23274 and not w23275;
w23277 <= not w23273 and w23276;
w23278 <= not w22395 and not w22398;
w23279 <= not w22396 and w22399;
w23280 <= not w23278 and not w23279;
w23281 <= w5601 and not w23280;
w23282 <= w23277 and not w23281;
w23283 <= a(17) and not w23282;
w23284 <= not w23282 and not w23283;
w23285 <= a(17) and not w23283;
w23286 <= not w23284 and not w23285;
w23287 <= not w23149 and not w23153;
w23288 <= not w23152 and not w23153;
w23289 <= not w23287 and not w23288;
w23290 <= not w23286 and not w23289;
w23291 <= not w23286 and not w23290;
w23292 <= not w23289 and not w23290;
w23293 <= not w23291 and not w23292;
w23294 <= w22953 and w23147;
w23295 <= not w23148 and not w23294;
w23296 <= w6168 and w22294;
w23297 <= w5598 and w22300;
w23298 <= w5874 and w22297;
w23299 <= not w23297 and not w23298;
w23300 <= not w23296 and w23299;
w23301 <= not w5601 and w23300;
w23302 <= w22391 and not w22393;
w23303 <= not w22394 and not w23302;
w23304 <= w23300 and not w23303;
w23305 <= not w23301 and not w23304;
w23306 <= a(17) and not w23305;
w23307 <= not a(17) and w23305;
w23308 <= not w23306 and not w23307;
w23309 <= w23295 and not w23308;
w23310 <= w22973 and w23145;
w23311 <= not w23146 and not w23310;
w23312 <= w6168 and w22297;
w23313 <= w5598 and w22303;
w23314 <= w5874 and w22300;
w23315 <= not w23313 and not w23314;
w23316 <= not w23312 and w23315;
w23317 <= not w5601 and w23316;
w23318 <= w23255 and w23316;
w23319 <= not w23317 and not w23318;
w23320 <= a(17) and not w23319;
w23321 <= not a(17) and w23319;
w23322 <= not w23320 and not w23321;
w23323 <= w23311 and not w23322;
w23324 <= w6168 and w22300;
w23325 <= w5598 and w22306;
w23326 <= w5874 and w22303;
w23327 <= not w23325 and not w23326;
w23328 <= not w23324 and w23327;
w23329 <= w5601 and not w22928;
w23330 <= w23328 and not w23329;
w23331 <= a(17) and not w23330;
w23332 <= not w23330 and not w23331;
w23333 <= a(17) and not w23331;
w23334 <= not w23332 and not w23333;
w23335 <= w23141 and not w23143;
w23336 <= not w23144 and not w23335;
w23337 <= not w23334 and w23336;
w23338 <= not w23334 and not w23337;
w23339 <= w23336 and not w23337;
w23340 <= not w23338 and not w23339;
w23341 <= w6168 and w22303;
w23342 <= w5598 and w22309;
w23343 <= w5874 and w22306;
w23344 <= not w23342 and not w23343;
w23345 <= not w23341 and w23344;
w23346 <= w5601 and w22941;
w23347 <= w23345 and not w23346;
w23348 <= a(17) and not w23347;
w23349 <= not w23347 and not w23348;
w23350 <= a(17) and not w23348;
w23351 <= not w23349 and not w23350;
w23352 <= not w23136 and not w23140;
w23353 <= not w23139 and not w23140;
w23354 <= not w23352 and not w23353;
w23355 <= not w23351 and not w23354;
w23356 <= not w23351 and not w23355;
w23357 <= not w23354 and not w23355;
w23358 <= not w23356 and not w23357;
w23359 <= w6168 and w22306;
w23360 <= w5598 and w22312;
w23361 <= w5874 and w22309;
w23362 <= not w23360 and not w23361;
w23363 <= not w23359 and w23362;
w23364 <= w5601 and w22960;
w23365 <= w23363 and not w23364;
w23366 <= a(17) and not w23365;
w23367 <= not w23365 and not w23366;
w23368 <= a(17) and not w23366;
w23369 <= not w23367 and not w23368;
w23370 <= not w23131 and not w23135;
w23371 <= not w23134 and not w23135;
w23372 <= not w23370 and not w23371;
w23373 <= not w23369 and not w23372;
w23374 <= not w23369 and not w23373;
w23375 <= not w23372 and not w23373;
w23376 <= not w23374 and not w23375;
w23377 <= w23032 and w23129;
w23378 <= not w23130 and not w23377;
w23379 <= w6168 and w22309;
w23380 <= w5598 and w22315;
w23381 <= w5874 and w22312;
w23382 <= not w23380 and not w23381;
w23383 <= not w23379 and w23382;
w23384 <= not w5601 and w23383;
w23385 <= not w22504 and w23383;
w23386 <= not w23384 and not w23385;
w23387 <= a(17) and not w23386;
w23388 <= not a(17) and w23386;
w23389 <= not w23387 and not w23388;
w23390 <= w23378 and not w23389;
w23391 <= w23125 and not w23127;
w23392 <= not w23128 and not w23391;
w23393 <= w6168 and w22312;
w23394 <= w5598 and w22319;
w23395 <= w5874 and w22315;
w23396 <= not w23394 and not w23395;
w23397 <= not w23393 and w23396;
w23398 <= not w5601 and w23397;
w23399 <= w22769 and w23397;
w23400 <= not w23398 and not w23399;
w23401 <= a(17) and not w23400;
w23402 <= not a(17) and w23400;
w23403 <= not w23401 and not w23402;
w23404 <= w23392 and not w23403;
w23405 <= w23064 and w23123;
w23406 <= not w23124 and not w23405;
w23407 <= w6168 and w22315;
w23408 <= w5598 and w22322;
w23409 <= w5874 and w22319;
w23410 <= not w23408 and not w23409;
w23411 <= not w23407 and w23410;
w23412 <= not w5601 and w23411;
w23413 <= not w22785 and w23411;
w23414 <= not w23412 and not w23413;
w23415 <= a(17) and not w23414;
w23416 <= not a(17) and w23414;
w23417 <= not w23415 and not w23416;
w23418 <= w23406 and not w23417;
w23419 <= w6168 and w22319;
w23420 <= w5598 and w22325;
w23421 <= w5874 and w22322;
w23422 <= not w23420 and not w23421;
w23423 <= not w23419 and w23422;
w23424 <= w5601 and w22741;
w23425 <= w23423 and not w23424;
w23426 <= a(17) and not w23425;
w23427 <= not w23425 and not w23426;
w23428 <= a(17) and not w23426;
w23429 <= not w23427 and not w23428;
w23430 <= w23119 and not w23121;
w23431 <= not w23122 and not w23430;
w23432 <= not w23429 and w23431;
w23433 <= not w23429 and not w23432;
w23434 <= w23431 and not w23432;
w23435 <= not w23433 and not w23434;
w23436 <= not w23106 and not w23118;
w23437 <= not w23117 and not w23118;
w23438 <= not w23436 and not w23437;
w23439 <= w6168 and w22322;
w23440 <= w5598 and w22328;
w23441 <= w5874 and w22325;
w23442 <= not w23440 and not w23441;
w23443 <= not w23439 and w23442;
w23444 <= not w5601 and w23443;
w23445 <= not w22517 and w23443;
w23446 <= not w23444 and not w23445;
w23447 <= a(17) and not w23446;
w23448 <= not a(17) and w23446;
w23449 <= not w23447 and not w23448;
w23450 <= not w23438 and not w23449;
w23451 <= w6168 and w22325;
w23452 <= w5598 and w22331;
w23453 <= w5874 and w22328;
w23454 <= not w23452 and not w23453;
w23455 <= not w23451 and w23454;
w23456 <= w5601 and w22584;
w23457 <= w23455 and not w23456;
w23458 <= a(17) and not w23457;
w23459 <= not w23457 and not w23458;
w23460 <= a(17) and not w23458;
w23461 <= not w23459 and not w23460;
w23462 <= not w23090 and w23101;
w23463 <= not w23102 and not w23462;
w23464 <= not w23461 and w23463;
w23465 <= not w23461 and not w23464;
w23466 <= w23463 and not w23464;
w23467 <= not w23465 and not w23466;
w23468 <= w23087 and not w23089;
w23469 <= not w23090 and not w23468;
w23470 <= w6168 and w22328;
w23471 <= w5598 and w22334;
w23472 <= w5874 and w22331;
w23473 <= not w23471 and not w23472;
w23474 <= not w23470 and w23473;
w23475 <= not w5601 and w23474;
w23476 <= not w22606 and w23474;
w23477 <= not w23475 and not w23476;
w23478 <= a(17) and not w23477;
w23479 <= not a(17) and w23477;
w23480 <= not w23478 and not w23479;
w23481 <= w23469 and not w23480;
w23482 <= w5874 and not w22341;
w23483 <= w6168 and w22337;
w23484 <= not w23482 and not w23483;
w23485 <= w5601 and not w22544;
w23486 <= w23484 and not w23485;
w23487 <= a(17) and not w23486;
w23488 <= a(17) and not w23487;
w23489 <= not w23486 and not w23487;
w23490 <= not w23488 and not w23489;
w23491 <= not w5593 and not w22341;
w23492 <= a(17) and not w23491;
w23493 <= not w23490 and w23492;
w23494 <= w6168 and w22334;
w23495 <= w5598 and not w22341;
w23496 <= w5874 and w22337;
w23497 <= not w23495 and not w23496;
w23498 <= not w23494 and w23497;
w23499 <= not w5601 and w23498;
w23500 <= w22560 and w23498;
w23501 <= not w23499 and not w23500;
w23502 <= a(17) and not w23501;
w23503 <= not a(17) and w23501;
w23504 <= not w23502 and not w23503;
w23505 <= w23493 and not w23504;
w23506 <= w23088 and w23505;
w23507 <= w23505 and not w23506;
w23508 <= w23088 and not w23506;
w23509 <= not w23507 and not w23508;
w23510 <= w6168 and w22331;
w23511 <= w5598 and w22337;
w23512 <= w5874 and w22334;
w23513 <= not w23511 and not w23512;
w23514 <= not w23510 and w23513;
w23515 <= w5601 and w22530;
w23516 <= w23514 and not w23515;
w23517 <= a(17) and not w23516;
w23518 <= a(17) and not w23517;
w23519 <= not w23516 and not w23517;
w23520 <= not w23518 and not w23519;
w23521 <= not w23509 and not w23520;
w23522 <= not w23506 and not w23521;
w23523 <= not w23469 and w23480;
w23524 <= not w23481 and not w23523;
w23525 <= not w23522 and w23524;
w23526 <= not w23481 and not w23525;
w23527 <= not w23467 and not w23526;
w23528 <= not w23464 and not w23527;
w23529 <= w23438 and w23449;
w23530 <= not w23450 and not w23529;
w23531 <= not w23528 and w23530;
w23532 <= not w23450 and not w23531;
w23533 <= not w23435 and not w23532;
w23534 <= not w23432 and not w23533;
w23535 <= w23406 and not w23418;
w23536 <= not w23417 and not w23418;
w23537 <= not w23535 and not w23536;
w23538 <= not w23534 and not w23537;
w23539 <= not w23418 and not w23538;
w23540 <= w23392 and not w23404;
w23541 <= not w23403 and not w23404;
w23542 <= not w23540 and not w23541;
w23543 <= not w23539 and not w23542;
w23544 <= not w23404 and not w23543;
w23545 <= not w23378 and w23389;
w23546 <= not w23390 and not w23545;
w23547 <= not w23544 and w23546;
w23548 <= not w23390 and not w23547;
w23549 <= not w23376 and not w23548;
w23550 <= not w23373 and not w23549;
w23551 <= not w23358 and not w23550;
w23552 <= not w23355 and not w23551;
w23553 <= not w23340 and not w23552;
w23554 <= not w23337 and not w23553;
w23555 <= w23311 and not w23323;
w23556 <= not w23322 and not w23323;
w23557 <= not w23555 and not w23556;
w23558 <= not w23554 and not w23557;
w23559 <= not w23323 and not w23558;
w23560 <= not w23295 and w23308;
w23561 <= not w23309 and not w23560;
w23562 <= not w23559 and w23561;
w23563 <= not w23309 and not w23562;
w23564 <= not w23293 and not w23563;
w23565 <= not w23290 and not w23564;
w23566 <= w23272 and w23565;
w23567 <= not w23272 and not w23565;
w23568 <= not w23566 and not w23567;
w23569 <= w7036 and w22279;
w23570 <= w6337 and w22285;
w23571 <= w6886 and w22282;
w23572 <= not w23570 and not w23571;
w23573 <= not w23569 and w23572;
w23574 <= not w6332 and w23573;
w23575 <= not w22411 and not w22414;
w23576 <= not w22412 and w22415;
w23577 <= not w23575 and not w23576;
w23578 <= w23573 and w23577;
w23579 <= not w23574 and not w23578;
w23580 <= a(14) and not w23579;
w23581 <= not a(14) and w23579;
w23582 <= not w23580 and not w23581;
w23583 <= w23568 and not w23582;
w23584 <= w23293 and w23563;
w23585 <= not w23564 and not w23584;
w23586 <= w7036 and w22282;
w23587 <= w6337 and w22288;
w23588 <= w6886 and w22285;
w23589 <= not w23587 and not w23588;
w23590 <= not w23586 and w23589;
w23591 <= not w6332 and w23590;
w23592 <= not w22407 and not w22410;
w23593 <= not w22408 and w22411;
w23594 <= not w23592 and not w23593;
w23595 <= w23590 and w23594;
w23596 <= not w23591 and not w23595;
w23597 <= a(14) and not w23596;
w23598 <= not a(14) and w23596;
w23599 <= not w23597 and not w23598;
w23600 <= w23585 and not w23599;
w23601 <= w7036 and w22285;
w23602 <= w6337 and w22291;
w23603 <= w6886 and w22288;
w23604 <= not w23602 and not w23603;
w23605 <= not w23601 and w23604;
w23606 <= w22403 and not w22405;
w23607 <= not w22406 and not w23606;
w23608 <= w6332 and w23607;
w23609 <= w23605 and not w23608;
w23610 <= a(14) and not w23609;
w23611 <= not w23609 and not w23610;
w23612 <= a(14) and not w23610;
w23613 <= not w23611 and not w23612;
w23614 <= w23559 and not w23561;
w23615 <= not w23562 and not w23614;
w23616 <= not w23613 and w23615;
w23617 <= not w23613 and not w23616;
w23618 <= w23615 and not w23616;
w23619 <= not w23617 and not w23618;
w23620 <= w7036 and w22288;
w23621 <= w6337 and w22294;
w23622 <= w6886 and w22291;
w23623 <= not w23621 and not w23622;
w23624 <= not w23620 and w23623;
w23625 <= w6332 and not w22491;
w23626 <= w23624 and not w23625;
w23627 <= a(14) and not w23626;
w23628 <= not w23626 and not w23627;
w23629 <= a(14) and not w23627;
w23630 <= not w23628 and not w23629;
w23631 <= not w23554 and not w23558;
w23632 <= not w23557 and not w23558;
w23633 <= not w23631 and not w23632;
w23634 <= not w23630 and not w23633;
w23635 <= not w23630 and not w23634;
w23636 <= not w23633 and not w23634;
w23637 <= not w23635 and not w23636;
w23638 <= w23340 and w23552;
w23639 <= not w23553 and not w23638;
w23640 <= w7036 and w22291;
w23641 <= w6337 and w22297;
w23642 <= w6886 and w22294;
w23643 <= not w23641 and not w23642;
w23644 <= not w23640 and w23643;
w23645 <= not w6332 and w23644;
w23646 <= w23280 and w23644;
w23647 <= not w23645 and not w23646;
w23648 <= a(14) and not w23647;
w23649 <= not a(14) and w23647;
w23650 <= not w23648 and not w23649;
w23651 <= w23639 and not w23650;
w23652 <= w23358 and w23550;
w23653 <= not w23551 and not w23652;
w23654 <= w7036 and w22294;
w23655 <= w6337 and w22300;
w23656 <= w6886 and w22297;
w23657 <= not w23655 and not w23656;
w23658 <= not w23654 and w23657;
w23659 <= not w6332 and w23658;
w23660 <= not w23303 and w23658;
w23661 <= not w23659 and not w23660;
w23662 <= a(14) and not w23661;
w23663 <= not a(14) and w23661;
w23664 <= not w23662 and not w23663;
w23665 <= w23653 and not w23664;
w23666 <= w23376 and w23548;
w23667 <= not w23549 and not w23666;
w23668 <= w7036 and w22297;
w23669 <= w6337 and w22303;
w23670 <= w6886 and w22300;
w23671 <= not w23669 and not w23670;
w23672 <= not w23668 and w23671;
w23673 <= not w6332 and w23672;
w23674 <= w23255 and w23672;
w23675 <= not w23673 and not w23674;
w23676 <= a(14) and not w23675;
w23677 <= not a(14) and w23675;
w23678 <= not w23676 and not w23677;
w23679 <= w23667 and not w23678;
w23680 <= w7036 and w22300;
w23681 <= w6337 and w22306;
w23682 <= w6886 and w22303;
w23683 <= not w23681 and not w23682;
w23684 <= not w23680 and w23683;
w23685 <= w6332 and not w22928;
w23686 <= w23684 and not w23685;
w23687 <= a(14) and not w23686;
w23688 <= not w23686 and not w23687;
w23689 <= a(14) and not w23687;
w23690 <= not w23688 and not w23689;
w23691 <= w23544 and not w23546;
w23692 <= not w23547 and not w23691;
w23693 <= not w23690 and w23692;
w23694 <= not w23690 and not w23693;
w23695 <= w23692 and not w23693;
w23696 <= not w23694 and not w23695;
w23697 <= w7036 and w22303;
w23698 <= w6337 and w22309;
w23699 <= w6886 and w22306;
w23700 <= not w23698 and not w23699;
w23701 <= not w23697 and w23700;
w23702 <= w6332 and w22941;
w23703 <= w23701 and not w23702;
w23704 <= a(14) and not w23703;
w23705 <= not w23703 and not w23704;
w23706 <= a(14) and not w23704;
w23707 <= not w23705 and not w23706;
w23708 <= not w23539 and not w23543;
w23709 <= not w23542 and not w23543;
w23710 <= not w23708 and not w23709;
w23711 <= not w23707 and not w23710;
w23712 <= not w23707 and not w23711;
w23713 <= not w23710 and not w23711;
w23714 <= not w23712 and not w23713;
w23715 <= w7036 and w22306;
w23716 <= w6337 and w22312;
w23717 <= w6886 and w22309;
w23718 <= not w23716 and not w23717;
w23719 <= not w23715 and w23718;
w23720 <= w6332 and w22960;
w23721 <= w23719 and not w23720;
w23722 <= a(14) and not w23721;
w23723 <= not w23721 and not w23722;
w23724 <= a(14) and not w23722;
w23725 <= not w23723 and not w23724;
w23726 <= not w23534 and not w23538;
w23727 <= not w23537 and not w23538;
w23728 <= not w23726 and not w23727;
w23729 <= not w23725 and not w23728;
w23730 <= not w23725 and not w23729;
w23731 <= not w23728 and not w23729;
w23732 <= not w23730 and not w23731;
w23733 <= w23435 and w23532;
w23734 <= not w23533 and not w23733;
w23735 <= w7036 and w22309;
w23736 <= w6337 and w22315;
w23737 <= w6886 and w22312;
w23738 <= not w23736 and not w23737;
w23739 <= not w23735 and w23738;
w23740 <= not w6332 and w23739;
w23741 <= not w22504 and w23739;
w23742 <= not w23740 and not w23741;
w23743 <= a(14) and not w23742;
w23744 <= not a(14) and w23742;
w23745 <= not w23743 and not w23744;
w23746 <= w23734 and not w23745;
w23747 <= w23528 and not w23530;
w23748 <= not w23531 and not w23747;
w23749 <= w7036 and w22312;
w23750 <= w6337 and w22319;
w23751 <= w6886 and w22315;
w23752 <= not w23750 and not w23751;
w23753 <= not w23749 and w23752;
w23754 <= not w6332 and w23753;
w23755 <= w22769 and w23753;
w23756 <= not w23754 and not w23755;
w23757 <= a(14) and not w23756;
w23758 <= not a(14) and w23756;
w23759 <= not w23757 and not w23758;
w23760 <= w23748 and not w23759;
w23761 <= w23467 and w23526;
w23762 <= not w23527 and not w23761;
w23763 <= w7036 and w22315;
w23764 <= w6337 and w22322;
w23765 <= w6886 and w22319;
w23766 <= not w23764 and not w23765;
w23767 <= not w23763 and w23766;
w23768 <= not w6332 and w23767;
w23769 <= not w22785 and w23767;
w23770 <= not w23768 and not w23769;
w23771 <= a(14) and not w23770;
w23772 <= not a(14) and w23770;
w23773 <= not w23771 and not w23772;
w23774 <= w23762 and not w23773;
w23775 <= w7036 and w22319;
w23776 <= w6337 and w22325;
w23777 <= w6886 and w22322;
w23778 <= not w23776 and not w23777;
w23779 <= not w23775 and w23778;
w23780 <= w6332 and w22741;
w23781 <= w23779 and not w23780;
w23782 <= a(14) and not w23781;
w23783 <= not w23781 and not w23782;
w23784 <= a(14) and not w23782;
w23785 <= not w23783 and not w23784;
w23786 <= w23522 and not w23524;
w23787 <= not w23525 and not w23786;
w23788 <= not w23785 and w23787;
w23789 <= not w23785 and not w23788;
w23790 <= w23787 and not w23788;
w23791 <= not w23789 and not w23790;
w23792 <= not w23509 and not w23521;
w23793 <= not w23520 and not w23521;
w23794 <= not w23792 and not w23793;
w23795 <= w7036 and w22322;
w23796 <= w6337 and w22328;
w23797 <= w6886 and w22325;
w23798 <= not w23796 and not w23797;
w23799 <= not w23795 and w23798;
w23800 <= not w6332 and w23799;
w23801 <= not w22517 and w23799;
w23802 <= not w23800 and not w23801;
w23803 <= a(14) and not w23802;
w23804 <= not a(14) and w23802;
w23805 <= not w23803 and not w23804;
w23806 <= not w23794 and not w23805;
w23807 <= w7036 and w22325;
w23808 <= w6337 and w22331;
w23809 <= w6886 and w22328;
w23810 <= not w23808 and not w23809;
w23811 <= not w23807 and w23810;
w23812 <= w6332 and w22584;
w23813 <= w23811 and not w23812;
w23814 <= a(14) and not w23813;
w23815 <= not w23813 and not w23814;
w23816 <= a(14) and not w23814;
w23817 <= not w23815 and not w23816;
w23818 <= not w23493 and w23504;
w23819 <= not w23505 and not w23818;
w23820 <= not w23817 and w23819;
w23821 <= not w23817 and not w23820;
w23822 <= w23819 and not w23820;
w23823 <= not w23821 and not w23822;
w23824 <= w23490 and not w23492;
w23825 <= not w23493 and not w23824;
w23826 <= w7036 and w22328;
w23827 <= w6337 and w22334;
w23828 <= w6886 and w22331;
w23829 <= not w23827 and not w23828;
w23830 <= not w23826 and w23829;
w23831 <= not w6332 and w23830;
w23832 <= not w22606 and w23830;
w23833 <= not w23831 and not w23832;
w23834 <= a(14) and not w23833;
w23835 <= not a(14) and w23833;
w23836 <= not w23834 and not w23835;
w23837 <= w23825 and not w23836;
w23838 <= w6886 and not w22341;
w23839 <= w7036 and w22337;
w23840 <= not w23838 and not w23839;
w23841 <= w6332 and not w22544;
w23842 <= w23840 and not w23841;
w23843 <= a(14) and not w23842;
w23844 <= a(14) and not w23843;
w23845 <= not w23842 and not w23843;
w23846 <= not w23844 and not w23845;
w23847 <= not w6328 and not w22341;
w23848 <= a(14) and not w23847;
w23849 <= not w23846 and w23848;
w23850 <= w7036 and w22334;
w23851 <= w6337 and not w22341;
w23852 <= w6886 and w22337;
w23853 <= not w23851 and not w23852;
w23854 <= not w23850 and w23853;
w23855 <= not w6332 and w23854;
w23856 <= w22560 and w23854;
w23857 <= not w23855 and not w23856;
w23858 <= a(14) and not w23857;
w23859 <= not a(14) and w23857;
w23860 <= not w23858 and not w23859;
w23861 <= w23849 and not w23860;
w23862 <= w23491 and w23861;
w23863 <= w23861 and not w23862;
w23864 <= w23491 and not w23862;
w23865 <= not w23863 and not w23864;
w23866 <= w7036 and w22331;
w23867 <= w6337 and w22337;
w23868 <= w6886 and w22334;
w23869 <= not w23867 and not w23868;
w23870 <= not w23866 and w23869;
w23871 <= w6332 and w22530;
w23872 <= w23870 and not w23871;
w23873 <= a(14) and not w23872;
w23874 <= a(14) and not w23873;
w23875 <= not w23872 and not w23873;
w23876 <= not w23874 and not w23875;
w23877 <= not w23865 and not w23876;
w23878 <= not w23862 and not w23877;
w23879 <= not w23825 and w23836;
w23880 <= not w23837 and not w23879;
w23881 <= not w23878 and w23880;
w23882 <= not w23837 and not w23881;
w23883 <= not w23823 and not w23882;
w23884 <= not w23820 and not w23883;
w23885 <= w23794 and w23805;
w23886 <= not w23806 and not w23885;
w23887 <= not w23884 and w23886;
w23888 <= not w23806 and not w23887;
w23889 <= not w23791 and not w23888;
w23890 <= not w23788 and not w23889;
w23891 <= w23762 and not w23774;
w23892 <= not w23773 and not w23774;
w23893 <= not w23891 and not w23892;
w23894 <= not w23890 and not w23893;
w23895 <= not w23774 and not w23894;
w23896 <= w23748 and not w23760;
w23897 <= not w23759 and not w23760;
w23898 <= not w23896 and not w23897;
w23899 <= not w23895 and not w23898;
w23900 <= not w23760 and not w23899;
w23901 <= not w23734 and w23745;
w23902 <= not w23746 and not w23901;
w23903 <= not w23900 and w23902;
w23904 <= not w23746 and not w23903;
w23905 <= not w23732 and not w23904;
w23906 <= not w23729 and not w23905;
w23907 <= not w23714 and not w23906;
w23908 <= not w23711 and not w23907;
w23909 <= not w23696 and not w23908;
w23910 <= not w23693 and not w23909;
w23911 <= w23667 and not w23679;
w23912 <= not w23678 and not w23679;
w23913 <= not w23911 and not w23912;
w23914 <= not w23910 and not w23913;
w23915 <= not w23679 and not w23914;
w23916 <= w23653 and not w23665;
w23917 <= not w23664 and not w23665;
w23918 <= not w23916 and not w23917;
w23919 <= not w23915 and not w23918;
w23920 <= not w23665 and not w23919;
w23921 <= not w23639 and w23650;
w23922 <= not w23651 and not w23921;
w23923 <= not w23920 and w23922;
w23924 <= not w23651 and not w23923;
w23925 <= not w23637 and not w23924;
w23926 <= not w23634 and not w23925;
w23927 <= not w23619 and not w23926;
w23928 <= not w23616 and not w23927;
w23929 <= w23585 and not w23600;
w23930 <= not w23599 and not w23600;
w23931 <= not w23929 and not w23930;
w23932 <= not w23928 and not w23931;
w23933 <= not w23600 and not w23932;
w23934 <= w23568 and not w23583;
w23935 <= not w23582 and not w23583;
w23936 <= not w23934 and not w23935;
w23937 <= not w23933 and not w23936;
w23938 <= not w23583 and not w23937;
w23939 <= w6168 and w22285;
w23940 <= w5598 and w22291;
w23941 <= w5874 and w22288;
w23942 <= not w23940 and not w23941;
w23943 <= not w23939 and w23942;
w23944 <= w5601 and w23607;
w23945 <= w23943 and not w23944;
w23946 <= a(17) and not w23945;
w23947 <= not w23945 and not w23946;
w23948 <= a(17) and not w23946;
w23949 <= not w23947 and not w23948;
w23950 <= not w23261 and not w23265;
w23951 <= w4629 and w22303;
w23952 <= w4468 and w22309;
w23953 <= w4539 and w22306;
w23954 <= not w23952 and not w23953;
w23955 <= not w23951 and w23954;
w23956 <= w4471 and w22941;
w23957 <= w23955 and not w23956;
w23958 <= a(23) and not w23957;
w23959 <= not w23957 and not w23958;
w23960 <= a(23) and not w23958;
w23961 <= not w23959 and not w23960;
w23962 <= not w23231 and not w23235;
w23963 <= w3392 and w22322;
w23964 <= w3477 and w22328;
w23965 <= w3541 and w22325;
w23966 <= not w23964 and not w23965;
w23967 <= not w23963 and w23966;
w23968 <= w3303 and w22517;
w23969 <= w23967 and not w23968;
w23970 <= a(29) and not w23969;
w23971 <= not w23969 and not w23970;
w23972 <= a(29) and not w23970;
w23973 <= not w23971 and not w23972;
w23974 <= not w23205 and not w23208;
w23975 <= w51 and not w446;
w23976 <= not w449 and w23975;
w23977 <= w1906 and w4937;
w23978 <= w23976 and w23977;
w23979 <= w4151 and w23978;
w23980 <= w1556 and w23979;
w23981 <= w5231 and w23980;
w23982 <= w851 and w23981;
w23983 <= w3225 and w23982;
w23984 <= w2281 and w23983;
w23985 <= w226 and w23984;
w23986 <= w406 and w23985;
w23987 <= w1466 and w23986;
w23988 <= w455 and w23987;
w23989 <= not w53 and w23988;
w23990 <= not w37 and w23989;
w23991 <= not w726 and w23990;
w23992 <= not w160 and w23991;
w23993 <= w2955 and w22331;
w23994 <= w2963 and w22334;
w23995 <= w2958 and w22337;
w23996 <= w10 and w22530;
w23997 <= not w23995 and not w23996;
w23998 <= not w23994 and w23997;
w23999 <= not w23993 and w23998;
w24000 <= not w23992 and not w23999;
w24001 <= not w23992 and not w24000;
w24002 <= not w23999 and not w24000;
w24003 <= not w24001 and not w24002;
w24004 <= not w23974 and not w24003;
w24005 <= not w23974 and not w24004;
w24006 <= not w24003 and not w24004;
w24007 <= not w24005 and not w24006;
w24008 <= not w23973 and not w24007;
w24009 <= not w23973 and not w24008;
w24010 <= not w24007 and not w24008;
w24011 <= not w24009 and not w24010;
w24012 <= not w23212 and not w23218;
w24013 <= w24011 and w24012;
w24014 <= not w24011 and not w24012;
w24015 <= not w24013 and not w24014;
w24016 <= w3819 and w22312;
w24017 <= w3902 and w22319;
w24018 <= w3981 and w22315;
w24019 <= not w24017 and not w24018;
w24020 <= not w24016 and w24019;
w24021 <= not w3985 and w24020;
w24022 <= w22769 and w24020;
w24023 <= not w24021 and not w24022;
w24024 <= a(26) and not w24023;
w24025 <= not a(26) and w24023;
w24026 <= not w24024 and not w24025;
w24027 <= w24015 and not w24026;
w24028 <= w24015 and not w24027;
w24029 <= not w24026 and not w24027;
w24030 <= not w24028 and not w24029;
w24031 <= not w23962 and not w24030;
w24032 <= not w23962 and not w24031;
w24033 <= not w24030 and not w24031;
w24034 <= not w24032 and not w24033;
w24035 <= not w23961 and not w24034;
w24036 <= not w23961 and not w24035;
w24037 <= not w24034 and not w24035;
w24038 <= not w24036 and not w24037;
w24039 <= not w23239 and not w23245;
w24040 <= w24038 and w24039;
w24041 <= not w24038 and not w24039;
w24042 <= not w24040 and not w24041;
w24043 <= w5431 and w22294;
w24044 <= w4870 and w22300;
w24045 <= w5342 and w22297;
w24046 <= not w24044 and not w24045;
w24047 <= not w24043 and w24046;
w24048 <= not w4873 and w24047;
w24049 <= not w23303 and w24047;
w24050 <= not w24048 and not w24049;
w24051 <= a(20) and not w24050;
w24052 <= not a(20) and w24050;
w24053 <= not w24051 and not w24052;
w24054 <= w24042 and not w24053;
w24055 <= w24042 and not w24054;
w24056 <= not w24053 and not w24054;
w24057 <= not w24055 and not w24056;
w24058 <= not w23950 and not w24057;
w24059 <= not w23950 and not w24058;
w24060 <= not w24057 and not w24058;
w24061 <= not w24059 and not w24060;
w24062 <= not w23949 and not w24061;
w24063 <= not w23949 and not w24062;
w24064 <= not w24061 and not w24062;
w24065 <= not w24063 and not w24064;
w24066 <= not w23269 and not w23567;
w24067 <= w24065 and w24066;
w24068 <= not w24065 and not w24066;
w24069 <= not w24067 and not w24068;
w24070 <= w7036 and w22276;
w24071 <= w6337 and w22282;
w24072 <= w6886 and w22279;
w24073 <= not w24071 and not w24072;
w24074 <= not w24070 and w24073;
w24075 <= not w6332 and w24074;
w24076 <= w22415 and not w22417;
w24077 <= not w22418 and not w24076;
w24078 <= w24074 and not w24077;
w24079 <= not w24075 and not w24078;
w24080 <= a(14) and not w24079;
w24081 <= not a(14) and w24079;
w24082 <= not w24080 and not w24081;
w24083 <= w24069 and not w24082;
w24084 <= w24069 and not w24083;
w24085 <= not w24082 and not w24083;
w24086 <= not w24084 and not w24085;
w24087 <= not w23938 and not w24086;
w24088 <= not w23938 and not w24087;
w24089 <= not w24086 and not w24087;
w24090 <= not w24088 and not w24089;
w24091 <= not w22483 and not w24090;
w24092 <= not w22483 and not w24091;
w24093 <= not w24090 and not w24091;
w24094 <= not w24092 and not w24093;
w24095 <= w7918 and w22270;
w24096 <= w7226 and w22276;
w24097 <= w7567 and w22273;
w24098 <= not w24096 and not w24097;
w24099 <= not w24095 and w24098;
w24100 <= not w22423 and not w22426;
w24101 <= not w22424 and w22427;
w24102 <= not w24100 and not w24101;
w24103 <= w7229 and not w24102;
w24104 <= w24099 and not w24103;
w24105 <= a(11) and not w24104;
w24106 <= not w24104 and not w24105;
w24107 <= a(11) and not w24105;
w24108 <= not w24106 and not w24107;
w24109 <= not w23933 and not w23937;
w24110 <= not w23936 and not w23937;
w24111 <= not w24109 and not w24110;
w24112 <= not w24108 and not w24111;
w24113 <= not w24108 and not w24112;
w24114 <= not w24111 and not w24112;
w24115 <= not w24113 and not w24114;
w24116 <= w7918 and w22273;
w24117 <= w7226 and w22279;
w24118 <= w7567 and w22276;
w24119 <= not w24117 and not w24118;
w24120 <= not w24116 and w24119;
w24121 <= not w22419 and not w22422;
w24122 <= not w22420 and w22423;
w24123 <= not w24121 and not w24122;
w24124 <= w7229 and not w24123;
w24125 <= w24120 and not w24124;
w24126 <= a(11) and not w24125;
w24127 <= not w24125 and not w24126;
w24128 <= a(11) and not w24126;
w24129 <= not w24127 and not w24128;
w24130 <= not w23928 and not w23932;
w24131 <= not w23931 and not w23932;
w24132 <= not w24130 and not w24131;
w24133 <= not w24129 and not w24132;
w24134 <= not w24129 and not w24133;
w24135 <= not w24132 and not w24133;
w24136 <= not w24134 and not w24135;
w24137 <= w23619 and w23926;
w24138 <= not w23927 and not w24137;
w24139 <= w7918 and w22276;
w24140 <= w7226 and w22282;
w24141 <= w7567 and w22279;
w24142 <= not w24140 and not w24141;
w24143 <= not w24139 and w24142;
w24144 <= not w7229 and w24143;
w24145 <= not w24077 and w24143;
w24146 <= not w24144 and not w24145;
w24147 <= a(11) and not w24146;
w24148 <= not a(11) and w24146;
w24149 <= not w24147 and not w24148;
w24150 <= w24138 and not w24149;
w24151 <= w23637 and w23924;
w24152 <= not w23925 and not w24151;
w24153 <= w7918 and w22279;
w24154 <= w7226 and w22285;
w24155 <= w7567 and w22282;
w24156 <= not w24154 and not w24155;
w24157 <= not w24153 and w24156;
w24158 <= not w7229 and w24157;
w24159 <= w23577 and w24157;
w24160 <= not w24158 and not w24159;
w24161 <= a(11) and not w24160;
w24162 <= not a(11) and w24160;
w24163 <= not w24161 and not w24162;
w24164 <= w24152 and not w24163;
w24165 <= w7918 and w22282;
w24166 <= w7226 and w22288;
w24167 <= w7567 and w22285;
w24168 <= not w24166 and not w24167;
w24169 <= not w24165 and w24168;
w24170 <= w7229 and not w23594;
w24171 <= w24169 and not w24170;
w24172 <= a(11) and not w24171;
w24173 <= not w24171 and not w24172;
w24174 <= a(11) and not w24172;
w24175 <= not w24173 and not w24174;
w24176 <= w23920 and not w23922;
w24177 <= not w23923 and not w24176;
w24178 <= not w24175 and w24177;
w24179 <= not w24175 and not w24178;
w24180 <= w24177 and not w24178;
w24181 <= not w24179 and not w24180;
w24182 <= w7918 and w22285;
w24183 <= w7226 and w22291;
w24184 <= w7567 and w22288;
w24185 <= not w24183 and not w24184;
w24186 <= not w24182 and w24185;
w24187 <= w7229 and w23607;
w24188 <= w24186 and not w24187;
w24189 <= a(11) and not w24188;
w24190 <= not w24188 and not w24189;
w24191 <= a(11) and not w24189;
w24192 <= not w24190 and not w24191;
w24193 <= not w23915 and not w23919;
w24194 <= not w23918 and not w23919;
w24195 <= not w24193 and not w24194;
w24196 <= not w24192 and not w24195;
w24197 <= not w24192 and not w24196;
w24198 <= not w24195 and not w24196;
w24199 <= not w24197 and not w24198;
w24200 <= w7918 and w22288;
w24201 <= w7226 and w22294;
w24202 <= w7567 and w22291;
w24203 <= not w24201 and not w24202;
w24204 <= not w24200 and w24203;
w24205 <= w7229 and not w22491;
w24206 <= w24204 and not w24205;
w24207 <= a(11) and not w24206;
w24208 <= not w24206 and not w24207;
w24209 <= a(11) and not w24207;
w24210 <= not w24208 and not w24209;
w24211 <= not w23910 and not w23914;
w24212 <= not w23913 and not w23914;
w24213 <= not w24211 and not w24212;
w24214 <= not w24210 and not w24213;
w24215 <= not w24210 and not w24214;
w24216 <= not w24213 and not w24214;
w24217 <= not w24215 and not w24216;
w24218 <= w23696 and w23908;
w24219 <= not w23909 and not w24218;
w24220 <= w7918 and w22291;
w24221 <= w7226 and w22297;
w24222 <= w7567 and w22294;
w24223 <= not w24221 and not w24222;
w24224 <= not w24220 and w24223;
w24225 <= not w7229 and w24224;
w24226 <= w23280 and w24224;
w24227 <= not w24225 and not w24226;
w24228 <= a(11) and not w24227;
w24229 <= not a(11) and w24227;
w24230 <= not w24228 and not w24229;
w24231 <= w24219 and not w24230;
w24232 <= w23714 and w23906;
w24233 <= not w23907 and not w24232;
w24234 <= w7918 and w22294;
w24235 <= w7226 and w22300;
w24236 <= w7567 and w22297;
w24237 <= not w24235 and not w24236;
w24238 <= not w24234 and w24237;
w24239 <= not w7229 and w24238;
w24240 <= not w23303 and w24238;
w24241 <= not w24239 and not w24240;
w24242 <= a(11) and not w24241;
w24243 <= not a(11) and w24241;
w24244 <= not w24242 and not w24243;
w24245 <= w24233 and not w24244;
w24246 <= w23732 and w23904;
w24247 <= not w23905 and not w24246;
w24248 <= w7918 and w22297;
w24249 <= w7226 and w22303;
w24250 <= w7567 and w22300;
w24251 <= not w24249 and not w24250;
w24252 <= not w24248 and w24251;
w24253 <= not w7229 and w24252;
w24254 <= w23255 and w24252;
w24255 <= not w24253 and not w24254;
w24256 <= a(11) and not w24255;
w24257 <= not a(11) and w24255;
w24258 <= not w24256 and not w24257;
w24259 <= w24247 and not w24258;
w24260 <= w7918 and w22300;
w24261 <= w7226 and w22306;
w24262 <= w7567 and w22303;
w24263 <= not w24261 and not w24262;
w24264 <= not w24260 and w24263;
w24265 <= w7229 and not w22928;
w24266 <= w24264 and not w24265;
w24267 <= a(11) and not w24266;
w24268 <= not w24266 and not w24267;
w24269 <= a(11) and not w24267;
w24270 <= not w24268 and not w24269;
w24271 <= w23900 and not w23902;
w24272 <= not w23903 and not w24271;
w24273 <= not w24270 and w24272;
w24274 <= not w24270 and not w24273;
w24275 <= w24272 and not w24273;
w24276 <= not w24274 and not w24275;
w24277 <= w7918 and w22303;
w24278 <= w7226 and w22309;
w24279 <= w7567 and w22306;
w24280 <= not w24278 and not w24279;
w24281 <= not w24277 and w24280;
w24282 <= w7229 and w22941;
w24283 <= w24281 and not w24282;
w24284 <= a(11) and not w24283;
w24285 <= not w24283 and not w24284;
w24286 <= a(11) and not w24284;
w24287 <= not w24285 and not w24286;
w24288 <= not w23895 and not w23899;
w24289 <= not w23898 and not w23899;
w24290 <= not w24288 and not w24289;
w24291 <= not w24287 and not w24290;
w24292 <= not w24287 and not w24291;
w24293 <= not w24290 and not w24291;
w24294 <= not w24292 and not w24293;
w24295 <= w7918 and w22306;
w24296 <= w7226 and w22312;
w24297 <= w7567 and w22309;
w24298 <= not w24296 and not w24297;
w24299 <= not w24295 and w24298;
w24300 <= w7229 and w22960;
w24301 <= w24299 and not w24300;
w24302 <= a(11) and not w24301;
w24303 <= not w24301 and not w24302;
w24304 <= a(11) and not w24302;
w24305 <= not w24303 and not w24304;
w24306 <= not w23890 and not w23894;
w24307 <= not w23893 and not w23894;
w24308 <= not w24306 and not w24307;
w24309 <= not w24305 and not w24308;
w24310 <= not w24305 and not w24309;
w24311 <= not w24308 and not w24309;
w24312 <= not w24310 and not w24311;
w24313 <= w23791 and w23888;
w24314 <= not w23889 and not w24313;
w24315 <= w7918 and w22309;
w24316 <= w7226 and w22315;
w24317 <= w7567 and w22312;
w24318 <= not w24316 and not w24317;
w24319 <= not w24315 and w24318;
w24320 <= not w7229 and w24319;
w24321 <= not w22504 and w24319;
w24322 <= not w24320 and not w24321;
w24323 <= a(11) and not w24322;
w24324 <= not a(11) and w24322;
w24325 <= not w24323 and not w24324;
w24326 <= w24314 and not w24325;
w24327 <= w23884 and not w23886;
w24328 <= not w23887 and not w24327;
w24329 <= w7918 and w22312;
w24330 <= w7226 and w22319;
w24331 <= w7567 and w22315;
w24332 <= not w24330 and not w24331;
w24333 <= not w24329 and w24332;
w24334 <= not w7229 and w24333;
w24335 <= w22769 and w24333;
w24336 <= not w24334 and not w24335;
w24337 <= a(11) and not w24336;
w24338 <= not a(11) and w24336;
w24339 <= not w24337 and not w24338;
w24340 <= w24328 and not w24339;
w24341 <= w23823 and w23882;
w24342 <= not w23883 and not w24341;
w24343 <= w7918 and w22315;
w24344 <= w7226 and w22322;
w24345 <= w7567 and w22319;
w24346 <= not w24344 and not w24345;
w24347 <= not w24343 and w24346;
w24348 <= not w7229 and w24347;
w24349 <= not w22785 and w24347;
w24350 <= not w24348 and not w24349;
w24351 <= a(11) and not w24350;
w24352 <= not a(11) and w24350;
w24353 <= not w24351 and not w24352;
w24354 <= w24342 and not w24353;
w24355 <= w7918 and w22319;
w24356 <= w7226 and w22325;
w24357 <= w7567 and w22322;
w24358 <= not w24356 and not w24357;
w24359 <= not w24355 and w24358;
w24360 <= w7229 and w22741;
w24361 <= w24359 and not w24360;
w24362 <= a(11) and not w24361;
w24363 <= not w24361 and not w24362;
w24364 <= a(11) and not w24362;
w24365 <= not w24363 and not w24364;
w24366 <= w23878 and not w23880;
w24367 <= not w23881 and not w24366;
w24368 <= not w24365 and w24367;
w24369 <= not w24365 and not w24368;
w24370 <= w24367 and not w24368;
w24371 <= not w24369 and not w24370;
w24372 <= not w23865 and not w23877;
w24373 <= not w23876 and not w23877;
w24374 <= not w24372 and not w24373;
w24375 <= w7918 and w22322;
w24376 <= w7226 and w22328;
w24377 <= w7567 and w22325;
w24378 <= not w24376 and not w24377;
w24379 <= not w24375 and w24378;
w24380 <= not w7229 and w24379;
w24381 <= not w22517 and w24379;
w24382 <= not w24380 and not w24381;
w24383 <= a(11) and not w24382;
w24384 <= not a(11) and w24382;
w24385 <= not w24383 and not w24384;
w24386 <= not w24374 and not w24385;
w24387 <= w7918 and w22325;
w24388 <= w7226 and w22331;
w24389 <= w7567 and w22328;
w24390 <= not w24388 and not w24389;
w24391 <= not w24387 and w24390;
w24392 <= w7229 and w22584;
w24393 <= w24391 and not w24392;
w24394 <= a(11) and not w24393;
w24395 <= not w24393 and not w24394;
w24396 <= a(11) and not w24394;
w24397 <= not w24395 and not w24396;
w24398 <= not w23849 and w23860;
w24399 <= not w23861 and not w24398;
w24400 <= not w24397 and w24399;
w24401 <= not w24397 and not w24400;
w24402 <= w24399 and not w24400;
w24403 <= not w24401 and not w24402;
w24404 <= w23846 and not w23848;
w24405 <= not w23849 and not w24404;
w24406 <= w7918 and w22328;
w24407 <= w7226 and w22334;
w24408 <= w7567 and w22331;
w24409 <= not w24407 and not w24408;
w24410 <= not w24406 and w24409;
w24411 <= not w7229 and w24410;
w24412 <= not w22606 and w24410;
w24413 <= not w24411 and not w24412;
w24414 <= a(11) and not w24413;
w24415 <= not a(11) and w24413;
w24416 <= not w24414 and not w24415;
w24417 <= w24405 and not w24416;
w24418 <= w7567 and not w22341;
w24419 <= w7918 and w22337;
w24420 <= not w24418 and not w24419;
w24421 <= w7229 and not w22544;
w24422 <= w24420 and not w24421;
w24423 <= a(11) and not w24422;
w24424 <= a(11) and not w24423;
w24425 <= not w24422 and not w24423;
w24426 <= not w24424 and not w24425;
w24427 <= not w7224 and not w22341;
w24428 <= a(11) and not w24427;
w24429 <= not w24426 and w24428;
w24430 <= w7918 and w22334;
w24431 <= w7226 and not w22341;
w24432 <= w7567 and w22337;
w24433 <= not w24431 and not w24432;
w24434 <= not w24430 and w24433;
w24435 <= not w7229 and w24434;
w24436 <= w22560 and w24434;
w24437 <= not w24435 and not w24436;
w24438 <= a(11) and not w24437;
w24439 <= not a(11) and w24437;
w24440 <= not w24438 and not w24439;
w24441 <= w24429 and not w24440;
w24442 <= w23847 and w24441;
w24443 <= w24441 and not w24442;
w24444 <= w23847 and not w24442;
w24445 <= not w24443 and not w24444;
w24446 <= w7918 and w22331;
w24447 <= w7226 and w22337;
w24448 <= w7567 and w22334;
w24449 <= not w24447 and not w24448;
w24450 <= not w24446 and w24449;
w24451 <= w7229 and w22530;
w24452 <= w24450 and not w24451;
w24453 <= a(11) and not w24452;
w24454 <= a(11) and not w24453;
w24455 <= not w24452 and not w24453;
w24456 <= not w24454 and not w24455;
w24457 <= not w24445 and not w24456;
w24458 <= not w24442 and not w24457;
w24459 <= not w24405 and w24416;
w24460 <= not w24417 and not w24459;
w24461 <= not w24458 and w24460;
w24462 <= not w24417 and not w24461;
w24463 <= not w24403 and not w24462;
w24464 <= not w24400 and not w24463;
w24465 <= w24374 and w24385;
w24466 <= not w24386 and not w24465;
w24467 <= not w24464 and w24466;
w24468 <= not w24386 and not w24467;
w24469 <= not w24371 and not w24468;
w24470 <= not w24368 and not w24469;
w24471 <= w24342 and not w24354;
w24472 <= not w24353 and not w24354;
w24473 <= not w24471 and not w24472;
w24474 <= not w24470 and not w24473;
w24475 <= not w24354 and not w24474;
w24476 <= w24328 and not w24340;
w24477 <= not w24339 and not w24340;
w24478 <= not w24476 and not w24477;
w24479 <= not w24475 and not w24478;
w24480 <= not w24340 and not w24479;
w24481 <= not w24314 and w24325;
w24482 <= not w24326 and not w24481;
w24483 <= not w24480 and w24482;
w24484 <= not w24326 and not w24483;
w24485 <= not w24312 and not w24484;
w24486 <= not w24309 and not w24485;
w24487 <= not w24294 and not w24486;
w24488 <= not w24291 and not w24487;
w24489 <= not w24276 and not w24488;
w24490 <= not w24273 and not w24489;
w24491 <= w24247 and not w24259;
w24492 <= not w24258 and not w24259;
w24493 <= not w24491 and not w24492;
w24494 <= not w24490 and not w24493;
w24495 <= not w24259 and not w24494;
w24496 <= w24233 and not w24245;
w24497 <= not w24244 and not w24245;
w24498 <= not w24496 and not w24497;
w24499 <= not w24495 and not w24498;
w24500 <= not w24245 and not w24499;
w24501 <= not w24219 and w24230;
w24502 <= not w24231 and not w24501;
w24503 <= not w24500 and w24502;
w24504 <= not w24231 and not w24503;
w24505 <= not w24217 and not w24504;
w24506 <= not w24214 and not w24505;
w24507 <= not w24199 and not w24506;
w24508 <= not w24196 and not w24507;
w24509 <= not w24181 and not w24508;
w24510 <= not w24178 and not w24509;
w24511 <= w24152 and not w24164;
w24512 <= not w24163 and not w24164;
w24513 <= not w24511 and not w24512;
w24514 <= not w24510 and not w24513;
w24515 <= not w24164 and not w24514;
w24516 <= not w24138 and w24149;
w24517 <= not w24150 and not w24516;
w24518 <= not w24515 and w24517;
w24519 <= not w24150 and not w24518;
w24520 <= not w24136 and not w24519;
w24521 <= not w24133 and not w24520;
w24522 <= not w24115 and not w24521;
w24523 <= not w24112 and not w24522;
w24524 <= w24094 and w24523;
w24525 <= not w24094 and not w24523;
w24526 <= not w24524 and not w24525;
w24527 <= w9266 and w22258;
w24528 <= w8353 and w22264;
w24529 <= w8795 and w22261;
w24530 <= not w24528 and not w24529;
w24531 <= not w24527 and w24530;
w24532 <= not w8356 and w24531;
w24533 <= w22439 and not w22441;
w24534 <= not w22442 and not w24533;
w24535 <= w24531 and not w24534;
w24536 <= not w24532 and not w24535;
w24537 <= a(8) and not w24536;
w24538 <= not a(8) and w24536;
w24539 <= not w24537 and not w24538;
w24540 <= w24526 and not w24539;
w24541 <= w24115 and w24521;
w24542 <= not w24522 and not w24541;
w24543 <= w9266 and w22261;
w24544 <= w8353 and w22267;
w24545 <= w8795 and w22264;
w24546 <= not w24544 and not w24545;
w24547 <= not w24543 and w24546;
w24548 <= not w8356 and w24547;
w24549 <= not w22435 and not w22438;
w24550 <= not w22436 and w22439;
w24551 <= not w24549 and not w24550;
w24552 <= w24547 and w24551;
w24553 <= not w24548 and not w24552;
w24554 <= a(8) and not w24553;
w24555 <= not a(8) and w24553;
w24556 <= not w24554 and not w24555;
w24557 <= w24542 and not w24556;
w24558 <= w24136 and w24519;
w24559 <= not w24520 and not w24558;
w24560 <= w9266 and w22264;
w24561 <= w8353 and w22270;
w24562 <= w8795 and w22267;
w24563 <= not w24561 and not w24562;
w24564 <= not w24560 and w24563;
w24565 <= not w8356 and w24564;
w24566 <= not w22431 and not w22434;
w24567 <= not w22432 and w22435;
w24568 <= not w24566 and not w24567;
w24569 <= w24564 and w24568;
w24570 <= not w24565 and not w24569;
w24571 <= a(8) and not w24570;
w24572 <= not a(8) and w24570;
w24573 <= not w24571 and not w24572;
w24574 <= w24559 and not w24573;
w24575 <= w9266 and w22267;
w24576 <= w8353 and w22273;
w24577 <= w8795 and w22270;
w24578 <= not w24576 and not w24577;
w24579 <= not w24575 and w24578;
w24580 <= w8356 and w22477;
w24581 <= w24579 and not w24580;
w24582 <= a(8) and not w24581;
w24583 <= not w24581 and not w24582;
w24584 <= a(8) and not w24582;
w24585 <= not w24583 and not w24584;
w24586 <= w24515 and not w24517;
w24587 <= not w24518 and not w24586;
w24588 <= not w24585 and w24587;
w24589 <= not w24585 and not w24588;
w24590 <= w24587 and not w24588;
w24591 <= not w24589 and not w24590;
w24592 <= w9266 and w22270;
w24593 <= w8353 and w22276;
w24594 <= w8795 and w22273;
w24595 <= not w24593 and not w24594;
w24596 <= not w24592 and w24595;
w24597 <= w8356 and not w24102;
w24598 <= w24596 and not w24597;
w24599 <= a(8) and not w24598;
w24600 <= not w24598 and not w24599;
w24601 <= a(8) and not w24599;
w24602 <= not w24600 and not w24601;
w24603 <= not w24510 and not w24514;
w24604 <= not w24513 and not w24514;
w24605 <= not w24603 and not w24604;
w24606 <= not w24602 and not w24605;
w24607 <= not w24602 and not w24606;
w24608 <= not w24605 and not w24606;
w24609 <= not w24607 and not w24608;
w24610 <= w24181 and w24508;
w24611 <= not w24509 and not w24610;
w24612 <= w9266 and w22273;
w24613 <= w8353 and w22279;
w24614 <= w8795 and w22276;
w24615 <= not w24613 and not w24614;
w24616 <= not w24612 and w24615;
w24617 <= not w8356 and w24616;
w24618 <= w24123 and w24616;
w24619 <= not w24617 and not w24618;
w24620 <= a(8) and not w24619;
w24621 <= not a(8) and w24619;
w24622 <= not w24620 and not w24621;
w24623 <= w24611 and not w24622;
w24624 <= w24199 and w24506;
w24625 <= not w24507 and not w24624;
w24626 <= w9266 and w22276;
w24627 <= w8353 and w22282;
w24628 <= w8795 and w22279;
w24629 <= not w24627 and not w24628;
w24630 <= not w24626 and w24629;
w24631 <= not w8356 and w24630;
w24632 <= not w24077 and w24630;
w24633 <= not w24631 and not w24632;
w24634 <= a(8) and not w24633;
w24635 <= not a(8) and w24633;
w24636 <= not w24634 and not w24635;
w24637 <= w24625 and not w24636;
w24638 <= w24217 and w24504;
w24639 <= not w24505 and not w24638;
w24640 <= w9266 and w22279;
w24641 <= w8353 and w22285;
w24642 <= w8795 and w22282;
w24643 <= not w24641 and not w24642;
w24644 <= not w24640 and w24643;
w24645 <= not w8356 and w24644;
w24646 <= w23577 and w24644;
w24647 <= not w24645 and not w24646;
w24648 <= a(8) and not w24647;
w24649 <= not a(8) and w24647;
w24650 <= not w24648 and not w24649;
w24651 <= w24639 and not w24650;
w24652 <= w9266 and w22282;
w24653 <= w8353 and w22288;
w24654 <= w8795 and w22285;
w24655 <= not w24653 and not w24654;
w24656 <= not w24652 and w24655;
w24657 <= w8356 and not w23594;
w24658 <= w24656 and not w24657;
w24659 <= a(8) and not w24658;
w24660 <= not w24658 and not w24659;
w24661 <= a(8) and not w24659;
w24662 <= not w24660 and not w24661;
w24663 <= w24500 and not w24502;
w24664 <= not w24503 and not w24663;
w24665 <= not w24662 and w24664;
w24666 <= not w24662 and not w24665;
w24667 <= w24664 and not w24665;
w24668 <= not w24666 and not w24667;
w24669 <= w9266 and w22285;
w24670 <= w8353 and w22291;
w24671 <= w8795 and w22288;
w24672 <= not w24670 and not w24671;
w24673 <= not w24669 and w24672;
w24674 <= w8356 and w23607;
w24675 <= w24673 and not w24674;
w24676 <= a(8) and not w24675;
w24677 <= not w24675 and not w24676;
w24678 <= a(8) and not w24676;
w24679 <= not w24677 and not w24678;
w24680 <= not w24495 and not w24499;
w24681 <= not w24498 and not w24499;
w24682 <= not w24680 and not w24681;
w24683 <= not w24679 and not w24682;
w24684 <= not w24679 and not w24683;
w24685 <= not w24682 and not w24683;
w24686 <= not w24684 and not w24685;
w24687 <= w9266 and w22288;
w24688 <= w8353 and w22294;
w24689 <= w8795 and w22291;
w24690 <= not w24688 and not w24689;
w24691 <= not w24687 and w24690;
w24692 <= w8356 and not w22491;
w24693 <= w24691 and not w24692;
w24694 <= a(8) and not w24693;
w24695 <= not w24693 and not w24694;
w24696 <= a(8) and not w24694;
w24697 <= not w24695 and not w24696;
w24698 <= not w24490 and not w24494;
w24699 <= not w24493 and not w24494;
w24700 <= not w24698 and not w24699;
w24701 <= not w24697 and not w24700;
w24702 <= not w24697 and not w24701;
w24703 <= not w24700 and not w24701;
w24704 <= not w24702 and not w24703;
w24705 <= w24276 and w24488;
w24706 <= not w24489 and not w24705;
w24707 <= w9266 and w22291;
w24708 <= w8353 and w22297;
w24709 <= w8795 and w22294;
w24710 <= not w24708 and not w24709;
w24711 <= not w24707 and w24710;
w24712 <= not w8356 and w24711;
w24713 <= w23280 and w24711;
w24714 <= not w24712 and not w24713;
w24715 <= a(8) and not w24714;
w24716 <= not a(8) and w24714;
w24717 <= not w24715 and not w24716;
w24718 <= w24706 and not w24717;
w24719 <= w24294 and w24486;
w24720 <= not w24487 and not w24719;
w24721 <= w9266 and w22294;
w24722 <= w8353 and w22300;
w24723 <= w8795 and w22297;
w24724 <= not w24722 and not w24723;
w24725 <= not w24721 and w24724;
w24726 <= not w8356 and w24725;
w24727 <= not w23303 and w24725;
w24728 <= not w24726 and not w24727;
w24729 <= a(8) and not w24728;
w24730 <= not a(8) and w24728;
w24731 <= not w24729 and not w24730;
w24732 <= w24720 and not w24731;
w24733 <= w24312 and w24484;
w24734 <= not w24485 and not w24733;
w24735 <= w9266 and w22297;
w24736 <= w8353 and w22303;
w24737 <= w8795 and w22300;
w24738 <= not w24736 and not w24737;
w24739 <= not w24735 and w24738;
w24740 <= not w8356 and w24739;
w24741 <= w23255 and w24739;
w24742 <= not w24740 and not w24741;
w24743 <= a(8) and not w24742;
w24744 <= not a(8) and w24742;
w24745 <= not w24743 and not w24744;
w24746 <= w24734 and not w24745;
w24747 <= w9266 and w22300;
w24748 <= w8353 and w22306;
w24749 <= w8795 and w22303;
w24750 <= not w24748 and not w24749;
w24751 <= not w24747 and w24750;
w24752 <= w8356 and not w22928;
w24753 <= w24751 and not w24752;
w24754 <= a(8) and not w24753;
w24755 <= not w24753 and not w24754;
w24756 <= a(8) and not w24754;
w24757 <= not w24755 and not w24756;
w24758 <= w24480 and not w24482;
w24759 <= not w24483 and not w24758;
w24760 <= not w24757 and w24759;
w24761 <= not w24757 and not w24760;
w24762 <= w24759 and not w24760;
w24763 <= not w24761 and not w24762;
w24764 <= w9266 and w22303;
w24765 <= w8353 and w22309;
w24766 <= w8795 and w22306;
w24767 <= not w24765 and not w24766;
w24768 <= not w24764 and w24767;
w24769 <= w8356 and w22941;
w24770 <= w24768 and not w24769;
w24771 <= a(8) and not w24770;
w24772 <= not w24770 and not w24771;
w24773 <= a(8) and not w24771;
w24774 <= not w24772 and not w24773;
w24775 <= not w24475 and not w24479;
w24776 <= not w24478 and not w24479;
w24777 <= not w24775 and not w24776;
w24778 <= not w24774 and not w24777;
w24779 <= not w24774 and not w24778;
w24780 <= not w24777 and not w24778;
w24781 <= not w24779 and not w24780;
w24782 <= w9266 and w22306;
w24783 <= w8353 and w22312;
w24784 <= w8795 and w22309;
w24785 <= not w24783 and not w24784;
w24786 <= not w24782 and w24785;
w24787 <= w8356 and w22960;
w24788 <= w24786 and not w24787;
w24789 <= a(8) and not w24788;
w24790 <= not w24788 and not w24789;
w24791 <= a(8) and not w24789;
w24792 <= not w24790 and not w24791;
w24793 <= not w24470 and not w24474;
w24794 <= not w24473 and not w24474;
w24795 <= not w24793 and not w24794;
w24796 <= not w24792 and not w24795;
w24797 <= not w24792 and not w24796;
w24798 <= not w24795 and not w24796;
w24799 <= not w24797 and not w24798;
w24800 <= w24371 and w24468;
w24801 <= not w24469 and not w24800;
w24802 <= w9266 and w22309;
w24803 <= w8353 and w22315;
w24804 <= w8795 and w22312;
w24805 <= not w24803 and not w24804;
w24806 <= not w24802 and w24805;
w24807 <= not w8356 and w24806;
w24808 <= not w22504 and w24806;
w24809 <= not w24807 and not w24808;
w24810 <= a(8) and not w24809;
w24811 <= not a(8) and w24809;
w24812 <= not w24810 and not w24811;
w24813 <= w24801 and not w24812;
w24814 <= w24464 and not w24466;
w24815 <= not w24467 and not w24814;
w24816 <= w9266 and w22312;
w24817 <= w8353 and w22319;
w24818 <= w8795 and w22315;
w24819 <= not w24817 and not w24818;
w24820 <= not w24816 and w24819;
w24821 <= not w8356 and w24820;
w24822 <= w22769 and w24820;
w24823 <= not w24821 and not w24822;
w24824 <= a(8) and not w24823;
w24825 <= not a(8) and w24823;
w24826 <= not w24824 and not w24825;
w24827 <= w24815 and not w24826;
w24828 <= w24403 and w24462;
w24829 <= not w24463 and not w24828;
w24830 <= w9266 and w22315;
w24831 <= w8353 and w22322;
w24832 <= w8795 and w22319;
w24833 <= not w24831 and not w24832;
w24834 <= not w24830 and w24833;
w24835 <= not w8356 and w24834;
w24836 <= not w22785 and w24834;
w24837 <= not w24835 and not w24836;
w24838 <= a(8) and not w24837;
w24839 <= not a(8) and w24837;
w24840 <= not w24838 and not w24839;
w24841 <= w24829 and not w24840;
w24842 <= w9266 and w22319;
w24843 <= w8353 and w22325;
w24844 <= w8795 and w22322;
w24845 <= not w24843 and not w24844;
w24846 <= not w24842 and w24845;
w24847 <= w8356 and w22741;
w24848 <= w24846 and not w24847;
w24849 <= a(8) and not w24848;
w24850 <= not w24848 and not w24849;
w24851 <= a(8) and not w24849;
w24852 <= not w24850 and not w24851;
w24853 <= w24458 and not w24460;
w24854 <= not w24461 and not w24853;
w24855 <= not w24852 and w24854;
w24856 <= not w24852 and not w24855;
w24857 <= w24854 and not w24855;
w24858 <= not w24856 and not w24857;
w24859 <= not w24445 and not w24457;
w24860 <= not w24456 and not w24457;
w24861 <= not w24859 and not w24860;
w24862 <= w9266 and w22322;
w24863 <= w8353 and w22328;
w24864 <= w8795 and w22325;
w24865 <= not w24863 and not w24864;
w24866 <= not w24862 and w24865;
w24867 <= not w8356 and w24866;
w24868 <= not w22517 and w24866;
w24869 <= not w24867 and not w24868;
w24870 <= a(8) and not w24869;
w24871 <= not a(8) and w24869;
w24872 <= not w24870 and not w24871;
w24873 <= not w24861 and not w24872;
w24874 <= w9266 and w22325;
w24875 <= w8353 and w22331;
w24876 <= w8795 and w22328;
w24877 <= not w24875 and not w24876;
w24878 <= not w24874 and w24877;
w24879 <= w8356 and w22584;
w24880 <= w24878 and not w24879;
w24881 <= a(8) and not w24880;
w24882 <= not w24880 and not w24881;
w24883 <= a(8) and not w24881;
w24884 <= not w24882 and not w24883;
w24885 <= not w24429 and w24440;
w24886 <= not w24441 and not w24885;
w24887 <= not w24884 and w24886;
w24888 <= not w24884 and not w24887;
w24889 <= w24886 and not w24887;
w24890 <= not w24888 and not w24889;
w24891 <= w24426 and not w24428;
w24892 <= not w24429 and not w24891;
w24893 <= w9266 and w22328;
w24894 <= w8353 and w22334;
w24895 <= w8795 and w22331;
w24896 <= not w24894 and not w24895;
w24897 <= not w24893 and w24896;
w24898 <= not w8356 and w24897;
w24899 <= not w22606 and w24897;
w24900 <= not w24898 and not w24899;
w24901 <= a(8) and not w24900;
w24902 <= not a(8) and w24900;
w24903 <= not w24901 and not w24902;
w24904 <= w24892 and not w24903;
w24905 <= w8795 and not w22341;
w24906 <= w9266 and w22337;
w24907 <= not w24905 and not w24906;
w24908 <= w8356 and not w22544;
w24909 <= w24907 and not w24908;
w24910 <= a(8) and not w24909;
w24911 <= a(8) and not w24910;
w24912 <= not w24909 and not w24910;
w24913 <= not w24911 and not w24912;
w24914 <= not w8351 and not w22341;
w24915 <= a(8) and not w24914;
w24916 <= not w24913 and w24915;
w24917 <= w9266 and w22334;
w24918 <= w8353 and not w22341;
w24919 <= w8795 and w22337;
w24920 <= not w24918 and not w24919;
w24921 <= not w24917 and w24920;
w24922 <= not w8356 and w24921;
w24923 <= w22560 and w24921;
w24924 <= not w24922 and not w24923;
w24925 <= a(8) and not w24924;
w24926 <= not a(8) and w24924;
w24927 <= not w24925 and not w24926;
w24928 <= w24916 and not w24927;
w24929 <= w24427 and w24928;
w24930 <= w24928 and not w24929;
w24931 <= w24427 and not w24929;
w24932 <= not w24930 and not w24931;
w24933 <= w9266 and w22331;
w24934 <= w8353 and w22337;
w24935 <= w8795 and w22334;
w24936 <= not w24934 and not w24935;
w24937 <= not w24933 and w24936;
w24938 <= w8356 and w22530;
w24939 <= w24937 and not w24938;
w24940 <= a(8) and not w24939;
w24941 <= a(8) and not w24940;
w24942 <= not w24939 and not w24940;
w24943 <= not w24941 and not w24942;
w24944 <= not w24932 and not w24943;
w24945 <= not w24929 and not w24944;
w24946 <= not w24892 and w24903;
w24947 <= not w24904 and not w24946;
w24948 <= not w24945 and w24947;
w24949 <= not w24904 and not w24948;
w24950 <= not w24890 and not w24949;
w24951 <= not w24887 and not w24950;
w24952 <= w24861 and w24872;
w24953 <= not w24873 and not w24952;
w24954 <= not w24951 and w24953;
w24955 <= not w24873 and not w24954;
w24956 <= not w24858 and not w24955;
w24957 <= not w24855 and not w24956;
w24958 <= w24829 and not w24841;
w24959 <= not w24840 and not w24841;
w24960 <= not w24958 and not w24959;
w24961 <= not w24957 and not w24960;
w24962 <= not w24841 and not w24961;
w24963 <= w24815 and not w24827;
w24964 <= not w24826 and not w24827;
w24965 <= not w24963 and not w24964;
w24966 <= not w24962 and not w24965;
w24967 <= not w24827 and not w24966;
w24968 <= not w24801 and w24812;
w24969 <= not w24813 and not w24968;
w24970 <= not w24967 and w24969;
w24971 <= not w24813 and not w24970;
w24972 <= not w24799 and not w24971;
w24973 <= not w24796 and not w24972;
w24974 <= not w24781 and not w24973;
w24975 <= not w24778 and not w24974;
w24976 <= not w24763 and not w24975;
w24977 <= not w24760 and not w24976;
w24978 <= w24734 and not w24746;
w24979 <= not w24745 and not w24746;
w24980 <= not w24978 and not w24979;
w24981 <= not w24977 and not w24980;
w24982 <= not w24746 and not w24981;
w24983 <= w24720 and not w24732;
w24984 <= not w24731 and not w24732;
w24985 <= not w24983 and not w24984;
w24986 <= not w24982 and not w24985;
w24987 <= not w24732 and not w24986;
w24988 <= not w24706 and w24717;
w24989 <= not w24718 and not w24988;
w24990 <= not w24987 and w24989;
w24991 <= not w24718 and not w24990;
w24992 <= not w24704 and not w24991;
w24993 <= not w24701 and not w24992;
w24994 <= not w24686 and not w24993;
w24995 <= not w24683 and not w24994;
w24996 <= not w24668 and not w24995;
w24997 <= not w24665 and not w24996;
w24998 <= w24639 and not w24651;
w24999 <= not w24650 and not w24651;
w25000 <= not w24998 and not w24999;
w25001 <= not w24997 and not w25000;
w25002 <= not w24651 and not w25001;
w25003 <= w24625 and not w24637;
w25004 <= not w24636 and not w24637;
w25005 <= not w25003 and not w25004;
w25006 <= not w25002 and not w25005;
w25007 <= not w24637 and not w25006;
w25008 <= not w24611 and w24622;
w25009 <= not w24623 and not w25008;
w25010 <= not w25007 and w25009;
w25011 <= not w24623 and not w25010;
w25012 <= not w24609 and not w25011;
w25013 <= not w24606 and not w25012;
w25014 <= not w24591 and not w25013;
w25015 <= not w24588 and not w25014;
w25016 <= w24559 and not w24574;
w25017 <= not w24573 and not w24574;
w25018 <= not w25016 and not w25017;
w25019 <= not w25015 and not w25018;
w25020 <= not w24574 and not w25019;
w25021 <= w24542 and not w24557;
w25022 <= not w24556 and not w24557;
w25023 <= not w25021 and not w25022;
w25024 <= not w25020 and not w25023;
w25025 <= not w24557 and not w25024;
w25026 <= w24526 and not w24540;
w25027 <= not w24539 and not w24540;
w25028 <= not w25026 and not w25027;
w25029 <= not w25025 and not w25028;
w25030 <= not w24540 and not w25029;
w25031 <= w7918 and w22264;
w25032 <= w7226 and w22270;
w25033 <= w7567 and w22267;
w25034 <= not w25032 and not w25033;
w25035 <= not w25031 and w25034;
w25036 <= w7229 and not w24568;
w25037 <= w25035 and not w25036;
w25038 <= a(11) and not w25037;
w25039 <= not w25037 and not w25038;
w25040 <= a(11) and not w25038;
w25041 <= not w25039 and not w25040;
w25042 <= not w24083 and not w24087;
w25043 <= w6168 and w22282;
w25044 <= w5598 and w22288;
w25045 <= w5874 and w22285;
w25046 <= not w25044 and not w25045;
w25047 <= not w25043 and w25046;
w25048 <= w5601 and not w23594;
w25049 <= w25047 and not w25048;
w25050 <= a(17) and not w25049;
w25051 <= not w25049 and not w25050;
w25052 <= a(17) and not w25050;
w25053 <= not w25051 and not w25052;
w25054 <= not w24054 and not w24058;
w25055 <= w4629 and w22300;
w25056 <= w4468 and w22306;
w25057 <= w4539 and w22303;
w25058 <= not w25056 and not w25057;
w25059 <= not w25055 and w25058;
w25060 <= w4471 and not w22928;
w25061 <= w25059 and not w25060;
w25062 <= a(23) and not w25061;
w25063 <= not w25061 and not w25062;
w25064 <= a(23) and not w25062;
w25065 <= not w25063 and not w25064;
w25066 <= not w24027 and not w24031;
w25067 <= w3392 and w22319;
w25068 <= w3477 and w22325;
w25069 <= w3541 and w22322;
w25070 <= not w25068 and not w25069;
w25071 <= not w25067 and w25070;
w25072 <= w3303 and w22741;
w25073 <= w25071 and not w25072;
w25074 <= a(29) and not w25073;
w25075 <= not w25073 and not w25074;
w25076 <= a(29) and not w25074;
w25077 <= not w25075 and not w25076;
w25078 <= not w24000 and not w24004;
w25079 <= w1546 and w5683;
w25080 <= w4204 and w25079;
w25081 <= w626 and w25080;
w25082 <= w139 and w25081;
w25083 <= w13495 and w25082;
w25084 <= w12867 and w25083;
w25085 <= w12844 and w25084;
w25086 <= w15859 and w25085;
w25087 <= w450 and w25086;
w25088 <= not w213 and w25087;
w25089 <= not w70 and w25088;
w25090 <= not w503 and w25089;
w25091 <= not w266 and w25090;
w25092 <= not w160 and w25091;
w25093 <= w2955 and w22328;
w25094 <= w2963 and w22331;
w25095 <= w2958 and w22334;
w25096 <= w10 and w22606;
w25097 <= not w25095 and not w25096;
w25098 <= not w25094 and w25097;
w25099 <= not w25093 and w25098;
w25100 <= not w25092 and not w25099;
w25101 <= not w25092 and not w25100;
w25102 <= not w25099 and not w25100;
w25103 <= not w25101 and not w25102;
w25104 <= not w25078 and not w25103;
w25105 <= not w25078 and not w25104;
w25106 <= not w25103 and not w25104;
w25107 <= not w25105 and not w25106;
w25108 <= not w25077 and not w25107;
w25109 <= not w25077 and not w25108;
w25110 <= not w25107 and not w25108;
w25111 <= not w25109 and not w25110;
w25112 <= not w24008 and not w24014;
w25113 <= w25111 and w25112;
w25114 <= not w25111 and not w25112;
w25115 <= not w25113 and not w25114;
w25116 <= w3819 and w22309;
w25117 <= w3902 and w22315;
w25118 <= w3981 and w22312;
w25119 <= not w25117 and not w25118;
w25120 <= not w25116 and w25119;
w25121 <= not w3985 and w25120;
w25122 <= not w22504 and w25120;
w25123 <= not w25121 and not w25122;
w25124 <= a(26) and not w25123;
w25125 <= not a(26) and w25123;
w25126 <= not w25124 and not w25125;
w25127 <= w25115 and not w25126;
w25128 <= w25115 and not w25127;
w25129 <= not w25126 and not w25127;
w25130 <= not w25128 and not w25129;
w25131 <= not w25066 and not w25130;
w25132 <= not w25066 and not w25131;
w25133 <= not w25130 and not w25131;
w25134 <= not w25132 and not w25133;
w25135 <= not w25065 and not w25134;
w25136 <= not w25065 and not w25135;
w25137 <= not w25134 and not w25135;
w25138 <= not w25136 and not w25137;
w25139 <= not w24035 and not w24041;
w25140 <= w25138 and w25139;
w25141 <= not w25138 and not w25139;
w25142 <= not w25140 and not w25141;
w25143 <= w5431 and w22291;
w25144 <= w4870 and w22297;
w25145 <= w5342 and w22294;
w25146 <= not w25144 and not w25145;
w25147 <= not w25143 and w25146;
w25148 <= not w4873 and w25147;
w25149 <= w23280 and w25147;
w25150 <= not w25148 and not w25149;
w25151 <= a(20) and not w25150;
w25152 <= not a(20) and w25150;
w25153 <= not w25151 and not w25152;
w25154 <= w25142 and not w25153;
w25155 <= w25142 and not w25154;
w25156 <= not w25153 and not w25154;
w25157 <= not w25155 and not w25156;
w25158 <= not w25054 and not w25157;
w25159 <= not w25054 and not w25158;
w25160 <= not w25157 and not w25158;
w25161 <= not w25159 and not w25160;
w25162 <= not w25053 and not w25161;
w25163 <= not w25053 and not w25162;
w25164 <= not w25161 and not w25162;
w25165 <= not w25163 and not w25164;
w25166 <= not w24062 and not w24068;
w25167 <= w25165 and w25166;
w25168 <= not w25165 and not w25166;
w25169 <= not w25167 and not w25168;
w25170 <= w7036 and w22273;
w25171 <= w6337 and w22279;
w25172 <= w6886 and w22276;
w25173 <= not w25171 and not w25172;
w25174 <= not w25170 and w25173;
w25175 <= not w6332 and w25174;
w25176 <= w24123 and w25174;
w25177 <= not w25175 and not w25176;
w25178 <= a(14) and not w25177;
w25179 <= not a(14) and w25177;
w25180 <= not w25178 and not w25179;
w25181 <= w25169 and not w25180;
w25182 <= w25169 and not w25181;
w25183 <= not w25180 and not w25181;
w25184 <= not w25182 and not w25183;
w25185 <= not w25042 and not w25184;
w25186 <= not w25042 and not w25185;
w25187 <= not w25184 and not w25185;
w25188 <= not w25186 and not w25187;
w25189 <= not w25041 and not w25188;
w25190 <= not w25041 and not w25189;
w25191 <= not w25188 and not w25189;
w25192 <= not w25190 and not w25191;
w25193 <= not w24091 and not w24525;
w25194 <= w25192 and w25193;
w25195 <= not w25192 and not w25193;
w25196 <= not w25194 and not w25195;
w25197 <= w9266 and w22255;
w25198 <= w8353 and w22261;
w25199 <= w8795 and w22258;
w25200 <= not w25198 and not w25199;
w25201 <= not w25197 and w25200;
w25202 <= not w8356 and w25201;
w25203 <= not w22443 and not w22446;
w25204 <= not w22444 and w22447;
w25205 <= not w25203 and not w25204;
w25206 <= w25201 and w25205;
w25207 <= not w25202 and not w25206;
w25208 <= a(8) and not w25207;
w25209 <= not a(8) and w25207;
w25210 <= not w25208 and not w25209;
w25211 <= w25196 and not w25210;
w25212 <= w25196 and not w25211;
w25213 <= not w25210 and not w25211;
w25214 <= not w25212 and not w25213;
w25215 <= not w25030 and not w25214;
w25216 <= not w25030 and not w25215;
w25217 <= not w25214 and not w25215;
w25218 <= not w25216 and not w25217;
w25219 <= not w22470 and not w25218;
w25220 <= not w22470 and not w25219;
w25221 <= not w25218 and not w25219;
w25222 <= not w25220 and not w25221;
w25223 <= w6 and w22250;
w25224 <= w9802 and w22255;
w25225 <= w10369 and w22247;
w25226 <= not w25224 and not w25225;
w25227 <= not w25223 and w25226;
w25228 <= w22451 and not w22454;
w25229 <= not w22455 and not w25228;
w25230 <= w9805 and w25229;
w25231 <= w25227 and not w25230;
w25232 <= a(5) and not w25231;
w25233 <= not w25231 and not w25232;
w25234 <= a(5) and not w25232;
w25235 <= not w25233 and not w25234;
w25236 <= not w25025 and not w25029;
w25237 <= not w25028 and not w25029;
w25238 <= not w25236 and not w25237;
w25239 <= not w25235 and not w25238;
w25240 <= not w25235 and not w25239;
w25241 <= not w25238 and not w25239;
w25242 <= not w25240 and not w25241;
w25243 <= w6 and w22247;
w25244 <= w9802 and w22258;
w25245 <= w10369 and w22255;
w25246 <= not w25244 and not w25245;
w25247 <= not w25243 and w25246;
w25248 <= not w22447 and not w22450;
w25249 <= not w22448 and w22451;
w25250 <= not w25248 and not w25249;
w25251 <= w9805 and not w25250;
w25252 <= w25247 and not w25251;
w25253 <= a(5) and not w25252;
w25254 <= not w25252 and not w25253;
w25255 <= a(5) and not w25253;
w25256 <= not w25254 and not w25255;
w25257 <= not w25020 and not w25024;
w25258 <= not w25023 and not w25024;
w25259 <= not w25257 and not w25258;
w25260 <= not w25256 and not w25259;
w25261 <= not w25256 and not w25260;
w25262 <= not w25259 and not w25260;
w25263 <= not w25261 and not w25262;
w25264 <= w6 and w22255;
w25265 <= w9802 and w22261;
w25266 <= w10369 and w22258;
w25267 <= not w25265 and not w25266;
w25268 <= not w25264 and w25267;
w25269 <= w9805 and not w25205;
w25270 <= w25268 and not w25269;
w25271 <= a(5) and not w25270;
w25272 <= not w25270 and not w25271;
w25273 <= a(5) and not w25271;
w25274 <= not w25272 and not w25273;
w25275 <= not w25015 and not w25019;
w25276 <= not w25018 and not w25019;
w25277 <= not w25275 and not w25276;
w25278 <= not w25274 and not w25277;
w25279 <= not w25274 and not w25278;
w25280 <= not w25277 and not w25278;
w25281 <= not w25279 and not w25280;
w25282 <= w24591 and w25013;
w25283 <= not w25014 and not w25282;
w25284 <= w6 and w22258;
w25285 <= w9802 and w22264;
w25286 <= w10369 and w22261;
w25287 <= not w25285 and not w25286;
w25288 <= not w25284 and w25287;
w25289 <= not w9805 and w25288;
w25290 <= not w24534 and w25288;
w25291 <= not w25289 and not w25290;
w25292 <= a(5) and not w25291;
w25293 <= not a(5) and w25291;
w25294 <= not w25292 and not w25293;
w25295 <= w25283 and not w25294;
w25296 <= w24609 and w25011;
w25297 <= not w25012 and not w25296;
w25298 <= w6 and w22261;
w25299 <= w9802 and w22267;
w25300 <= w10369 and w22264;
w25301 <= not w25299 and not w25300;
w25302 <= not w25298 and w25301;
w25303 <= not w9805 and w25302;
w25304 <= w24551 and w25302;
w25305 <= not w25303 and not w25304;
w25306 <= a(5) and not w25305;
w25307 <= not a(5) and w25305;
w25308 <= not w25306 and not w25307;
w25309 <= w25297 and not w25308;
w25310 <= w6 and w22264;
w25311 <= w9802 and w22270;
w25312 <= w10369 and w22267;
w25313 <= not w25311 and not w25312;
w25314 <= not w25310 and w25313;
w25315 <= w9805 and not w24568;
w25316 <= w25314 and not w25315;
w25317 <= a(5) and not w25316;
w25318 <= not w25316 and not w25317;
w25319 <= a(5) and not w25317;
w25320 <= not w25318 and not w25319;
w25321 <= w25007 and not w25009;
w25322 <= not w25010 and not w25321;
w25323 <= not w25320 and w25322;
w25324 <= not w25320 and not w25323;
w25325 <= w25322 and not w25323;
w25326 <= not w25324 and not w25325;
w25327 <= w6 and w22267;
w25328 <= w9802 and w22273;
w25329 <= w10369 and w22270;
w25330 <= not w25328 and not w25329;
w25331 <= not w25327 and w25330;
w25332 <= w9805 and w22477;
w25333 <= w25331 and not w25332;
w25334 <= a(5) and not w25333;
w25335 <= not w25333 and not w25334;
w25336 <= a(5) and not w25334;
w25337 <= not w25335 and not w25336;
w25338 <= not w25002 and not w25006;
w25339 <= not w25005 and not w25006;
w25340 <= not w25338 and not w25339;
w25341 <= not w25337 and not w25340;
w25342 <= not w25337 and not w25341;
w25343 <= not w25340 and not w25341;
w25344 <= not w25342 and not w25343;
w25345 <= w6 and w22270;
w25346 <= w9802 and w22276;
w25347 <= w10369 and w22273;
w25348 <= not w25346 and not w25347;
w25349 <= not w25345 and w25348;
w25350 <= w9805 and not w24102;
w25351 <= w25349 and not w25350;
w25352 <= a(5) and not w25351;
w25353 <= not w25351 and not w25352;
w25354 <= a(5) and not w25352;
w25355 <= not w25353 and not w25354;
w25356 <= not w24997 and not w25001;
w25357 <= not w25000 and not w25001;
w25358 <= not w25356 and not w25357;
w25359 <= not w25355 and not w25358;
w25360 <= not w25355 and not w25359;
w25361 <= not w25358 and not w25359;
w25362 <= not w25360 and not w25361;
w25363 <= w24668 and w24995;
w25364 <= not w24996 and not w25363;
w25365 <= w6 and w22273;
w25366 <= w9802 and w22279;
w25367 <= w10369 and w22276;
w25368 <= not w25366 and not w25367;
w25369 <= not w25365 and w25368;
w25370 <= not w9805 and w25369;
w25371 <= w24123 and w25369;
w25372 <= not w25370 and not w25371;
w25373 <= a(5) and not w25372;
w25374 <= not a(5) and w25372;
w25375 <= not w25373 and not w25374;
w25376 <= w25364 and not w25375;
w25377 <= w24686 and w24993;
w25378 <= not w24994 and not w25377;
w25379 <= w6 and w22276;
w25380 <= w9802 and w22282;
w25381 <= w10369 and w22279;
w25382 <= not w25380 and not w25381;
w25383 <= not w25379 and w25382;
w25384 <= not w9805 and w25383;
w25385 <= not w24077 and w25383;
w25386 <= not w25384 and not w25385;
w25387 <= a(5) and not w25386;
w25388 <= not a(5) and w25386;
w25389 <= not w25387 and not w25388;
w25390 <= w25378 and not w25389;
w25391 <= w24704 and w24991;
w25392 <= not w24992 and not w25391;
w25393 <= w6 and w22279;
w25394 <= w9802 and w22285;
w25395 <= w10369 and w22282;
w25396 <= not w25394 and not w25395;
w25397 <= not w25393 and w25396;
w25398 <= not w9805 and w25397;
w25399 <= w23577 and w25397;
w25400 <= not w25398 and not w25399;
w25401 <= a(5) and not w25400;
w25402 <= not a(5) and w25400;
w25403 <= not w25401 and not w25402;
w25404 <= w25392 and not w25403;
w25405 <= w6 and w22282;
w25406 <= w9802 and w22288;
w25407 <= w10369 and w22285;
w25408 <= not w25406 and not w25407;
w25409 <= not w25405 and w25408;
w25410 <= w9805 and not w23594;
w25411 <= w25409 and not w25410;
w25412 <= a(5) and not w25411;
w25413 <= not w25411 and not w25412;
w25414 <= a(5) and not w25412;
w25415 <= not w25413 and not w25414;
w25416 <= w24987 and not w24989;
w25417 <= not w24990 and not w25416;
w25418 <= not w25415 and w25417;
w25419 <= not w25415 and not w25418;
w25420 <= w25417 and not w25418;
w25421 <= not w25419 and not w25420;
w25422 <= w6 and w22285;
w25423 <= w9802 and w22291;
w25424 <= w10369 and w22288;
w25425 <= not w25423 and not w25424;
w25426 <= not w25422 and w25425;
w25427 <= w9805 and w23607;
w25428 <= w25426 and not w25427;
w25429 <= a(5) and not w25428;
w25430 <= not w25428 and not w25429;
w25431 <= a(5) and not w25429;
w25432 <= not w25430 and not w25431;
w25433 <= not w24982 and not w24986;
w25434 <= not w24985 and not w24986;
w25435 <= not w25433 and not w25434;
w25436 <= not w25432 and not w25435;
w25437 <= not w25432 and not w25436;
w25438 <= not w25435 and not w25436;
w25439 <= not w25437 and not w25438;
w25440 <= w6 and w22288;
w25441 <= w9802 and w22294;
w25442 <= w10369 and w22291;
w25443 <= not w25441 and not w25442;
w25444 <= not w25440 and w25443;
w25445 <= w9805 and not w22491;
w25446 <= w25444 and not w25445;
w25447 <= a(5) and not w25446;
w25448 <= not w25446 and not w25447;
w25449 <= a(5) and not w25447;
w25450 <= not w25448 and not w25449;
w25451 <= not w24977 and not w24981;
w25452 <= not w24980 and not w24981;
w25453 <= not w25451 and not w25452;
w25454 <= not w25450 and not w25453;
w25455 <= not w25450 and not w25454;
w25456 <= not w25453 and not w25454;
w25457 <= not w25455 and not w25456;
w25458 <= w24763 and w24975;
w25459 <= not w24976 and not w25458;
w25460 <= w6 and w22291;
w25461 <= w9802 and w22297;
w25462 <= w10369 and w22294;
w25463 <= not w25461 and not w25462;
w25464 <= not w25460 and w25463;
w25465 <= not w9805 and w25464;
w25466 <= w23280 and w25464;
w25467 <= not w25465 and not w25466;
w25468 <= a(5) and not w25467;
w25469 <= not a(5) and w25467;
w25470 <= not w25468 and not w25469;
w25471 <= w25459 and not w25470;
w25472 <= w24781 and w24973;
w25473 <= not w24974 and not w25472;
w25474 <= w6 and w22294;
w25475 <= w9802 and w22300;
w25476 <= w10369 and w22297;
w25477 <= not w25475 and not w25476;
w25478 <= not w25474 and w25477;
w25479 <= not w9805 and w25478;
w25480 <= not w23303 and w25478;
w25481 <= not w25479 and not w25480;
w25482 <= a(5) and not w25481;
w25483 <= not a(5) and w25481;
w25484 <= not w25482 and not w25483;
w25485 <= w25473 and not w25484;
w25486 <= w24799 and w24971;
w25487 <= not w24972 and not w25486;
w25488 <= w6 and w22297;
w25489 <= w9802 and w22303;
w25490 <= w10369 and w22300;
w25491 <= not w25489 and not w25490;
w25492 <= not w25488 and w25491;
w25493 <= not w9805 and w25492;
w25494 <= w23255 and w25492;
w25495 <= not w25493 and not w25494;
w25496 <= a(5) and not w25495;
w25497 <= not a(5) and w25495;
w25498 <= not w25496 and not w25497;
w25499 <= w25487 and not w25498;
w25500 <= w6 and w22300;
w25501 <= w9802 and w22306;
w25502 <= w10369 and w22303;
w25503 <= not w25501 and not w25502;
w25504 <= not w25500 and w25503;
w25505 <= w9805 and not w22928;
w25506 <= w25504 and not w25505;
w25507 <= a(5) and not w25506;
w25508 <= not w25506 and not w25507;
w25509 <= a(5) and not w25507;
w25510 <= not w25508 and not w25509;
w25511 <= w24967 and not w24969;
w25512 <= not w24970 and not w25511;
w25513 <= not w25510 and w25512;
w25514 <= not w25510 and not w25513;
w25515 <= w25512 and not w25513;
w25516 <= not w25514 and not w25515;
w25517 <= w6 and w22303;
w25518 <= w9802 and w22309;
w25519 <= w10369 and w22306;
w25520 <= not w25518 and not w25519;
w25521 <= not w25517 and w25520;
w25522 <= w9805 and w22941;
w25523 <= w25521 and not w25522;
w25524 <= a(5) and not w25523;
w25525 <= not w25523 and not w25524;
w25526 <= a(5) and not w25524;
w25527 <= not w25525 and not w25526;
w25528 <= not w24962 and not w24966;
w25529 <= not w24965 and not w24966;
w25530 <= not w25528 and not w25529;
w25531 <= not w25527 and not w25530;
w25532 <= not w25527 and not w25531;
w25533 <= not w25530 and not w25531;
w25534 <= not w25532 and not w25533;
w25535 <= w6 and w22306;
w25536 <= w9802 and w22312;
w25537 <= w10369 and w22309;
w25538 <= not w25536 and not w25537;
w25539 <= not w25535 and w25538;
w25540 <= w9805 and w22960;
w25541 <= w25539 and not w25540;
w25542 <= a(5) and not w25541;
w25543 <= not w25541 and not w25542;
w25544 <= a(5) and not w25542;
w25545 <= not w25543 and not w25544;
w25546 <= not w24957 and not w24961;
w25547 <= not w24960 and not w24961;
w25548 <= not w25546 and not w25547;
w25549 <= not w25545 and not w25548;
w25550 <= not w25545 and not w25549;
w25551 <= not w25548 and not w25549;
w25552 <= not w25550 and not w25551;
w25553 <= w24858 and w24955;
w25554 <= not w24956 and not w25553;
w25555 <= w6 and w22309;
w25556 <= w9802 and w22315;
w25557 <= w10369 and w22312;
w25558 <= not w25556 and not w25557;
w25559 <= not w25555 and w25558;
w25560 <= not w9805 and w25559;
w25561 <= not w22504 and w25559;
w25562 <= not w25560 and not w25561;
w25563 <= a(5) and not w25562;
w25564 <= not a(5) and w25562;
w25565 <= not w25563 and not w25564;
w25566 <= w25554 and not w25565;
w25567 <= w24951 and not w24953;
w25568 <= not w24954 and not w25567;
w25569 <= w6 and w22312;
w25570 <= w9802 and w22319;
w25571 <= w10369 and w22315;
w25572 <= not w25570 and not w25571;
w25573 <= not w25569 and w25572;
w25574 <= not w9805 and w25573;
w25575 <= w22769 and w25573;
w25576 <= not w25574 and not w25575;
w25577 <= a(5) and not w25576;
w25578 <= not a(5) and w25576;
w25579 <= not w25577 and not w25578;
w25580 <= w25568 and not w25579;
w25581 <= w24890 and w24949;
w25582 <= not w24950 and not w25581;
w25583 <= w6 and w22315;
w25584 <= w9802 and w22322;
w25585 <= w10369 and w22319;
w25586 <= not w25584 and not w25585;
w25587 <= not w25583 and w25586;
w25588 <= not w9805 and w25587;
w25589 <= not w22785 and w25587;
w25590 <= not w25588 and not w25589;
w25591 <= a(5) and not w25590;
w25592 <= not a(5) and w25590;
w25593 <= not w25591 and not w25592;
w25594 <= w25582 and not w25593;
w25595 <= w6 and w22319;
w25596 <= w9802 and w22325;
w25597 <= w10369 and w22322;
w25598 <= not w25596 and not w25597;
w25599 <= not w25595 and w25598;
w25600 <= w9805 and w22741;
w25601 <= w25599 and not w25600;
w25602 <= a(5) and not w25601;
w25603 <= not w25601 and not w25602;
w25604 <= a(5) and not w25602;
w25605 <= not w25603 and not w25604;
w25606 <= w24945 and not w24947;
w25607 <= not w24948 and not w25606;
w25608 <= not w25605 and w25607;
w25609 <= not w25605 and not w25608;
w25610 <= w25607 and not w25608;
w25611 <= not w25609 and not w25610;
w25612 <= not w24932 and not w24944;
w25613 <= not w24943 and not w24944;
w25614 <= not w25612 and not w25613;
w25615 <= w6 and w22322;
w25616 <= w9802 and w22328;
w25617 <= w10369 and w22325;
w25618 <= not w25616 and not w25617;
w25619 <= not w25615 and w25618;
w25620 <= not w9805 and w25619;
w25621 <= not w22517 and w25619;
w25622 <= not w25620 and not w25621;
w25623 <= a(5) and not w25622;
w25624 <= not a(5) and w25622;
w25625 <= not w25623 and not w25624;
w25626 <= not w25614 and not w25625;
w25627 <= w6 and w22325;
w25628 <= w9802 and w22331;
w25629 <= w10369 and w22328;
w25630 <= not w25628 and not w25629;
w25631 <= not w25627 and w25630;
w25632 <= w9805 and w22584;
w25633 <= w25631 and not w25632;
w25634 <= a(5) and not w25633;
w25635 <= not w25633 and not w25634;
w25636 <= a(5) and not w25634;
w25637 <= not w25635 and not w25636;
w25638 <= not w24916 and w24927;
w25639 <= not w24928 and not w25638;
w25640 <= not w25637 and w25639;
w25641 <= not w25637 and not w25640;
w25642 <= w25639 and not w25640;
w25643 <= not w25641 and not w25642;
w25644 <= w24913 and not w24915;
w25645 <= not w24916 and not w25644;
w25646 <= w6 and w22328;
w25647 <= w9802 and w22334;
w25648 <= w10369 and w22331;
w25649 <= not w25647 and not w25648;
w25650 <= not w25646 and w25649;
w25651 <= not w9805 and w25650;
w25652 <= not w22606 and w25650;
w25653 <= not w25651 and not w25652;
w25654 <= a(5) and not w25653;
w25655 <= not a(5) and w25653;
w25656 <= not w25654 and not w25655;
w25657 <= w25645 and not w25656;
w25658 <= w10369 and not w22341;
w25659 <= w6 and w22337;
w25660 <= not w25658 and not w25659;
w25661 <= w9805 and not w22544;
w25662 <= w25660 and not w25661;
w25663 <= a(5) and not w25662;
w25664 <= a(5) and not w25663;
w25665 <= not w25662 and not w25663;
w25666 <= not w25664 and not w25665;
w25667 <= not w5 and not w22341;
w25668 <= a(5) and not w25667;
w25669 <= not w25666 and w25668;
w25670 <= w6 and w22334;
w25671 <= w9802 and not w22341;
w25672 <= w10369 and w22337;
w25673 <= not w25671 and not w25672;
w25674 <= not w25670 and w25673;
w25675 <= not w9805 and w25674;
w25676 <= w22560 and w25674;
w25677 <= not w25675 and not w25676;
w25678 <= a(5) and not w25677;
w25679 <= not a(5) and w25677;
w25680 <= not w25678 and not w25679;
w25681 <= w25669 and not w25680;
w25682 <= w24914 and w25681;
w25683 <= w25681 and not w25682;
w25684 <= w24914 and not w25682;
w25685 <= not w25683 and not w25684;
w25686 <= w6 and w22331;
w25687 <= w9802 and w22337;
w25688 <= w10369 and w22334;
w25689 <= not w25687 and not w25688;
w25690 <= not w25686 and w25689;
w25691 <= w9805 and w22530;
w25692 <= w25690 and not w25691;
w25693 <= a(5) and not w25692;
w25694 <= a(5) and not w25693;
w25695 <= not w25692 and not w25693;
w25696 <= not w25694 and not w25695;
w25697 <= not w25685 and not w25696;
w25698 <= not w25682 and not w25697;
w25699 <= not w25645 and w25656;
w25700 <= not w25657 and not w25699;
w25701 <= not w25698 and w25700;
w25702 <= not w25657 and not w25701;
w25703 <= not w25643 and not w25702;
w25704 <= not w25640 and not w25703;
w25705 <= w25614 and w25625;
w25706 <= not w25626 and not w25705;
w25707 <= not w25704 and w25706;
w25708 <= not w25626 and not w25707;
w25709 <= not w25611 and not w25708;
w25710 <= not w25608 and not w25709;
w25711 <= w25582 and not w25594;
w25712 <= not w25593 and not w25594;
w25713 <= not w25711 and not w25712;
w25714 <= not w25710 and not w25713;
w25715 <= not w25594 and not w25714;
w25716 <= w25568 and not w25580;
w25717 <= not w25579 and not w25580;
w25718 <= not w25716 and not w25717;
w25719 <= not w25715 and not w25718;
w25720 <= not w25580 and not w25719;
w25721 <= not w25554 and w25565;
w25722 <= not w25566 and not w25721;
w25723 <= not w25720 and w25722;
w25724 <= not w25566 and not w25723;
w25725 <= not w25552 and not w25724;
w25726 <= not w25549 and not w25725;
w25727 <= not w25534 and not w25726;
w25728 <= not w25531 and not w25727;
w25729 <= not w25516 and not w25728;
w25730 <= not w25513 and not w25729;
w25731 <= w25487 and not w25499;
w25732 <= not w25498 and not w25499;
w25733 <= not w25731 and not w25732;
w25734 <= not w25730 and not w25733;
w25735 <= not w25499 and not w25734;
w25736 <= w25473 and not w25485;
w25737 <= not w25484 and not w25485;
w25738 <= not w25736 and not w25737;
w25739 <= not w25735 and not w25738;
w25740 <= not w25485 and not w25739;
w25741 <= not w25459 and w25470;
w25742 <= not w25471 and not w25741;
w25743 <= not w25740 and w25742;
w25744 <= not w25471 and not w25743;
w25745 <= not w25457 and not w25744;
w25746 <= not w25454 and not w25745;
w25747 <= not w25439 and not w25746;
w25748 <= not w25436 and not w25747;
w25749 <= not w25421 and not w25748;
w25750 <= not w25418 and not w25749;
w25751 <= w25392 and not w25404;
w25752 <= not w25403 and not w25404;
w25753 <= not w25751 and not w25752;
w25754 <= not w25750 and not w25753;
w25755 <= not w25404 and not w25754;
w25756 <= w25378 and not w25390;
w25757 <= not w25389 and not w25390;
w25758 <= not w25756 and not w25757;
w25759 <= not w25755 and not w25758;
w25760 <= not w25390 and not w25759;
w25761 <= not w25364 and w25375;
w25762 <= not w25376 and not w25761;
w25763 <= not w25760 and w25762;
w25764 <= not w25376 and not w25763;
w25765 <= not w25362 and not w25764;
w25766 <= not w25359 and not w25765;
w25767 <= not w25344 and not w25766;
w25768 <= not w25341 and not w25767;
w25769 <= not w25326 and not w25768;
w25770 <= not w25323 and not w25769;
w25771 <= w25297 and not w25309;
w25772 <= not w25308 and not w25309;
w25773 <= not w25771 and not w25772;
w25774 <= not w25770 and not w25773;
w25775 <= not w25309 and not w25774;
w25776 <= not w25283 and w25294;
w25777 <= not w25295 and not w25776;
w25778 <= not w25775 and w25777;
w25779 <= not w25295 and not w25778;
w25780 <= not w25281 and not w25779;
w25781 <= not w25278 and not w25780;
w25782 <= not w25263 and not w25781;
w25783 <= not w25260 and not w25782;
w25784 <= not w25242 and not w25783;
w25785 <= not w25239 and not w25784;
w25786 <= w25222 and w25785;
w25787 <= not w25222 and not w25785;
w25788 <= not w25786 and not w25787;
w25789 <= not w22219 and not w22232;
w25790 <= not w22210 and not w22213;
w25791 <= not w22205 and not w22207;
w25792 <= w709 and w6651;
w25793 <= w1759 and w25792;
w25794 <= w3821 and w25793;
w25795 <= not w554 and w25794;
w25796 <= not w387 and w25795;
w25797 <= not w1138 and w25796;
w25798 <= not w172 and w25797;
w25799 <= w727 and w12998;
w25800 <= w3367 and w25799;
w25801 <= w3699 and w25800;
w25802 <= w3340 and w25801;
w25803 <= w1536 and w25802;
w25804 <= w25798 and w25803;
w25805 <= w2211 and w25804;
w25806 <= w1302 and w25805;
w25807 <= not w299 and w25806;
w25808 <= not w430 and w25807;
w25809 <= not w231 and w25808;
w25810 <= not w25791 and w25809;
w25811 <= w25791 and not w25809;
w25812 <= not w25810 and not w25811;
w25813 <= w2955 and w13450;
w25814 <= w2963 and w13456;
w25815 <= w2958 and w13453;
w25816 <= w10 and w13476;
w25817 <= not w25815 and not w25816;
w25818 <= not w25814 and w25817;
w25819 <= not w25813 and w25818;
w25820 <= w25812 and not w25819;
w25821 <= not w25812 and w25819;
w25822 <= not w25820 and not w25821;
w25823 <= not w25790 and w25822;
w25824 <= w25790 and not w25822;
w25825 <= not w25823 and not w25824;
w25826 <= w3392 and w13568;
w25827 <= w3477 and w13532;
w25828 <= w3541 and w13565;
w25829 <= not w25827 and not w25828;
w25830 <= not w25826 and w25829;
w25831 <= not w3303 and w25830;
w25832 <= not w13864 and w25830;
w25833 <= not w25831 and not w25832;
w25834 <= a(29) and not w25833;
w25835 <= not a(29) and w25833;
w25836 <= not w25834 and not w25835;
w25837 <= w25825 and not w25836;
w25838 <= not w25825 and w25836;
w25839 <= not w25837 and not w25838;
w25840 <= not w25789 and w25839;
w25841 <= w25789 and not w25839;
w25842 <= not w25840 and not w25841;
w25843 <= w3819 and not w13373;
w25844 <= w3902 and not w13562;
w25845 <= w3981 and w13876;
w25846 <= not w25844 and not w25845;
w25847 <= not w25843 and w25846;
w25848 <= w3985 and w13963;
w25849 <= w25847 and not w25848;
w25850 <= a(26) and not w25849;
w25851 <= a(26) and not w25850;
w25852 <= not w25849 and not w25850;
w25853 <= not w25851 and not w25852;
w25854 <= w25842 and not w25853;
w25855 <= not w25840 and not w25854;
w25856 <= w10 and not w13547;
w25857 <= w2955 and w13532;
w25858 <= w2958 and w13456;
w25859 <= w2963 and w13450;
w25860 <= not w25858 and not w25859;
w25861 <= not w25857 and w25860;
w25862 <= not w25856 and w25861;
w25863 <= w408 and w982;
w25864 <= w3913 and w25863;
w25865 <= w3717 and w25864;
w25866 <= w12998 and w25865;
w25867 <= w1666 and w25866;
w25868 <= w2105 and w25867;
w25869 <= w3692 and w25868;
w25870 <= not w681 and w25869;
w25871 <= not w231 and w25870;
w25872 <= not w108 and w25871;
w25873 <= not w536 and w25872;
w25874 <= not w180 and w25873;
w25875 <= not w77 and w25874;
w25876 <= not w25809 and w25875;
w25877 <= w25809 and not w25875;
w25878 <= not w25862 and not w25877;
w25879 <= not w25876 and w25878;
w25880 <= not w25862 and not w25879;
w25881 <= not w25877 and not w25879;
w25882 <= not w25876 and w25881;
w25883 <= not w25880 and not w25882;
w25884 <= not w25810 and not w25820;
w25885 <= w25883 and w25884;
w25886 <= not w25883 and not w25884;
w25887 <= not w25885 and not w25886;
w25888 <= not w25823 and not w25837;
w25889 <= not w25887 and w25888;
w25890 <= w25887 and not w25888;
w25891 <= not w25889 and not w25890;
w25892 <= not w3819 and not w3981;
w25893 <= not w13373 and not w25892;
w25894 <= w3902 and w13876;
w25895 <= not w25893 and not w25894;
w25896 <= w3985 and not w13886;
w25897 <= w25895 and not w25896;
w25898 <= a(26) and not w25897;
w25899 <= not w25897 and not w25898;
w25900 <= a(26) and not w25898;
w25901 <= not w25899 and not w25900;
w25902 <= w3392 and not w13562;
w25903 <= w3477 and w13565;
w25904 <= w3541 and w13568;
w25905 <= not w25903 and not w25904;
w25906 <= not w25902 and w25905;
w25907 <= w3303 and not w13589;
w25908 <= w25906 and not w25907;
w25909 <= a(29) and not w25908;
w25910 <= a(29) and not w25909;
w25911 <= not w25908 and not w25909;
w25912 <= not w25910 and not w25911;
w25913 <= not w25901 and not w25912;
w25914 <= not w25901 and not w25913;
w25915 <= not w25912 and not w25913;
w25916 <= not w25914 and not w25915;
w25917 <= not w25891 and w25916;
w25918 <= w25891 and not w25916;
w25919 <= not w25917 and not w25918;
w25920 <= not w25855 and w25919;
w25921 <= w25842 and not w25854;
w25922 <= not w25853 and not w25854;
w25923 <= not w25921 and not w25922;
w25924 <= not w22174 and not w22235;
w25925 <= not w22171 and not w25924;
w25926 <= not w25923 and not w25925;
w25927 <= not w25923 and not w25926;
w25928 <= not w25925 and not w25926;
w25929 <= not w25927 and not w25928;
w25930 <= not w22239 and not w22242;
w25931 <= not w25929 and not w25930;
w25932 <= not w25926 and not w25931;
w25933 <= w25855 and not w25919;
w25934 <= not w25920 and not w25933;
w25935 <= not w25932 and w25934;
w25936 <= not w25920 and not w25935;
w25937 <= w10 and w13911;
w25938 <= w2955 and w13565;
w25939 <= w2958 and w13450;
w25940 <= w2963 and w13532;
w25941 <= not w25939 and not w25940;
w25942 <= not w25938 and w25941;
w25943 <= not w25937 and w25942;
w25944 <= not w3902 and w25892;
w25945 <= not w3985 and w25944;
w25946 <= not w13373 and not w25945;
w25947 <= a(26) and not w25946;
w25948 <= not a(26) and w25946;
w25949 <= not w25947 and not w25948;
w25950 <= w3808 and w3907;
w25951 <= not w231 and w25950;
w25952 <= w3952 and w3975;
w25953 <= w2675 and w25952;
w25954 <= w25951 and w25953;
w25955 <= not w263 and w25954;
w25956 <= not w536 and w25955;
w25957 <= w25809 and w25956;
w25958 <= not w25809 and not w25956;
w25959 <= not w25957 and not w25958;
w25960 <= w25949 and w25959;
w25961 <= not w25949 and not w25959;
w25962 <= not w25960 and not w25961;
w25963 <= not w25881 and w25962;
w25964 <= w25881 and not w25962;
w25965 <= not w25963 and not w25964;
w25966 <= not w25943 and w25965;
w25967 <= w25965 and not w25966;
w25968 <= not w25943 and not w25966;
w25969 <= not w25967 and not w25968;
w25970 <= w3392 and w13876;
w25971 <= w3477 and w13568;
w25972 <= w3541 and not w13562;
w25973 <= not w25971 and not w25972;
w25974 <= not w25970 and w25973;
w25975 <= w3303 and w14071;
w25976 <= w25974 and not w25975;
w25977 <= a(29) and not w25976;
w25978 <= a(29) and not w25977;
w25979 <= not w25976 and not w25977;
w25980 <= not w25978 and not w25979;
w25981 <= not w25969 and not w25980;
w25982 <= not w25969 and not w25981;
w25983 <= not w25980 and not w25981;
w25984 <= not w25982 and not w25983;
w25985 <= not w25886 and not w25890;
w25986 <= w25984 and w25985;
w25987 <= not w25984 and not w25985;
w25988 <= not w25986 and not w25987;
w25989 <= not w25913 and not w25918;
w25990 <= w25988 and not w25989;
w25991 <= not w25988 and w25989;
w25992 <= not w25990 and not w25991;
w25993 <= w25936 and not w25992;
w25994 <= not w25936 and w25992;
w25995 <= not w25993 and not w25994;
w25996 <= w11662 and w25995;
w25997 <= w25929 and w25930;
w25998 <= not w25931 and not w25997;
w25999 <= w10990 and w25998;
w26000 <= w25932 and not w25934;
w26001 <= not w25935 and not w26000;
w26002 <= w11650 and w26001;
w26003 <= not w25999 and not w26002;
w26004 <= not w25996 and w26003;
w26005 <= not w10992 and w26004;
w26006 <= w25998 and w26001;
w26007 <= w22244 and w25998;
w26008 <= not w22244 and not w25998;
w26009 <= not w22462 and not w26008;
w26010 <= not w26007 and w26009;
w26011 <= not w26007 and not w26010;
w26012 <= not w25998 and not w26001;
w26013 <= not w26011 and not w26012;
w26014 <= not w26006 and w26013;
w26015 <= not w26006 and not w26014;
w26016 <= w25995 and w26001;
w26017 <= not w25995 and not w26001;
w26018 <= not w26015 and not w26017;
w26019 <= not w26016 and w26018;
w26020 <= not w26015 and not w26019;
w26021 <= not w26016 and not w26019;
w26022 <= not w26017 and w26021;
w26023 <= not w26020 and not w26022;
w26024 <= w26004 and w26023;
w26025 <= not w26005 and not w26024;
w26026 <= a(2) and not w26025;
w26027 <= not a(2) and w26025;
w26028 <= not w26026 and not w26027;
w26029 <= w25788 and not w26028;
w26030 <= w25775 and not w25777;
w26031 <= not w25778 and not w26030;
w26032 <= w25760 and not w25762;
w26033 <= not w25763 and not w26032;
w26034 <= w25740 and not w25742;
w26035 <= not w25743 and not w26034;
w26036 <= w25720 and not w25722;
w26037 <= not w25723 and not w26036;
w26038 <= w25698 and not w25700;
w26039 <= not w25701 and not w26038;
w26040 <= not w25669 and w25680;
w26041 <= not w25681 and not w26040;
w26042 <= not w11729 and not w22341;
w26043 <= w11731 and not w22560;
w26044 <= w11662 and w22334;
w26045 <= w10990 and not w22341;
w26046 <= w11650 and w22337;
w26047 <= not w26045 and not w26046;
w26048 <= not w26044 and w26047;
w26049 <= a(2) and not w26048;
w26050 <= w11731 and not w22544;
w26051 <= w11740 and not w22341;
w26052 <= w11742 and w22337;
w26053 <= a(2) and not w26052;
w26054 <= not w26051 and w26053;
w26055 <= not w26050 and w26054;
w26056 <= not w26049 and w26055;
w26057 <= not w26043 and w26056;
w26058 <= not w26042 and w26057;
w26059 <= w25667 and w26058;
w26060 <= not w25667 and not w26058;
w26061 <= w11662 and w22331;
w26062 <= w10990 and w22337;
w26063 <= w11650 and w22334;
w26064 <= not w26062 and not w26063;
w26065 <= not w26061 and w26064;
w26066 <= w10992 and w22530;
w26067 <= w26065 and not w26066;
w26068 <= not a(2) and not w26067;
w26069 <= a(2) and w26067;
w26070 <= not w26068 and not w26069;
w26071 <= not w26060 and not w26070;
w26072 <= not w26059 and not w26071;
w26073 <= w11662 and w22328;
w26074 <= w10990 and w22334;
w26075 <= w11650 and w22331;
w26076 <= not w26074 and not w26075;
w26077 <= not w26073 and w26076;
w26078 <= not w10992 and w26077;
w26079 <= not w22606 and w26077;
w26080 <= not w26078 and not w26079;
w26081 <= a(2) and not w26080;
w26082 <= not a(2) and w26080;
w26083 <= not w26081 and not w26082;
w26084 <= w26072 and w26083;
w26085 <= w25666 and not w25668;
w26086 <= not w25669 and not w26085;
w26087 <= not w26084 and w26086;
w26088 <= not w26072 and not w26083;
w26089 <= not w26087 and not w26088;
w26090 <= w26041 and not w26089;
w26091 <= not w26041 and w26089;
w26092 <= w11662 and w22325;
w26093 <= w10990 and w22331;
w26094 <= w11650 and w22328;
w26095 <= not w26093 and not w26094;
w26096 <= not w26092 and w26095;
w26097 <= w10992 and w22584;
w26098 <= w26096 and not w26097;
w26099 <= not a(2) and not w26098;
w26100 <= a(2) and w26098;
w26101 <= not w26099 and not w26100;
w26102 <= not w26091 and not w26101;
w26103 <= not w26090 and not w26102;
w26104 <= w11662 and w22322;
w26105 <= w10990 and w22328;
w26106 <= w11650 and w22325;
w26107 <= not w26105 and not w26106;
w26108 <= not w26104 and w26107;
w26109 <= not w10992 and w26108;
w26110 <= not w22517 and w26108;
w26111 <= not w26109 and not w26110;
w26112 <= a(2) and not w26111;
w26113 <= not a(2) and w26111;
w26114 <= not w26112 and not w26113;
w26115 <= not w26103 and not w26114;
w26116 <= w26103 and w26114;
w26117 <= w25685 and w25696;
w26118 <= not w25697 and not w26117;
w26119 <= not w26116 and w26118;
w26120 <= not w26115 and not w26119;
w26121 <= w26039 and not w26120;
w26122 <= not w26039 and w26120;
w26123 <= w11662 and w22319;
w26124 <= w10990 and w22325;
w26125 <= w11650 and w22322;
w26126 <= not w26124 and not w26125;
w26127 <= not w26123 and w26126;
w26128 <= w10992 and w22741;
w26129 <= w26127 and not w26128;
w26130 <= not a(2) and not w26129;
w26131 <= a(2) and w26129;
w26132 <= not w26130 and not w26131;
w26133 <= not w26122 and not w26132;
w26134 <= not w26121 and not w26133;
w26135 <= w11662 and w22315;
w26136 <= w10990 and w22322;
w26137 <= w11650 and w22319;
w26138 <= not w26136 and not w26137;
w26139 <= not w26135 and w26138;
w26140 <= not w10992 and w26139;
w26141 <= not w22785 and w26139;
w26142 <= not w26140 and not w26141;
w26143 <= a(2) and not w26142;
w26144 <= not a(2) and w26142;
w26145 <= not w26143 and not w26144;
w26146 <= w26134 and w26145;
w26147 <= w25643 and w25702;
w26148 <= not w25703 and not w26147;
w26149 <= not w26146 and w26148;
w26150 <= not w26134 and not w26145;
w26151 <= not w26149 and not w26150;
w26152 <= w11662 and w22312;
w26153 <= w10990 and w22319;
w26154 <= w11650 and w22315;
w26155 <= not w26153 and not w26154;
w26156 <= not w26152 and w26155;
w26157 <= not w10992 and w26156;
w26158 <= w22769 and w26156;
w26159 <= not w26157 and not w26158;
w26160 <= a(2) and not w26159;
w26161 <= not a(2) and w26159;
w26162 <= not w26160 and not w26161;
w26163 <= w26151 and w26162;
w26164 <= w25704 and not w25706;
w26165 <= not w25707 and not w26164;
w26166 <= not w26163 and w26165;
w26167 <= not w26151 and not w26162;
w26168 <= not w26166 and not w26167;
w26169 <= w11662 and w22309;
w26170 <= w10990 and w22315;
w26171 <= w11650 and w22312;
w26172 <= not w26170 and not w26171;
w26173 <= not w26169 and w26172;
w26174 <= not w10992 and w26173;
w26175 <= not w22504 and w26173;
w26176 <= not w26174 and not w26175;
w26177 <= a(2) and not w26176;
w26178 <= not a(2) and w26176;
w26179 <= not w26177 and not w26178;
w26180 <= w26168 and w26179;
w26181 <= w25611 and w25708;
w26182 <= not w25709 and not w26181;
w26183 <= not w26180 and w26182;
w26184 <= not w26168 and not w26179;
w26185 <= not w26183 and not w26184;
w26186 <= w25710 and not w25712;
w26187 <= not w25711 and w26186;
w26188 <= not w25714 and not w26187;
w26189 <= not w26185 and w26188;
w26190 <= w26185 and not w26188;
w26191 <= w11662 and w22306;
w26192 <= w10990 and w22312;
w26193 <= w11650 and w22309;
w26194 <= not w26192 and not w26193;
w26195 <= not w26191 and w26194;
w26196 <= w10992 and w22960;
w26197 <= w26195 and not w26196;
w26198 <= not a(2) and not w26197;
w26199 <= a(2) and w26197;
w26200 <= not w26198 and not w26199;
w26201 <= not w26190 and not w26200;
w26202 <= not w26189 and not w26201;
w26203 <= w25715 and not w25717;
w26204 <= not w25716 and w26203;
w26205 <= not w25719 and not w26204;
w26206 <= not w26202 and w26205;
w26207 <= w26202 and not w26205;
w26208 <= w11662 and w22303;
w26209 <= w10990 and w22309;
w26210 <= w11650 and w22306;
w26211 <= not w26209 and not w26210;
w26212 <= not w26208 and w26211;
w26213 <= w10992 and w22941;
w26214 <= w26212 and not w26213;
w26215 <= not a(2) and not w26214;
w26216 <= a(2) and w26214;
w26217 <= not w26215 and not w26216;
w26218 <= not w26207 and not w26217;
w26219 <= not w26206 and not w26218;
w26220 <= w26037 and not w26219;
w26221 <= not w26037 and w26219;
w26222 <= w11662 and w22300;
w26223 <= w10990 and w22306;
w26224 <= w11650 and w22303;
w26225 <= not w26223 and not w26224;
w26226 <= not w26222 and w26225;
w26227 <= w10992 and not w22928;
w26228 <= w26226 and not w26227;
w26229 <= not a(2) and not w26228;
w26230 <= a(2) and w26228;
w26231 <= not w26229 and not w26230;
w26232 <= not w26221 and not w26231;
w26233 <= not w26220 and not w26232;
w26234 <= w11662 and w22297;
w26235 <= w10990 and w22303;
w26236 <= w11650 and w22300;
w26237 <= not w26235 and not w26236;
w26238 <= not w26234 and w26237;
w26239 <= not w10992 and w26238;
w26240 <= w23255 and w26238;
w26241 <= not w26239 and not w26240;
w26242 <= a(2) and not w26241;
w26243 <= not a(2) and w26241;
w26244 <= not w26242 and not w26243;
w26245 <= w26233 and w26244;
w26246 <= w25552 and w25724;
w26247 <= not w25725 and not w26246;
w26248 <= not w26245 and w26247;
w26249 <= not w26233 and not w26244;
w26250 <= not w26248 and not w26249;
w26251 <= w11662 and w22294;
w26252 <= w10990 and w22300;
w26253 <= w11650 and w22297;
w26254 <= not w26252 and not w26253;
w26255 <= not w26251 and w26254;
w26256 <= not w10992 and w26255;
w26257 <= not w23303 and w26255;
w26258 <= not w26256 and not w26257;
w26259 <= a(2) and not w26258;
w26260 <= not a(2) and w26258;
w26261 <= not w26259 and not w26260;
w26262 <= w26250 and w26261;
w26263 <= w25534 and w25726;
w26264 <= not w25727 and not w26263;
w26265 <= not w26262 and w26264;
w26266 <= not w26250 and not w26261;
w26267 <= not w26265 and not w26266;
w26268 <= w11662 and w22291;
w26269 <= w10990 and w22297;
w26270 <= w11650 and w22294;
w26271 <= not w26269 and not w26270;
w26272 <= not w26268 and w26271;
w26273 <= not w10992 and w26272;
w26274 <= w23280 and w26272;
w26275 <= not w26273 and not w26274;
w26276 <= a(2) and not w26275;
w26277 <= not a(2) and w26275;
w26278 <= not w26276 and not w26277;
w26279 <= w26267 and w26278;
w26280 <= w25516 and w25728;
w26281 <= not w25729 and not w26280;
w26282 <= not w26279 and w26281;
w26283 <= not w26267 and not w26278;
w26284 <= not w26282 and not w26283;
w26285 <= w25730 and not w25732;
w26286 <= not w25731 and w26285;
w26287 <= not w25734 and not w26286;
w26288 <= not w26284 and w26287;
w26289 <= w26284 and not w26287;
w26290 <= w11662 and w22288;
w26291 <= w10990 and w22294;
w26292 <= w11650 and w22291;
w26293 <= not w26291 and not w26292;
w26294 <= not w26290 and w26293;
w26295 <= w10992 and not w22491;
w26296 <= w26294 and not w26295;
w26297 <= not a(2) and not w26296;
w26298 <= a(2) and w26296;
w26299 <= not w26297 and not w26298;
w26300 <= not w26289 and not w26299;
w26301 <= not w26288 and not w26300;
w26302 <= w25735 and not w25737;
w26303 <= not w25736 and w26302;
w26304 <= not w25739 and not w26303;
w26305 <= not w26301 and w26304;
w26306 <= w26301 and not w26304;
w26307 <= w11662 and w22285;
w26308 <= w10990 and w22291;
w26309 <= w11650 and w22288;
w26310 <= not w26308 and not w26309;
w26311 <= not w26307 and w26310;
w26312 <= w10992 and w23607;
w26313 <= w26311 and not w26312;
w26314 <= not a(2) and not w26313;
w26315 <= a(2) and w26313;
w26316 <= not w26314 and not w26315;
w26317 <= not w26306 and not w26316;
w26318 <= not w26305 and not w26317;
w26319 <= w26035 and not w26318;
w26320 <= not w26035 and w26318;
w26321 <= w11662 and w22282;
w26322 <= w10990 and w22288;
w26323 <= w11650 and w22285;
w26324 <= not w26322 and not w26323;
w26325 <= not w26321 and w26324;
w26326 <= w10992 and not w23594;
w26327 <= w26325 and not w26326;
w26328 <= not a(2) and not w26327;
w26329 <= a(2) and w26327;
w26330 <= not w26328 and not w26329;
w26331 <= not w26320 and not w26330;
w26332 <= not w26319 and not w26331;
w26333 <= w11662 and w22279;
w26334 <= w10990 and w22285;
w26335 <= w11650 and w22282;
w26336 <= not w26334 and not w26335;
w26337 <= not w26333 and w26336;
w26338 <= not w10992 and w26337;
w26339 <= w23577 and w26337;
w26340 <= not w26338 and not w26339;
w26341 <= a(2) and not w26340;
w26342 <= not a(2) and w26340;
w26343 <= not w26341 and not w26342;
w26344 <= w26332 and w26343;
w26345 <= w25457 and w25744;
w26346 <= not w25745 and not w26345;
w26347 <= not w26344 and w26346;
w26348 <= not w26332 and not w26343;
w26349 <= not w26347 and not w26348;
w26350 <= w11662 and w22276;
w26351 <= w10990 and w22282;
w26352 <= w11650 and w22279;
w26353 <= not w26351 and not w26352;
w26354 <= not w26350 and w26353;
w26355 <= not w10992 and w26354;
w26356 <= not w24077 and w26354;
w26357 <= not w26355 and not w26356;
w26358 <= a(2) and not w26357;
w26359 <= not a(2) and w26357;
w26360 <= not w26358 and not w26359;
w26361 <= w26349 and w26360;
w26362 <= w25439 and w25746;
w26363 <= not w25747 and not w26362;
w26364 <= not w26361 and w26363;
w26365 <= not w26349 and not w26360;
w26366 <= not w26364 and not w26365;
w26367 <= w11662 and w22273;
w26368 <= w10990 and w22279;
w26369 <= w11650 and w22276;
w26370 <= not w26368 and not w26369;
w26371 <= not w26367 and w26370;
w26372 <= not w10992 and w26371;
w26373 <= w24123 and w26371;
w26374 <= not w26372 and not w26373;
w26375 <= a(2) and not w26374;
w26376 <= not a(2) and w26374;
w26377 <= not w26375 and not w26376;
w26378 <= w26366 and w26377;
w26379 <= w25421 and w25748;
w26380 <= not w25749 and not w26379;
w26381 <= not w26378 and w26380;
w26382 <= not w26366 and not w26377;
w26383 <= not w26381 and not w26382;
w26384 <= w25750 and not w25752;
w26385 <= not w25751 and w26384;
w26386 <= not w25754 and not w26385;
w26387 <= not w26383 and w26386;
w26388 <= w26383 and not w26386;
w26389 <= w11662 and w22270;
w26390 <= w10990 and w22276;
w26391 <= w11650 and w22273;
w26392 <= not w26390 and not w26391;
w26393 <= not w26389 and w26392;
w26394 <= w10992 and not w24102;
w26395 <= w26393 and not w26394;
w26396 <= not a(2) and not w26395;
w26397 <= a(2) and w26395;
w26398 <= not w26396 and not w26397;
w26399 <= not w26388 and not w26398;
w26400 <= not w26387 and not w26399;
w26401 <= w25755 and not w25757;
w26402 <= not w25756 and w26401;
w26403 <= not w25759 and not w26402;
w26404 <= not w26400 and w26403;
w26405 <= w26400 and not w26403;
w26406 <= w11662 and w22267;
w26407 <= w10990 and w22273;
w26408 <= w11650 and w22270;
w26409 <= not w26407 and not w26408;
w26410 <= not w26406 and w26409;
w26411 <= w10992 and w22477;
w26412 <= w26410 and not w26411;
w26413 <= not a(2) and not w26412;
w26414 <= a(2) and w26412;
w26415 <= not w26413 and not w26414;
w26416 <= not w26405 and not w26415;
w26417 <= not w26404 and not w26416;
w26418 <= w26033 and not w26417;
w26419 <= not w26033 and w26417;
w26420 <= w11662 and w22264;
w26421 <= w10990 and w22270;
w26422 <= w11650 and w22267;
w26423 <= not w26421 and not w26422;
w26424 <= not w26420 and w26423;
w26425 <= w10992 and not w24568;
w26426 <= w26424 and not w26425;
w26427 <= not a(2) and not w26426;
w26428 <= a(2) and w26426;
w26429 <= not w26427 and not w26428;
w26430 <= not w26419 and not w26429;
w26431 <= not w26418 and not w26430;
w26432 <= w11662 and w22261;
w26433 <= w10990 and w22267;
w26434 <= w11650 and w22264;
w26435 <= not w26433 and not w26434;
w26436 <= not w26432 and w26435;
w26437 <= not w10992 and w26436;
w26438 <= w24551 and w26436;
w26439 <= not w26437 and not w26438;
w26440 <= a(2) and not w26439;
w26441 <= not a(2) and w26439;
w26442 <= not w26440 and not w26441;
w26443 <= w26431 and w26442;
w26444 <= w25362 and w25764;
w26445 <= not w25765 and not w26444;
w26446 <= not w26443 and w26445;
w26447 <= not w26431 and not w26442;
w26448 <= not w26446 and not w26447;
w26449 <= w11662 and w22258;
w26450 <= w10990 and w22264;
w26451 <= w11650 and w22261;
w26452 <= not w26450 and not w26451;
w26453 <= not w26449 and w26452;
w26454 <= not w10992 and w26453;
w26455 <= not w24534 and w26453;
w26456 <= not w26454 and not w26455;
w26457 <= a(2) and not w26456;
w26458 <= not a(2) and w26456;
w26459 <= not w26457 and not w26458;
w26460 <= w26448 and w26459;
w26461 <= w25344 and w25766;
w26462 <= not w25767 and not w26461;
w26463 <= not w26460 and w26462;
w26464 <= not w26448 and not w26459;
w26465 <= not w26463 and not w26464;
w26466 <= w11662 and w22255;
w26467 <= w10990 and w22261;
w26468 <= w11650 and w22258;
w26469 <= not w26467 and not w26468;
w26470 <= not w26466 and w26469;
w26471 <= not w10992 and w26470;
w26472 <= w25205 and w26470;
w26473 <= not w26471 and not w26472;
w26474 <= a(2) and not w26473;
w26475 <= not a(2) and w26473;
w26476 <= not w26474 and not w26475;
w26477 <= w26465 and w26476;
w26478 <= w25326 and w25768;
w26479 <= not w25769 and not w26478;
w26480 <= not w26477 and w26479;
w26481 <= not w26465 and not w26476;
w26482 <= not w26480 and not w26481;
w26483 <= w25770 and not w25772;
w26484 <= not w25771 and w26483;
w26485 <= not w25774 and not w26484;
w26486 <= not w26482 and w26485;
w26487 <= w26482 and not w26485;
w26488 <= w11662 and w22247;
w26489 <= w10990 and w22258;
w26490 <= w11650 and w22255;
w26491 <= not w26489 and not w26490;
w26492 <= not w26488 and w26491;
w26493 <= w10992 and not w25250;
w26494 <= w26492 and not w26493;
w26495 <= not a(2) and not w26494;
w26496 <= a(2) and w26494;
w26497 <= not w26495 and not w26496;
w26498 <= not w26487 and not w26497;
w26499 <= not w26486 and not w26498;
w26500 <= w26031 and not w26499;
w26501 <= not w26031 and w26499;
w26502 <= w11662 and w22250;
w26503 <= w10990 and w22255;
w26504 <= w11650 and w22247;
w26505 <= not w26503 and not w26504;
w26506 <= not w26502 and w26505;
w26507 <= w10992 and w25229;
w26508 <= w26506 and not w26507;
w26509 <= not a(2) and not w26508;
w26510 <= a(2) and w26508;
w26511 <= not w26509 and not w26510;
w26512 <= not w26501 and not w26511;
w26513 <= not w26500 and not w26512;
w26514 <= w11662 and w22244;
w26515 <= w10990 and w22247;
w26516 <= w11650 and w22250;
w26517 <= not w26515 and not w26516;
w26518 <= not w26514 and w26517;
w26519 <= not w10992 and w26518;
w26520 <= w22464 and w26518;
w26521 <= not w26519 and not w26520;
w26522 <= a(2) and not w26521;
w26523 <= not a(2) and w26521;
w26524 <= not w26522 and not w26523;
w26525 <= w26513 and w26524;
w26526 <= w25281 and w25779;
w26527 <= not w25780 and not w26526;
w26528 <= not w26525 and w26527;
w26529 <= not w26513 and not w26524;
w26530 <= not w26528 and not w26529;
w26531 <= w11662 and w25998;
w26532 <= w10990 and w22250;
w26533 <= w11650 and w22244;
w26534 <= not w26532 and not w26533;
w26535 <= not w26531 and w26534;
w26536 <= not w10992 and w26535;
w26537 <= not w22462 and not w26010;
w26538 <= not w26008 and w26011;
w26539 <= not w26537 and not w26538;
w26540 <= w26535 and w26539;
w26541 <= not w26536 and not w26540;
w26542 <= a(2) and not w26541;
w26543 <= not a(2) and w26541;
w26544 <= not w26542 and not w26543;
w26545 <= w26530 and w26544;
w26546 <= w25263 and w25781;
w26547 <= not w25782 and not w26546;
w26548 <= not w26545 and w26547;
w26549 <= not w26530 and not w26544;
w26550 <= not w26548 and not w26549;
w26551 <= w11662 and w26001;
w26552 <= w10990 and w22244;
w26553 <= w11650 and w25998;
w26554 <= not w26552 and not w26553;
w26555 <= not w26551 and w26554;
w26556 <= not w10992 and w26555;
w26557 <= not w26011 and not w26014;
w26558 <= not w26012 and w26015;
w26559 <= not w26557 and not w26558;
w26560 <= w26555 and w26559;
w26561 <= not w26556 and not w26560;
w26562 <= a(2) and not w26561;
w26563 <= not a(2) and w26561;
w26564 <= not w26562 and not w26563;
w26565 <= w26550 and w26564;
w26566 <= w25242 and w25783;
w26567 <= not w25784 and not w26566;
w26568 <= not w26565 and w26567;
w26569 <= not w26550 and not w26564;
w26570 <= not w26568 and not w26569;
w26571 <= w25788 and not w26029;
w26572 <= not w26028 and not w26029;
w26573 <= not w26571 and not w26572;
w26574 <= not w26570 and not w26573;
w26575 <= not w26029 and not w26574;
w26576 <= w6 and w25998;
w26577 <= w9802 and w22250;
w26578 <= w10369 and w22244;
w26579 <= not w26577 and not w26578;
w26580 <= not w26576 and w26579;
w26581 <= w9805 and not w26539;
w26582 <= w26580 and not w26581;
w26583 <= a(5) and not w26582;
w26584 <= not w26582 and not w26583;
w26585 <= a(5) and not w26583;
w26586 <= not w26584 and not w26585;
w26587 <= not w25211 and not w25215;
w26588 <= w7918 and w22261;
w26589 <= w7226 and w22267;
w26590 <= w7567 and w22264;
w26591 <= not w26589 and not w26590;
w26592 <= not w26588 and w26591;
w26593 <= w7229 and not w24551;
w26594 <= w26592 and not w26593;
w26595 <= a(11) and not w26594;
w26596 <= not w26594 and not w26595;
w26597 <= a(11) and not w26595;
w26598 <= not w26596 and not w26597;
w26599 <= not w25181 and not w25185;
w26600 <= w6168 and w22279;
w26601 <= w5598 and w22285;
w26602 <= w5874 and w22282;
w26603 <= not w26601 and not w26602;
w26604 <= not w26600 and w26603;
w26605 <= w5601 and not w23577;
w26606 <= w26604 and not w26605;
w26607 <= a(17) and not w26606;
w26608 <= not w26606 and not w26607;
w26609 <= a(17) and not w26607;
w26610 <= not w26608 and not w26609;
w26611 <= not w25154 and not w25158;
w26612 <= w4629 and w22297;
w26613 <= w4468 and w22303;
w26614 <= w4539 and w22300;
w26615 <= not w26613 and not w26614;
w26616 <= not w26612 and w26615;
w26617 <= w4471 and not w23255;
w26618 <= w26616 and not w26617;
w26619 <= a(23) and not w26618;
w26620 <= not w26618 and not w26619;
w26621 <= a(23) and not w26619;
w26622 <= not w26620 and not w26621;
w26623 <= not w25127 and not w25131;
w26624 <= w3392 and w22315;
w26625 <= w3477 and w22322;
w26626 <= w3541 and w22319;
w26627 <= not w26625 and not w26626;
w26628 <= not w26624 and w26627;
w26629 <= w3303 and w22785;
w26630 <= w26628 and not w26629;
w26631 <= a(29) and not w26630;
w26632 <= not w26630 and not w26631;
w26633 <= a(29) and not w26631;
w26634 <= not w26632 and not w26633;
w26635 <= not w25100 and not w25104;
w26636 <= w12332 and w13724;
w26637 <= w4706 and w26636;
w26638 <= w1822 and w26637;
w26639 <= w725 and w26638;
w26640 <= w13612 and w26639;
w26641 <= w4246 and w26640;
w26642 <= w3090 and w26641;
w26643 <= w179 and w26642;
w26644 <= w868 and w26643;
w26645 <= w1172 and w26644;
w26646 <= w51 and w26645;
w26647 <= not w1036 and w26646;
w26648 <= not w357 and w26647;
w26649 <= not w428 and w26648;
w26650 <= not w363 and w26649;
w26651 <= w2955 and w22325;
w26652 <= w2963 and w22328;
w26653 <= w2958 and w22331;
w26654 <= w10 and w22584;
w26655 <= not w26653 and not w26654;
w26656 <= not w26652 and w26655;
w26657 <= not w26651 and w26656;
w26658 <= not w26650 and not w26657;
w26659 <= not w26650 and not w26658;
w26660 <= not w26657 and not w26658;
w26661 <= not w26659 and not w26660;
w26662 <= not w26635 and not w26661;
w26663 <= not w26635 and not w26662;
w26664 <= not w26661 and not w26662;
w26665 <= not w26663 and not w26664;
w26666 <= not w26634 and not w26665;
w26667 <= not w26634 and not w26666;
w26668 <= not w26665 and not w26666;
w26669 <= not w26667 and not w26668;
w26670 <= not w25108 and not w25114;
w26671 <= w26669 and w26670;
w26672 <= not w26669 and not w26670;
w26673 <= not w26671 and not w26672;
w26674 <= w3819 and w22306;
w26675 <= w3902 and w22312;
w26676 <= w3981 and w22309;
w26677 <= not w26675 and not w26676;
w26678 <= not w26674 and w26677;
w26679 <= not w3985 and w26678;
w26680 <= not w22960 and w26678;
w26681 <= not w26679 and not w26680;
w26682 <= a(26) and not w26681;
w26683 <= not a(26) and w26681;
w26684 <= not w26682 and not w26683;
w26685 <= w26673 and not w26684;
w26686 <= w26673 and not w26685;
w26687 <= not w26684 and not w26685;
w26688 <= not w26686 and not w26687;
w26689 <= not w26623 and not w26688;
w26690 <= not w26623 and not w26689;
w26691 <= not w26688 and not w26689;
w26692 <= not w26690 and not w26691;
w26693 <= not w26622 and not w26692;
w26694 <= not w26622 and not w26693;
w26695 <= not w26692 and not w26693;
w26696 <= not w26694 and not w26695;
w26697 <= not w25135 and not w25141;
w26698 <= w26696 and w26697;
w26699 <= not w26696 and not w26697;
w26700 <= not w26698 and not w26699;
w26701 <= w5431 and w22288;
w26702 <= w4870 and w22294;
w26703 <= w5342 and w22291;
w26704 <= not w26702 and not w26703;
w26705 <= not w26701 and w26704;
w26706 <= not w4873 and w26705;
w26707 <= w22491 and w26705;
w26708 <= not w26706 and not w26707;
w26709 <= a(20) and not w26708;
w26710 <= not a(20) and w26708;
w26711 <= not w26709 and not w26710;
w26712 <= w26700 and not w26711;
w26713 <= w26700 and not w26712;
w26714 <= not w26711 and not w26712;
w26715 <= not w26713 and not w26714;
w26716 <= not w26611 and not w26715;
w26717 <= not w26611 and not w26716;
w26718 <= not w26715 and not w26716;
w26719 <= not w26717 and not w26718;
w26720 <= not w26610 and not w26719;
w26721 <= not w26610 and not w26720;
w26722 <= not w26719 and not w26720;
w26723 <= not w26721 and not w26722;
w26724 <= not w25162 and not w25168;
w26725 <= w26723 and w26724;
w26726 <= not w26723 and not w26724;
w26727 <= not w26725 and not w26726;
w26728 <= w7036 and w22270;
w26729 <= w6337 and w22276;
w26730 <= w6886 and w22273;
w26731 <= not w26729 and not w26730;
w26732 <= not w26728 and w26731;
w26733 <= not w6332 and w26732;
w26734 <= w24102 and w26732;
w26735 <= not w26733 and not w26734;
w26736 <= a(14) and not w26735;
w26737 <= not a(14) and w26735;
w26738 <= not w26736 and not w26737;
w26739 <= w26727 and not w26738;
w26740 <= w26727 and not w26739;
w26741 <= not w26738 and not w26739;
w26742 <= not w26740 and not w26741;
w26743 <= not w26599 and not w26742;
w26744 <= not w26599 and not w26743;
w26745 <= not w26742 and not w26743;
w26746 <= not w26744 and not w26745;
w26747 <= not w26598 and not w26746;
w26748 <= not w26598 and not w26747;
w26749 <= not w26746 and not w26747;
w26750 <= not w26748 and not w26749;
w26751 <= not w25189 and not w25195;
w26752 <= w26750 and w26751;
w26753 <= not w26750 and not w26751;
w26754 <= not w26752 and not w26753;
w26755 <= w9266 and w22247;
w26756 <= w8353 and w22258;
w26757 <= w8795 and w22255;
w26758 <= not w26756 and not w26757;
w26759 <= not w26755 and w26758;
w26760 <= not w8356 and w26759;
w26761 <= w25250 and w26759;
w26762 <= not w26760 and not w26761;
w26763 <= a(8) and not w26762;
w26764 <= not a(8) and w26762;
w26765 <= not w26763 and not w26764;
w26766 <= w26754 and not w26765;
w26767 <= w26754 and not w26766;
w26768 <= not w26765 and not w26766;
w26769 <= not w26767 and not w26768;
w26770 <= not w26587 and not w26769;
w26771 <= not w26587 and not w26770;
w26772 <= not w26769 and not w26770;
w26773 <= not w26771 and not w26772;
w26774 <= not w26586 and not w26773;
w26775 <= not w26586 and not w26774;
w26776 <= not w26773 and not w26774;
w26777 <= not w26775 and not w26776;
w26778 <= not w25219 and not w25787;
w26779 <= w26777 and w26778;
w26780 <= not w26777 and not w26778;
w26781 <= not w26779 and not w26780;
w26782 <= not w25990 and not w25994;
w26783 <= not w25981 and not w25987;
w26784 <= w10 and w13864;
w26785 <= w2955 and w13568;
w26786 <= w2958 and w13532;
w26787 <= w2963 and w13565;
w26788 <= not w26786 and not w26787;
w26789 <= not w26785 and w26788;
w26790 <= not w26784 and w26789;
w26791 <= not w25958 and not w25960;
w26792 <= w3965 and w4446;
w26793 <= w25951 and w26792;
w26794 <= not w263 and w26793;
w26795 <= not w26791 and w26794;
w26796 <= w26791 and not w26794;
w26797 <= not w26795 and not w26796;
w26798 <= not w26790 and w26797;
w26799 <= not w26790 and not w26798;
w26800 <= w26797 and not w26798;
w26801 <= not w26799 and not w26800;
w26802 <= not w25963 and not w25966;
w26803 <= w26801 and w26802;
w26804 <= not w26801 and not w26802;
w26805 <= not w26803 and not w26804;
w26806 <= w3392 and not w13373;
w26807 <= w3477 and not w13562;
w26808 <= w3541 and w13876;
w26809 <= not w26807 and not w26808;
w26810 <= not w26806 and w26809;
w26811 <= not w3303 and w26810;
w26812 <= not w13963 and w26810;
w26813 <= not w26811 and not w26812;
w26814 <= a(29) and not w26813;
w26815 <= not a(29) and w26813;
w26816 <= not w26814 and not w26815;
w26817 <= w26805 and not w26816;
w26818 <= not w26805 and w26816;
w26819 <= not w26817 and not w26818;
w26820 <= not w26783 and w26819;
w26821 <= w26783 and not w26819;
w26822 <= not w26820 and not w26821;
w26823 <= not w26782 and w26822;
w26824 <= w26782 and not w26822;
w26825 <= not w26823 and not w26824;
w26826 <= w11662 and w26825;
w26827 <= w10990 and w26001;
w26828 <= w11650 and w25995;
w26829 <= not w26827 and not w26828;
w26830 <= not w26826 and w26829;
w26831 <= not w10992 and w26830;
w26832 <= w25995 and w26825;
w26833 <= not w25995 and not w26825;
w26834 <= not w26021 and not w26833;
w26835 <= not w26832 and w26834;
w26836 <= not w26021 and not w26835;
w26837 <= not w26832 and not w26835;
w26838 <= not w26833 and w26837;
w26839 <= not w26836 and not w26838;
w26840 <= w26830 and w26839;
w26841 <= not w26831 and not w26840;
w26842 <= a(2) and not w26841;
w26843 <= not a(2) and w26841;
w26844 <= not w26842 and not w26843;
w26845 <= w26781 and not w26844;
w26846 <= not w26781 and w26844;
w26847 <= not w26845 and not w26846;
w26848 <= not w26575 and w26847;
w26849 <= w26575 and not w26847;
w26850 <= not w26848 and not w26849;
w26851 <= not w26570 and not w26574;
w26852 <= not w26573 and not w26574;
w26853 <= not w26851 and not w26852;
w26854 <= w26850 and w26853;
w26855 <= not w26850 and not w26853;
w26856 <= not w26854 and not w26855;
w26857 <= w26850 and not w26853;
w26858 <= not w26845 and not w26848;
w26859 <= w6 and w26001;
w26860 <= w9802 and w22244;
w26861 <= w10369 and w25998;
w26862 <= not w26860 and not w26861;
w26863 <= not w26859 and w26862;
w26864 <= w9805 and not w26559;
w26865 <= w26863 and not w26864;
w26866 <= a(5) and not w26865;
w26867 <= not w26865 and not w26866;
w26868 <= a(5) and not w26866;
w26869 <= not w26867 and not w26868;
w26870 <= not w26766 and not w26770;
w26871 <= w7918 and w22258;
w26872 <= w7226 and w22264;
w26873 <= w7567 and w22261;
w26874 <= not w26872 and not w26873;
w26875 <= not w26871 and w26874;
w26876 <= w7229 and w24534;
w26877 <= w26875 and not w26876;
w26878 <= a(11) and not w26877;
w26879 <= not w26877 and not w26878;
w26880 <= a(11) and not w26878;
w26881 <= not w26879 and not w26880;
w26882 <= not w26739 and not w26743;
w26883 <= w6168 and w22276;
w26884 <= w5598 and w22282;
w26885 <= w5874 and w22279;
w26886 <= not w26884 and not w26885;
w26887 <= not w26883 and w26886;
w26888 <= w5601 and w24077;
w26889 <= w26887 and not w26888;
w26890 <= a(17) and not w26889;
w26891 <= not w26889 and not w26890;
w26892 <= a(17) and not w26890;
w26893 <= not w26891 and not w26892;
w26894 <= not w26712 and not w26716;
w26895 <= w4629 and w22294;
w26896 <= w4468 and w22300;
w26897 <= w4539 and w22297;
w26898 <= not w26896 and not w26897;
w26899 <= not w26895 and w26898;
w26900 <= w4471 and w23303;
w26901 <= w26899 and not w26900;
w26902 <= a(23) and not w26901;
w26903 <= not w26901 and not w26902;
w26904 <= a(23) and not w26902;
w26905 <= not w26903 and not w26904;
w26906 <= not w26685 and not w26689;
w26907 <= not w26666 and not w26672;
w26908 <= not w26658 and not w26662;
w26909 <= w1538 and w3449;
w26910 <= w1960 and w26909;
w26911 <= w6563 and w26910;
w26912 <= w14479 and w26911;
w26913 <= w6690 and w26912;
w26914 <= w2914 and w26913;
w26915 <= w3479 and w26914;
w26916 <= w1510 and w26915;
w26917 <= w2518 and w26916;
w26918 <= w1172 and w26917;
w26919 <= w2340 and w26918;
w26920 <= w1457 and w26919;
w26921 <= not w1181 and w26920;
w26922 <= not w265 and w26921;
w26923 <= not w231 and w26922;
w26924 <= not w307 and w26923;
w26925 <= not w867 and w26924;
w26926 <= not w706 and w26925;
w26927 <= w2955 and w22322;
w26928 <= w2963 and w22325;
w26929 <= w2958 and w22328;
w26930 <= w10 and w22517;
w26931 <= not w26929 and not w26930;
w26932 <= not w26928 and w26931;
w26933 <= not w26927 and w26932;
w26934 <= not w26926 and not w26933;
w26935 <= not w26926 and not w26934;
w26936 <= not w26933 and not w26934;
w26937 <= not w26935 and not w26936;
w26938 <= not w26908 and not w26937;
w26939 <= not w26908 and not w26938;
w26940 <= not w26937 and not w26938;
w26941 <= not w26939 and not w26940;
w26942 <= w3392 and w22312;
w26943 <= w3477 and w22319;
w26944 <= w3541 and w22315;
w26945 <= not w26943 and not w26944;
w26946 <= not w26942 and w26945;
w26947 <= not w3303 and w26946;
w26948 <= w22769 and w26946;
w26949 <= not w26947 and not w26948;
w26950 <= a(29) and not w26949;
w26951 <= not a(29) and w26949;
w26952 <= not w26950 and not w26951;
w26953 <= not w26941 and not w26952;
w26954 <= w26941 and w26952;
w26955 <= not w26953 and not w26954;
w26956 <= not w26907 and w26955;
w26957 <= w26907 and not w26955;
w26958 <= not w26956 and not w26957;
w26959 <= w3819 and w22303;
w26960 <= w3902 and w22309;
w26961 <= w3981 and w22306;
w26962 <= not w26960 and not w26961;
w26963 <= not w26959 and w26962;
w26964 <= not w3985 and w26963;
w26965 <= not w22941 and w26963;
w26966 <= not w26964 and not w26965;
w26967 <= a(26) and not w26966;
w26968 <= not a(26) and w26966;
w26969 <= not w26967 and not w26968;
w26970 <= w26958 and not w26969;
w26971 <= w26958 and not w26970;
w26972 <= not w26969 and not w26970;
w26973 <= not w26971 and not w26972;
w26974 <= not w26906 and not w26973;
w26975 <= not w26906 and not w26974;
w26976 <= not w26973 and not w26974;
w26977 <= not w26975 and not w26976;
w26978 <= not w26905 and not w26977;
w26979 <= not w26905 and not w26978;
w26980 <= not w26977 and not w26978;
w26981 <= not w26979 and not w26980;
w26982 <= not w26693 and not w26699;
w26983 <= w26981 and w26982;
w26984 <= not w26981 and not w26982;
w26985 <= not w26983 and not w26984;
w26986 <= w5431 and w22285;
w26987 <= w4870 and w22291;
w26988 <= w5342 and w22288;
w26989 <= not w26987 and not w26988;
w26990 <= not w26986 and w26989;
w26991 <= not w4873 and w26990;
w26992 <= not w23607 and w26990;
w26993 <= not w26991 and not w26992;
w26994 <= a(20) and not w26993;
w26995 <= not a(20) and w26993;
w26996 <= not w26994 and not w26995;
w26997 <= w26985 and not w26996;
w26998 <= w26985 and not w26997;
w26999 <= not w26996 and not w26997;
w27000 <= not w26998 and not w26999;
w27001 <= not w26894 and not w27000;
w27002 <= not w26894 and not w27001;
w27003 <= not w27000 and not w27001;
w27004 <= not w27002 and not w27003;
w27005 <= not w26893 and not w27004;
w27006 <= not w26893 and not w27005;
w27007 <= not w27004 and not w27005;
w27008 <= not w27006 and not w27007;
w27009 <= not w26720 and not w26726;
w27010 <= w27008 and w27009;
w27011 <= not w27008 and not w27009;
w27012 <= not w27010 and not w27011;
w27013 <= w7036 and w22267;
w27014 <= w6337 and w22273;
w27015 <= w6886 and w22270;
w27016 <= not w27014 and not w27015;
w27017 <= not w27013 and w27016;
w27018 <= not w6332 and w27017;
w27019 <= not w22477 and w27017;
w27020 <= not w27018 and not w27019;
w27021 <= a(14) and not w27020;
w27022 <= not a(14) and w27020;
w27023 <= not w27021 and not w27022;
w27024 <= w27012 and not w27023;
w27025 <= w27012 and not w27024;
w27026 <= not w27023 and not w27024;
w27027 <= not w27025 and not w27026;
w27028 <= not w26882 and not w27027;
w27029 <= not w26882 and not w27028;
w27030 <= not w27027 and not w27028;
w27031 <= not w27029 and not w27030;
w27032 <= not w26881 and not w27031;
w27033 <= not w26881 and not w27032;
w27034 <= not w27031 and not w27032;
w27035 <= not w27033 and not w27034;
w27036 <= not w26747 and not w26753;
w27037 <= w27035 and w27036;
w27038 <= not w27035 and not w27036;
w27039 <= not w27037 and not w27038;
w27040 <= w9266 and w22250;
w27041 <= w8353 and w22255;
w27042 <= w8795 and w22247;
w27043 <= not w27041 and not w27042;
w27044 <= not w27040 and w27043;
w27045 <= not w8356 and w27044;
w27046 <= not w25229 and w27044;
w27047 <= not w27045 and not w27046;
w27048 <= a(8) and not w27047;
w27049 <= not a(8) and w27047;
w27050 <= not w27048 and not w27049;
w27051 <= w27039 and not w27050;
w27052 <= w27039 and not w27051;
w27053 <= not w27050 and not w27051;
w27054 <= not w27052 and not w27053;
w27055 <= not w26870 and not w27054;
w27056 <= not w26870 and not w27055;
w27057 <= not w27054 and not w27055;
w27058 <= not w27056 and not w27057;
w27059 <= not w26869 and not w27058;
w27060 <= not w26869 and not w27059;
w27061 <= not w27058 and not w27059;
w27062 <= not w27060 and not w27061;
w27063 <= not w26774 and not w26780;
w27064 <= w27062 and w27063;
w27065 <= not w27062 and not w27063;
w27066 <= not w27064 and not w27065;
w27067 <= not w26820 and not w26823;
w27068 <= not w26804 and not w26817;
w27069 <= not w26795 and not w26798;
w27070 <= w3791 and w4449;
w27071 <= w26794 and not w27070;
w27072 <= not w26794 and w27070;
w27073 <= not w27069 and not w27072;
w27074 <= not w27071 and w27073;
w27075 <= not w27069 and not w27074;
w27076 <= not w27072 and not w27074;
w27077 <= not w27071 and w27076;
w27078 <= not w27075 and not w27077;
w27079 <= not w3392 and not w3541;
w27080 <= not w13373 and not w27079;
w27081 <= w3477 and w13876;
w27082 <= not w27080 and not w27081;
w27083 <= w3303 and not w13886;
w27084 <= w27082 and not w27083;
w27085 <= a(29) and not w27084;
w27086 <= not w27084 and not w27085;
w27087 <= a(29) and not w27085;
w27088 <= not w27086 and not w27087;
w27089 <= w10 and not w13589;
w27090 <= w2955 and not w13562;
w27091 <= w2958 and w13565;
w27092 <= w2963 and w13568;
w27093 <= not w27091 and not w27092;
w27094 <= not w27090 and w27093;
w27095 <= not w27089 and w27094;
w27096 <= not w27088 and not w27095;
w27097 <= not w27088 and not w27096;
w27098 <= not w27095 and not w27096;
w27099 <= not w27097 and not w27098;
w27100 <= not w27078 and w27099;
w27101 <= w27078 and not w27099;
w27102 <= not w27100 and not w27101;
w27103 <= not w27068 and not w27102;
w27104 <= w27068 and w27102;
w27105 <= not w27103 and not w27104;
w27106 <= not w27067 and w27105;
w27107 <= w27067 and not w27105;
w27108 <= not w27106 and not w27107;
w27109 <= w11662 and w27108;
w27110 <= w10990 and w25995;
w27111 <= w11650 and w26825;
w27112 <= not w27110 and not w27111;
w27113 <= not w27109 and w27112;
w27114 <= not w10992 and w27113;
w27115 <= not w26825 and not w27108;
w27116 <= w26825 and w27108;
w27117 <= not w27115 and not w27116;
w27118 <= not w26837 and w27117;
w27119 <= w26837 and not w27117;
w27120 <= not w27118 and not w27119;
w27121 <= w27113 and not w27120;
w27122 <= not w27114 and not w27121;
w27123 <= a(2) and not w27122;
w27124 <= not a(2) and w27122;
w27125 <= not w27123 and not w27124;
w27126 <= w27066 and not w27125;
w27127 <= not w27066 and w27125;
w27128 <= not w27126 and not w27127;
w27129 <= not w26858 and w27128;
w27130 <= w26858 and not w27128;
w27131 <= not w27129 and not w27130;
w27132 <= w26857 and w27131;
w27133 <= not w26857 and not w27131;
w27134 <= not w27132 and not w27133;
w27135 <= not w27126 and not w27129;
w27136 <= w6 and w25995;
w27137 <= w9802 and w25998;
w27138 <= w10369 and w26001;
w27139 <= not w27137 and not w27138;
w27140 <= not w27136 and w27139;
w27141 <= w9805 and not w26023;
w27142 <= w27140 and not w27141;
w27143 <= a(5) and not w27142;
w27144 <= not w27142 and not w27143;
w27145 <= a(5) and not w27143;
w27146 <= not w27144 and not w27145;
w27147 <= not w27051 and not w27055;
w27148 <= w7918 and w22255;
w27149 <= w7226 and w22261;
w27150 <= w7567 and w22258;
w27151 <= not w27149 and not w27150;
w27152 <= not w27148 and w27151;
w27153 <= w7229 and not w25205;
w27154 <= w27152 and not w27153;
w27155 <= a(11) and not w27154;
w27156 <= not w27154 and not w27155;
w27157 <= a(11) and not w27155;
w27158 <= not w27156 and not w27157;
w27159 <= not w27024 and not w27028;
w27160 <= w6168 and w22273;
w27161 <= w5598 and w22279;
w27162 <= w5874 and w22276;
w27163 <= not w27161 and not w27162;
w27164 <= not w27160 and w27163;
w27165 <= w5601 and not w24123;
w27166 <= w27164 and not w27165;
w27167 <= a(17) and not w27166;
w27168 <= not w27166 and not w27167;
w27169 <= a(17) and not w27167;
w27170 <= not w27168 and not w27169;
w27171 <= not w26997 and not w27001;
w27172 <= w4629 and w22291;
w27173 <= w4468 and w22297;
w27174 <= w4539 and w22294;
w27175 <= not w27173 and not w27174;
w27176 <= not w27172 and w27175;
w27177 <= w4471 and not w23280;
w27178 <= w27176 and not w27177;
w27179 <= a(23) and not w27178;
w27180 <= not w27178 and not w27179;
w27181 <= a(23) and not w27179;
w27182 <= not w27180 and not w27181;
w27183 <= not w26970 and not w26974;
w27184 <= not w26953 and not w26956;
w27185 <= not w26934 and not w26938;
w27186 <= w13762 and w14496;
w27187 <= w6652 and w27186;
w27188 <= w2345 and w27187;
w27189 <= w551 and w27188;
w27190 <= w3115 and w27189;
w27191 <= w3126 and w27190;
w27192 <= w1535 and w27191;
w27193 <= w1414 and w27192;
w27194 <= w1779 and w27193;
w27195 <= w450 and w27194;
w27196 <= w1661 and w27195;
w27197 <= w1204 and w27196;
w27198 <= not w42 and w27197;
w27199 <= not w425 and w27198;
w27200 <= not w221 and w27199;
w27201 <= not w180 and w27200;
w27202 <= not w405 and w27201;
w27203 <= w2955 and w22319;
w27204 <= w2963 and w22322;
w27205 <= w2958 and w22325;
w27206 <= w10 and w22741;
w27207 <= not w27205 and not w27206;
w27208 <= not w27204 and w27207;
w27209 <= not w27203 and w27208;
w27210 <= not w27202 and not w27209;
w27211 <= not w27202 and not w27210;
w27212 <= not w27209 and not w27210;
w27213 <= not w27211 and not w27212;
w27214 <= not w27185 and not w27213;
w27215 <= not w27185 and not w27214;
w27216 <= not w27213 and not w27214;
w27217 <= not w27215 and not w27216;
w27218 <= w3392 and w22309;
w27219 <= w3477 and w22315;
w27220 <= w3541 and w22312;
w27221 <= not w27219 and not w27220;
w27222 <= not w27218 and w27221;
w27223 <= not w3303 and w27222;
w27224 <= not w22504 and w27222;
w27225 <= not w27223 and not w27224;
w27226 <= a(29) and not w27225;
w27227 <= not a(29) and w27225;
w27228 <= not w27226 and not w27227;
w27229 <= not w27217 and not w27228;
w27230 <= w27217 and w27228;
w27231 <= not w27229 and not w27230;
w27232 <= not w27184 and w27231;
w27233 <= w27184 and not w27231;
w27234 <= not w27232 and not w27233;
w27235 <= w3819 and w22300;
w27236 <= w3902 and w22306;
w27237 <= w3981 and w22303;
w27238 <= not w27236 and not w27237;
w27239 <= not w27235 and w27238;
w27240 <= not w3985 and w27239;
w27241 <= w22928 and w27239;
w27242 <= not w27240 and not w27241;
w27243 <= a(26) and not w27242;
w27244 <= not a(26) and w27242;
w27245 <= not w27243 and not w27244;
w27246 <= w27234 and not w27245;
w27247 <= w27234 and not w27246;
w27248 <= not w27245 and not w27246;
w27249 <= not w27247 and not w27248;
w27250 <= not w27183 and not w27249;
w27251 <= not w27183 and not w27250;
w27252 <= not w27249 and not w27250;
w27253 <= not w27251 and not w27252;
w27254 <= not w27182 and not w27253;
w27255 <= not w27182 and not w27254;
w27256 <= not w27253 and not w27254;
w27257 <= not w27255 and not w27256;
w27258 <= not w26978 and not w26984;
w27259 <= w27257 and w27258;
w27260 <= not w27257 and not w27258;
w27261 <= not w27259 and not w27260;
w27262 <= w5431 and w22282;
w27263 <= w4870 and w22288;
w27264 <= w5342 and w22285;
w27265 <= not w27263 and not w27264;
w27266 <= not w27262 and w27265;
w27267 <= not w4873 and w27266;
w27268 <= w23594 and w27266;
w27269 <= not w27267 and not w27268;
w27270 <= a(20) and not w27269;
w27271 <= not a(20) and w27269;
w27272 <= not w27270 and not w27271;
w27273 <= w27261 and not w27272;
w27274 <= w27261 and not w27273;
w27275 <= not w27272 and not w27273;
w27276 <= not w27274 and not w27275;
w27277 <= not w27171 and not w27276;
w27278 <= not w27171 and not w27277;
w27279 <= not w27276 and not w27277;
w27280 <= not w27278 and not w27279;
w27281 <= not w27170 and not w27280;
w27282 <= not w27170 and not w27281;
w27283 <= not w27280 and not w27281;
w27284 <= not w27282 and not w27283;
w27285 <= not w27005 and not w27011;
w27286 <= w27284 and w27285;
w27287 <= not w27284 and not w27285;
w27288 <= not w27286 and not w27287;
w27289 <= w7036 and w22264;
w27290 <= w6337 and w22270;
w27291 <= w6886 and w22267;
w27292 <= not w27290 and not w27291;
w27293 <= not w27289 and w27292;
w27294 <= not w6332 and w27293;
w27295 <= w24568 and w27293;
w27296 <= not w27294 and not w27295;
w27297 <= a(14) and not w27296;
w27298 <= not a(14) and w27296;
w27299 <= not w27297 and not w27298;
w27300 <= w27288 and not w27299;
w27301 <= w27288 and not w27300;
w27302 <= not w27299 and not w27300;
w27303 <= not w27301 and not w27302;
w27304 <= not w27159 and not w27303;
w27305 <= not w27159 and not w27304;
w27306 <= not w27303 and not w27304;
w27307 <= not w27305 and not w27306;
w27308 <= not w27158 and not w27307;
w27309 <= not w27158 and not w27308;
w27310 <= not w27307 and not w27308;
w27311 <= not w27309 and not w27310;
w27312 <= not w27032 and not w27038;
w27313 <= w27311 and w27312;
w27314 <= not w27311 and not w27312;
w27315 <= not w27313 and not w27314;
w27316 <= w9266 and w22244;
w27317 <= w8353 and w22247;
w27318 <= w8795 and w22250;
w27319 <= not w27317 and not w27318;
w27320 <= not w27316 and w27319;
w27321 <= not w8356 and w27320;
w27322 <= w22464 and w27320;
w27323 <= not w27321 and not w27322;
w27324 <= a(8) and not w27323;
w27325 <= not a(8) and w27323;
w27326 <= not w27324 and not w27325;
w27327 <= w27315 and not w27326;
w27328 <= w27315 and not w27327;
w27329 <= not w27326 and not w27327;
w27330 <= not w27328 and not w27329;
w27331 <= not w27147 and not w27330;
w27332 <= not w27147 and not w27331;
w27333 <= not w27330 and not w27331;
w27334 <= not w27332 and not w27333;
w27335 <= not w27146 and not w27334;
w27336 <= not w27146 and not w27335;
w27337 <= not w27334 and not w27335;
w27338 <= not w27336 and not w27337;
w27339 <= not w27059 and not w27065;
w27340 <= w27338 and w27339;
w27341 <= not w27338 and not w27339;
w27342 <= not w27340 and not w27341;
w27343 <= not w27103 and not w27106;
w27344 <= not w27078 and not w27099;
w27345 <= not w27096 and not w27344;
w27346 <= w10 and w14071;
w27347 <= w2955 and w13876;
w27348 <= w2958 and w13568;
w27349 <= w2963 and not w13562;
w27350 <= not w27348 and not w27349;
w27351 <= not w27347 and w27350;
w27352 <= not w27346 and w27351;
w27353 <= not w3477 and not w3541;
w27354 <= w3302 and w27353;
w27355 <= not w13373 and not w27354;
w27356 <= a(29) and not w27355;
w27357 <= not a(29) and w27355;
w27358 <= not w27356 and not w27357;
w27359 <= w12991 and w27070;
w27360 <= not w12991 and not w27070;
w27361 <= not w27359 and not w27360;
w27362 <= w27358 and w27361;
w27363 <= not w27358 and not w27361;
w27364 <= not w27362 and not w27363;
w27365 <= not w27352 and w27364;
w27366 <= w27364 and not w27365;
w27367 <= not w27352 and not w27365;
w27368 <= not w27366 and not w27367;
w27369 <= not w27076 and not w27368;
w27370 <= w27076 and w27368;
w27371 <= not w27369 and not w27370;
w27372 <= not w27345 and w27371;
w27373 <= w27345 and not w27371;
w27374 <= not w27372 and not w27373;
w27375 <= not w27343 and w27374;
w27376 <= w27343 and not w27374;
w27377 <= not w27375 and not w27376;
w27378 <= w11662 and w27377;
w27379 <= w10990 and w26825;
w27380 <= w11650 and w27108;
w27381 <= not w27379 and not w27380;
w27382 <= not w27378 and w27381;
w27383 <= not w10992 and w27382;
w27384 <= not w27116 and not w27118;
w27385 <= not w27108 and not w27377;
w27386 <= w27108 and w27377;
w27387 <= not w27385 and not w27386;
w27388 <= not w27384 and w27387;
w27389 <= w27384 and not w27387;
w27390 <= not w27388 and not w27389;
w27391 <= w27382 and not w27390;
w27392 <= not w27383 and not w27391;
w27393 <= a(2) and not w27392;
w27394 <= not a(2) and w27392;
w27395 <= not w27393 and not w27394;
w27396 <= w27342 and not w27395;
w27397 <= not w27342 and w27395;
w27398 <= not w27396 and not w27397;
w27399 <= not w27135 and w27398;
w27400 <= w27135 and not w27398;
w27401 <= not w27399 and not w27400;
w27402 <= w27132 and w27401;
w27403 <= not w27132 and not w27401;
w27404 <= not w27402 and not w27403;
w27405 <= not w27396 and not w27399;
w27406 <= w6 and w26825;
w27407 <= w9802 and w26001;
w27408 <= w10369 and w25995;
w27409 <= not w27407 and not w27408;
w27410 <= not w27406 and w27409;
w27411 <= w9805 and not w26839;
w27412 <= w27410 and not w27411;
w27413 <= a(5) and not w27412;
w27414 <= not w27412 and not w27413;
w27415 <= a(5) and not w27413;
w27416 <= not w27414 and not w27415;
w27417 <= not w27327 and not w27331;
w27418 <= w7918 and w22247;
w27419 <= w7226 and w22258;
w27420 <= w7567 and w22255;
w27421 <= not w27419 and not w27420;
w27422 <= not w27418 and w27421;
w27423 <= w7229 and not w25250;
w27424 <= w27422 and not w27423;
w27425 <= a(11) and not w27424;
w27426 <= not w27424 and not w27425;
w27427 <= a(11) and not w27425;
w27428 <= not w27426 and not w27427;
w27429 <= not w27300 and not w27304;
w27430 <= w6168 and w22270;
w27431 <= w5598 and w22276;
w27432 <= w5874 and w22273;
w27433 <= not w27431 and not w27432;
w27434 <= not w27430 and w27433;
w27435 <= w5601 and not w24102;
w27436 <= w27434 and not w27435;
w27437 <= a(17) and not w27436;
w27438 <= not w27436 and not w27437;
w27439 <= a(17) and not w27437;
w27440 <= not w27438 and not w27439;
w27441 <= not w27273 and not w27277;
w27442 <= w4629 and w22288;
w27443 <= w4468 and w22294;
w27444 <= w4539 and w22291;
w27445 <= not w27443 and not w27444;
w27446 <= not w27442 and w27445;
w27447 <= w4471 and not w22491;
w27448 <= w27446 and not w27447;
w27449 <= a(23) and not w27448;
w27450 <= not w27448 and not w27449;
w27451 <= a(23) and not w27449;
w27452 <= not w27450 and not w27451;
w27453 <= not w27246 and not w27250;
w27454 <= not w27229 and not w27232;
w27455 <= not w27210 and not w27214;
w27456 <= w91 and w2401;
w27457 <= w2928 and w27456;
w27458 <= w1656 and w1672;
w27459 <= w27457 and w27458;
w27460 <= w2345 and w27459;
w27461 <= w4704 and w27460;
w27462 <= w15678 and w27461;
w27463 <= w6667 and w27462;
w27464 <= w6704 and w27463;
w27465 <= w2164 and w27464;
w27466 <= w445 and w27465;
w27467 <= w1761 and w27466;
w27468 <= w1117 and w27467;
w27469 <= not w126 and w27468;
w27470 <= not w275 and w27469;
w27471 <= w2955 and w22315;
w27472 <= w2963 and w22319;
w27473 <= w2958 and w22322;
w27474 <= w10 and w22785;
w27475 <= not w27473 and not w27474;
w27476 <= not w27472 and w27475;
w27477 <= not w27471 and w27476;
w27478 <= not w27470 and not w27477;
w27479 <= not w27470 and not w27478;
w27480 <= not w27477 and not w27478;
w27481 <= not w27479 and not w27480;
w27482 <= not w27455 and not w27481;
w27483 <= not w27455 and not w27482;
w27484 <= not w27481 and not w27482;
w27485 <= not w27483 and not w27484;
w27486 <= w3392 and w22306;
w27487 <= w3477 and w22312;
w27488 <= w3541 and w22309;
w27489 <= not w27487 and not w27488;
w27490 <= not w27486 and w27489;
w27491 <= not w3303 and w27490;
w27492 <= not w22960 and w27490;
w27493 <= not w27491 and not w27492;
w27494 <= a(29) and not w27493;
w27495 <= not a(29) and w27493;
w27496 <= not w27494 and not w27495;
w27497 <= not w27485 and not w27496;
w27498 <= w27485 and w27496;
w27499 <= not w27497 and not w27498;
w27500 <= not w27454 and w27499;
w27501 <= w27454 and not w27499;
w27502 <= not w27500 and not w27501;
w27503 <= w3819 and w22297;
w27504 <= w3902 and w22303;
w27505 <= w3981 and w22300;
w27506 <= not w27504 and not w27505;
w27507 <= not w27503 and w27506;
w27508 <= not w3985 and w27507;
w27509 <= w23255 and w27507;
w27510 <= not w27508 and not w27509;
w27511 <= a(26) and not w27510;
w27512 <= not a(26) and w27510;
w27513 <= not w27511 and not w27512;
w27514 <= w27502 and not w27513;
w27515 <= w27502 and not w27514;
w27516 <= not w27513 and not w27514;
w27517 <= not w27515 and not w27516;
w27518 <= not w27453 and not w27517;
w27519 <= not w27453 and not w27518;
w27520 <= not w27517 and not w27518;
w27521 <= not w27519 and not w27520;
w27522 <= not w27452 and not w27521;
w27523 <= not w27452 and not w27522;
w27524 <= not w27521 and not w27522;
w27525 <= not w27523 and not w27524;
w27526 <= not w27254 and not w27260;
w27527 <= w27525 and w27526;
w27528 <= not w27525 and not w27526;
w27529 <= not w27527 and not w27528;
w27530 <= w5431 and w22279;
w27531 <= w4870 and w22285;
w27532 <= w5342 and w22282;
w27533 <= not w27531 and not w27532;
w27534 <= not w27530 and w27533;
w27535 <= not w4873 and w27534;
w27536 <= w23577 and w27534;
w27537 <= not w27535 and not w27536;
w27538 <= a(20) and not w27537;
w27539 <= not a(20) and w27537;
w27540 <= not w27538 and not w27539;
w27541 <= w27529 and not w27540;
w27542 <= w27529 and not w27541;
w27543 <= not w27540 and not w27541;
w27544 <= not w27542 and not w27543;
w27545 <= not w27441 and not w27544;
w27546 <= not w27441 and not w27545;
w27547 <= not w27544 and not w27545;
w27548 <= not w27546 and not w27547;
w27549 <= not w27440 and not w27548;
w27550 <= not w27440 and not w27549;
w27551 <= not w27548 and not w27549;
w27552 <= not w27550 and not w27551;
w27553 <= not w27281 and not w27287;
w27554 <= w27552 and w27553;
w27555 <= not w27552 and not w27553;
w27556 <= not w27554 and not w27555;
w27557 <= w7036 and w22261;
w27558 <= w6337 and w22267;
w27559 <= w6886 and w22264;
w27560 <= not w27558 and not w27559;
w27561 <= not w27557 and w27560;
w27562 <= not w6332 and w27561;
w27563 <= w24551 and w27561;
w27564 <= not w27562 and not w27563;
w27565 <= a(14) and not w27564;
w27566 <= not a(14) and w27564;
w27567 <= not w27565 and not w27566;
w27568 <= w27556 and not w27567;
w27569 <= w27556 and not w27568;
w27570 <= not w27567 and not w27568;
w27571 <= not w27569 and not w27570;
w27572 <= not w27429 and not w27571;
w27573 <= not w27429 and not w27572;
w27574 <= not w27571 and not w27572;
w27575 <= not w27573 and not w27574;
w27576 <= not w27428 and not w27575;
w27577 <= not w27428 and not w27576;
w27578 <= not w27575 and not w27576;
w27579 <= not w27577 and not w27578;
w27580 <= not w27308 and not w27314;
w27581 <= w27579 and w27580;
w27582 <= not w27579 and not w27580;
w27583 <= not w27581 and not w27582;
w27584 <= w9266 and w25998;
w27585 <= w8353 and w22250;
w27586 <= w8795 and w22244;
w27587 <= not w27585 and not w27586;
w27588 <= not w27584 and w27587;
w27589 <= not w8356 and w27588;
w27590 <= w26539 and w27588;
w27591 <= not w27589 and not w27590;
w27592 <= a(8) and not w27591;
w27593 <= not a(8) and w27591;
w27594 <= not w27592 and not w27593;
w27595 <= w27583 and not w27594;
w27596 <= w27583 and not w27595;
w27597 <= not w27594 and not w27595;
w27598 <= not w27596 and not w27597;
w27599 <= not w27417 and not w27598;
w27600 <= not w27417 and not w27599;
w27601 <= not w27598 and not w27599;
w27602 <= not w27600 and not w27601;
w27603 <= not w27416 and not w27602;
w27604 <= not w27416 and not w27603;
w27605 <= not w27602 and not w27603;
w27606 <= not w27604 and not w27605;
w27607 <= not w27335 and not w27341;
w27608 <= w27606 and w27607;
w27609 <= not w27606 and not w27607;
w27610 <= not w27608 and not w27609;
w27611 <= w10 and w13963;
w27612 <= w2955 and not w13373;
w27613 <= w2958 and not w13562;
w27614 <= w2963 and w13876;
w27615 <= not w27613 and not w27614;
w27616 <= not w27612 and w27615;
w27617 <= not w27611 and w27616;
w27618 <= not w27360 and not w27362;
w27619 <= w3774 and not w27618;
w27620 <= not w3774 and w27618;
w27621 <= not w27619 and not w27620;
w27622 <= not w27617 and w27621;
w27623 <= not w27617 and not w27622;
w27624 <= w27621 and not w27622;
w27625 <= not w27623 and not w27624;
w27626 <= not w27365 and not w27369;
w27627 <= w27625 and w27626;
w27628 <= not w27625 and not w27626;
w27629 <= not w27627 and not w27628;
w27630 <= not w27372 and not w27375;
w27631 <= not w27629 and w27630;
w27632 <= w27629 and not w27630;
w27633 <= not w27631 and not w27632;
w27634 <= w11662 and w27633;
w27635 <= w10990 and w27108;
w27636 <= w11650 and w27377;
w27637 <= not w27635 and not w27636;
w27638 <= not w27634 and w27637;
w27639 <= not w10992 and w27638;
w27640 <= not w27386 and not w27388;
w27641 <= w27377 and w27633;
w27642 <= not w27377 and not w27633;
w27643 <= not w27640 and not w27642;
w27644 <= not w27641 and w27643;
w27645 <= not w27640 and not w27644;
w27646 <= not w27641 and not w27644;
w27647 <= not w27642 and w27646;
w27648 <= not w27645 and not w27647;
w27649 <= w27638 and w27648;
w27650 <= not w27639 and not w27649;
w27651 <= a(2) and not w27650;
w27652 <= not a(2) and w27650;
w27653 <= not w27651 and not w27652;
w27654 <= w27610 and not w27653;
w27655 <= not w27610 and w27653;
w27656 <= not w27654 and not w27655;
w27657 <= not w27405 and w27656;
w27658 <= w27405 and not w27656;
w27659 <= not w27657 and not w27658;
w27660 <= w27402 and w27659;
w27661 <= not w27402 and not w27659;
w27662 <= not w27660 and not w27661;
w27663 <= not w27654 and not w27657;
w27664 <= w6 and w27108;
w27665 <= w9802 and w25995;
w27666 <= w10369 and w26825;
w27667 <= not w27665 and not w27666;
w27668 <= not w27664 and w27667;
w27669 <= w9805 and w27120;
w27670 <= w27668 and not w27669;
w27671 <= a(5) and not w27670;
w27672 <= not w27670 and not w27671;
w27673 <= a(5) and not w27671;
w27674 <= not w27672 and not w27673;
w27675 <= not w27595 and not w27599;
w27676 <= w7918 and w22250;
w27677 <= w7226 and w22255;
w27678 <= w7567 and w22247;
w27679 <= not w27677 and not w27678;
w27680 <= not w27676 and w27679;
w27681 <= w7229 and w25229;
w27682 <= w27680 and not w27681;
w27683 <= a(11) and not w27682;
w27684 <= not w27682 and not w27683;
w27685 <= a(11) and not w27683;
w27686 <= not w27684 and not w27685;
w27687 <= not w27568 and not w27572;
w27688 <= w6168 and w22267;
w27689 <= w5598 and w22273;
w27690 <= w5874 and w22270;
w27691 <= not w27689 and not w27690;
w27692 <= not w27688 and w27691;
w27693 <= w5601 and w22477;
w27694 <= w27692 and not w27693;
w27695 <= a(17) and not w27694;
w27696 <= not w27694 and not w27695;
w27697 <= a(17) and not w27695;
w27698 <= not w27696 and not w27697;
w27699 <= not w27541 and not w27545;
w27700 <= w4629 and w22285;
w27701 <= w4468 and w22291;
w27702 <= w4539 and w22288;
w27703 <= not w27701 and not w27702;
w27704 <= not w27700 and w27703;
w27705 <= w4471 and w23607;
w27706 <= w27704 and not w27705;
w27707 <= a(23) and not w27706;
w27708 <= not w27706 and not w27707;
w27709 <= a(23) and not w27707;
w27710 <= not w27708 and not w27709;
w27711 <= not w27514 and not w27518;
w27712 <= not w27497 and not w27500;
w27713 <= not w27478 and not w27482;
w27714 <= w1358 and w2028;
w27715 <= w3479 and w27714;
w27716 <= w1510 and w27715;
w27717 <= not w46 and w27716;
w27718 <= not w335 and w27717;
w27719 <= not w161 and w27718;
w27720 <= not w141 and w27719;
w27721 <= not w425 and w27720;
w27722 <= not w100 and w27721;
w27723 <= not w726 and w27722;
w27724 <= not w821 and w27723;
w27725 <= w1075 and w2027;
w27726 <= w1616 and w27725;
w27727 <= w1175 and w27726;
w27728 <= w461 and w27727;
w27729 <= w2975 and w27728;
w27730 <= w1644 and w27729;
w27731 <= w3062 and w27730;
w27732 <= w4323 and w27731;
w27733 <= w1947 and w27732;
w27734 <= w27724 and w27733;
w27735 <= w55 and w27734;
w27736 <= w913 and w27735;
w27737 <= w505 and w27736;
w27738 <= not w265 and w27737;
w27739 <= not w537 and w27738;
w27740 <= not w42 and w27739;
w27741 <= not w180 and w27740;
w27742 <= not w364 and w27741;
w27743 <= w2955 and w22312;
w27744 <= w2963 and w22315;
w27745 <= w2958 and w22319;
w27746 <= w10 and not w22769;
w27747 <= not w27745 and not w27746;
w27748 <= not w27744 and w27747;
w27749 <= not w27743 and w27748;
w27750 <= not w27742 and not w27749;
w27751 <= not w27742 and not w27750;
w27752 <= not w27749 and not w27750;
w27753 <= not w27751 and not w27752;
w27754 <= not w27713 and not w27753;
w27755 <= not w27713 and not w27754;
w27756 <= not w27753 and not w27754;
w27757 <= not w27755 and not w27756;
w27758 <= w3392 and w22303;
w27759 <= w3477 and w22309;
w27760 <= w3541 and w22306;
w27761 <= not w27759 and not w27760;
w27762 <= not w27758 and w27761;
w27763 <= not w3303 and w27762;
w27764 <= not w22941 and w27762;
w27765 <= not w27763 and not w27764;
w27766 <= a(29) and not w27765;
w27767 <= not a(29) and w27765;
w27768 <= not w27766 and not w27767;
w27769 <= not w27757 and not w27768;
w27770 <= w27757 and w27768;
w27771 <= not w27769 and not w27770;
w27772 <= not w27712 and w27771;
w27773 <= w27712 and not w27771;
w27774 <= not w27772 and not w27773;
w27775 <= w3819 and w22294;
w27776 <= w3902 and w22300;
w27777 <= w3981 and w22297;
w27778 <= not w27776 and not w27777;
w27779 <= not w27775 and w27778;
w27780 <= not w3985 and w27779;
w27781 <= not w23303 and w27779;
w27782 <= not w27780 and not w27781;
w27783 <= a(26) and not w27782;
w27784 <= not a(26) and w27782;
w27785 <= not w27783 and not w27784;
w27786 <= w27774 and not w27785;
w27787 <= w27774 and not w27786;
w27788 <= not w27785 and not w27786;
w27789 <= not w27787 and not w27788;
w27790 <= not w27711 and not w27789;
w27791 <= not w27711 and not w27790;
w27792 <= not w27789 and not w27790;
w27793 <= not w27791 and not w27792;
w27794 <= not w27710 and not w27793;
w27795 <= not w27710 and not w27794;
w27796 <= not w27793 and not w27794;
w27797 <= not w27795 and not w27796;
w27798 <= not w27522 and not w27528;
w27799 <= w27797 and w27798;
w27800 <= not w27797 and not w27798;
w27801 <= not w27799 and not w27800;
w27802 <= w5431 and w22276;
w27803 <= w4870 and w22282;
w27804 <= w5342 and w22279;
w27805 <= not w27803 and not w27804;
w27806 <= not w27802 and w27805;
w27807 <= not w4873 and w27806;
w27808 <= not w24077 and w27806;
w27809 <= not w27807 and not w27808;
w27810 <= a(20) and not w27809;
w27811 <= not a(20) and w27809;
w27812 <= not w27810 and not w27811;
w27813 <= w27801 and not w27812;
w27814 <= w27801 and not w27813;
w27815 <= not w27812 and not w27813;
w27816 <= not w27814 and not w27815;
w27817 <= not w27699 and not w27816;
w27818 <= not w27699 and not w27817;
w27819 <= not w27816 and not w27817;
w27820 <= not w27818 and not w27819;
w27821 <= not w27698 and not w27820;
w27822 <= not w27698 and not w27821;
w27823 <= not w27820 and not w27821;
w27824 <= not w27822 and not w27823;
w27825 <= not w27549 and not w27555;
w27826 <= w27824 and w27825;
w27827 <= not w27824 and not w27825;
w27828 <= not w27826 and not w27827;
w27829 <= w7036 and w22258;
w27830 <= w6337 and w22264;
w27831 <= w6886 and w22261;
w27832 <= not w27830 and not w27831;
w27833 <= not w27829 and w27832;
w27834 <= not w6332 and w27833;
w27835 <= not w24534 and w27833;
w27836 <= not w27834 and not w27835;
w27837 <= a(14) and not w27836;
w27838 <= not a(14) and w27836;
w27839 <= not w27837 and not w27838;
w27840 <= w27828 and not w27839;
w27841 <= w27828 and not w27840;
w27842 <= not w27839 and not w27840;
w27843 <= not w27841 and not w27842;
w27844 <= not w27687 and not w27843;
w27845 <= not w27687 and not w27844;
w27846 <= not w27843 and not w27844;
w27847 <= not w27845 and not w27846;
w27848 <= not w27686 and not w27847;
w27849 <= not w27686 and not w27848;
w27850 <= not w27847 and not w27848;
w27851 <= not w27849 and not w27850;
w27852 <= not w27576 and not w27582;
w27853 <= w27851 and w27852;
w27854 <= not w27851 and not w27852;
w27855 <= not w27853 and not w27854;
w27856 <= w9266 and w26001;
w27857 <= w8353 and w22244;
w27858 <= w8795 and w25998;
w27859 <= not w27857 and not w27858;
w27860 <= not w27856 and w27859;
w27861 <= not w8356 and w27860;
w27862 <= w26559 and w27860;
w27863 <= not w27861 and not w27862;
w27864 <= a(8) and not w27863;
w27865 <= not a(8) and w27863;
w27866 <= not w27864 and not w27865;
w27867 <= w27855 and not w27866;
w27868 <= w27855 and not w27867;
w27869 <= not w27866 and not w27867;
w27870 <= not w27868 and not w27869;
w27871 <= not w27675 and not w27870;
w27872 <= not w27675 and not w27871;
w27873 <= not w27870 and not w27871;
w27874 <= not w27872 and not w27873;
w27875 <= not w27674 and not w27874;
w27876 <= not w27674 and not w27875;
w27877 <= not w27874 and not w27875;
w27878 <= not w27876 and not w27877;
w27879 <= not w27603 and not w27609;
w27880 <= w27878 and w27879;
w27881 <= not w27878 and not w27879;
w27882 <= not w27880 and not w27881;
w27883 <= w10 and not w13886;
w27884 <= not w2955 and not w2963;
w27885 <= not w13373 and not w27884;
w27886 <= w2958 and w13876;
w27887 <= not w27885 and not w27886;
w27888 <= not w27883 and w27887;
w27889 <= w3774 and w27888;
w27890 <= not w3774 and not w27888;
w27891 <= not w27889 and not w27890;
w27892 <= not w27619 and not w27622;
w27893 <= w27891 and w27892;
w27894 <= not w27891 and not w27892;
w27895 <= not w27893 and not w27894;
w27896 <= not w27628 and not w27632;
w27897 <= not w27895 and w27896;
w27898 <= w27895 and not w27896;
w27899 <= not w27897 and not w27898;
w27900 <= w11662 and w27899;
w27901 <= w10990 and w27377;
w27902 <= w11650 and w27633;
w27903 <= not w27901 and not w27902;
w27904 <= not w27900 and w27903;
w27905 <= not w10992 and w27904;
w27906 <= not w27633 and not w27899;
w27907 <= w27633 and w27899;
w27908 <= not w27906 and not w27907;
w27909 <= not w27646 and w27908;
w27910 <= w27646 and not w27908;
w27911 <= not w27909 and not w27910;
w27912 <= w27904 and not w27911;
w27913 <= not w27905 and not w27912;
w27914 <= a(2) and not w27913;
w27915 <= not a(2) and w27913;
w27916 <= not w27914 and not w27915;
w27917 <= w27882 and not w27916;
w27918 <= not w27882 and w27916;
w27919 <= not w27917 and not w27918;
w27920 <= not w27663 and w27919;
w27921 <= w27663 and not w27919;
w27922 <= not w27920 and not w27921;
w27923 <= w27660 and w27922;
w27924 <= not w27660 and not w27922;
w27925 <= not w27923 and not w27924;
w27926 <= not w27917 and not w27920;
w27927 <= w6 and w27377;
w27928 <= w9802 and w26825;
w27929 <= w10369 and w27108;
w27930 <= not w27928 and not w27929;
w27931 <= not w27927 and w27930;
w27932 <= w9805 and w27390;
w27933 <= w27931 and not w27932;
w27934 <= a(5) and not w27933;
w27935 <= not w27933 and not w27934;
w27936 <= a(5) and not w27934;
w27937 <= not w27935 and not w27936;
w27938 <= not w27867 and not w27871;
w27939 <= w7918 and w22244;
w27940 <= w7226 and w22247;
w27941 <= w7567 and w22250;
w27942 <= not w27940 and not w27941;
w27943 <= not w27939 and w27942;
w27944 <= w7229 and not w22464;
w27945 <= w27943 and not w27944;
w27946 <= a(11) and not w27945;
w27947 <= not w27945 and not w27946;
w27948 <= a(11) and not w27946;
w27949 <= not w27947 and not w27948;
w27950 <= not w27840 and not w27844;
w27951 <= w6168 and w22264;
w27952 <= w5598 and w22270;
w27953 <= w5874 and w22267;
w27954 <= not w27952 and not w27953;
w27955 <= not w27951 and w27954;
w27956 <= w5601 and not w24568;
w27957 <= w27955 and not w27956;
w27958 <= a(17) and not w27957;
w27959 <= not w27957 and not w27958;
w27960 <= a(17) and not w27958;
w27961 <= not w27959 and not w27960;
w27962 <= not w27813 and not w27817;
w27963 <= w4629 and w22282;
w27964 <= w4468 and w22288;
w27965 <= w4539 and w22285;
w27966 <= not w27964 and not w27965;
w27967 <= not w27963 and w27966;
w27968 <= w4471 and not w23594;
w27969 <= w27967 and not w27968;
w27970 <= a(23) and not w27969;
w27971 <= not w27969 and not w27970;
w27972 <= a(23) and not w27970;
w27973 <= not w27971 and not w27972;
w27974 <= not w27786 and not w27790;
w27975 <= not w27769 and not w27772;
w27976 <= not w27750 and not w27754;
w27977 <= w142 and w3522;
w27978 <= w625 and w27977;
w27979 <= w12344 and w27978;
w27980 <= w15905 and w27979;
w27981 <= w3579 and w27980;
w27982 <= w5221 and w27981;
w27983 <= w981 and w27982;
w27984 <= not w404 and w27983;
w27985 <= not w46 and w27984;
w27986 <= not w177 and w27985;
w27987 <= not w106 and w27986;
w27988 <= not w536 and w27987;
w27989 <= not w310 and w27988;
w27990 <= not w428 and w27989;
w27991 <= not w96 and w27990;
w27992 <= not w186 and w27991;
w27993 <= not w93 and w27992;
w27994 <= not w157 and w27993;
w27995 <= w2955 and w22309;
w27996 <= w2963 and w22312;
w27997 <= w2958 and w22315;
w27998 <= w10 and w22504;
w27999 <= not w27997 and not w27998;
w28000 <= not w27996 and w27999;
w28001 <= not w27995 and w28000;
w28002 <= not w27994 and not w28001;
w28003 <= not w27994 and not w28002;
w28004 <= not w28001 and not w28002;
w28005 <= not w28003 and not w28004;
w28006 <= not w27976 and not w28005;
w28007 <= not w27976 and not w28006;
w28008 <= not w28005 and not w28006;
w28009 <= not w28007 and not w28008;
w28010 <= w3392 and w22300;
w28011 <= w3477 and w22306;
w28012 <= w3541 and w22303;
w28013 <= not w28011 and not w28012;
w28014 <= not w28010 and w28013;
w28015 <= not w3303 and w28014;
w28016 <= w22928 and w28014;
w28017 <= not w28015 and not w28016;
w28018 <= a(29) and not w28017;
w28019 <= not a(29) and w28017;
w28020 <= not w28018 and not w28019;
w28021 <= not w28009 and not w28020;
w28022 <= w28009 and w28020;
w28023 <= not w28021 and not w28022;
w28024 <= not w27975 and w28023;
w28025 <= w27975 and not w28023;
w28026 <= not w28024 and not w28025;
w28027 <= w3819 and w22291;
w28028 <= w3902 and w22297;
w28029 <= w3981 and w22294;
w28030 <= not w28028 and not w28029;
w28031 <= not w28027 and w28030;
w28032 <= not w3985 and w28031;
w28033 <= w23280 and w28031;
w28034 <= not w28032 and not w28033;
w28035 <= a(26) and not w28034;
w28036 <= not a(26) and w28034;
w28037 <= not w28035 and not w28036;
w28038 <= w28026 and not w28037;
w28039 <= w28026 and not w28038;
w28040 <= not w28037 and not w28038;
w28041 <= not w28039 and not w28040;
w28042 <= not w27974 and not w28041;
w28043 <= not w27974 and not w28042;
w28044 <= not w28041 and not w28042;
w28045 <= not w28043 and not w28044;
w28046 <= not w27973 and not w28045;
w28047 <= not w27973 and not w28046;
w28048 <= not w28045 and not w28046;
w28049 <= not w28047 and not w28048;
w28050 <= not w27794 and not w27800;
w28051 <= w28049 and w28050;
w28052 <= not w28049 and not w28050;
w28053 <= not w28051 and not w28052;
w28054 <= w5431 and w22273;
w28055 <= w4870 and w22279;
w28056 <= w5342 and w22276;
w28057 <= not w28055 and not w28056;
w28058 <= not w28054 and w28057;
w28059 <= not w4873 and w28058;
w28060 <= w24123 and w28058;
w28061 <= not w28059 and not w28060;
w28062 <= a(20) and not w28061;
w28063 <= not a(20) and w28061;
w28064 <= not w28062 and not w28063;
w28065 <= w28053 and not w28064;
w28066 <= w28053 and not w28065;
w28067 <= not w28064 and not w28065;
w28068 <= not w28066 and not w28067;
w28069 <= not w27962 and not w28068;
w28070 <= not w27962 and not w28069;
w28071 <= not w28068 and not w28069;
w28072 <= not w28070 and not w28071;
w28073 <= not w27961 and not w28072;
w28074 <= not w27961 and not w28073;
w28075 <= not w28072 and not w28073;
w28076 <= not w28074 and not w28075;
w28077 <= not w27821 and not w27827;
w28078 <= w28076 and w28077;
w28079 <= not w28076 and not w28077;
w28080 <= not w28078 and not w28079;
w28081 <= w7036 and w22255;
w28082 <= w6337 and w22261;
w28083 <= w6886 and w22258;
w28084 <= not w28082 and not w28083;
w28085 <= not w28081 and w28084;
w28086 <= not w6332 and w28085;
w28087 <= w25205 and w28085;
w28088 <= not w28086 and not w28087;
w28089 <= a(14) and not w28088;
w28090 <= not a(14) and w28088;
w28091 <= not w28089 and not w28090;
w28092 <= w28080 and not w28091;
w28093 <= w28080 and not w28092;
w28094 <= not w28091 and not w28092;
w28095 <= not w28093 and not w28094;
w28096 <= not w27950 and not w28095;
w28097 <= not w27950 and not w28096;
w28098 <= not w28095 and not w28096;
w28099 <= not w28097 and not w28098;
w28100 <= not w27949 and not w28099;
w28101 <= not w27949 and not w28100;
w28102 <= not w28099 and not w28100;
w28103 <= not w28101 and not w28102;
w28104 <= not w27848 and not w27854;
w28105 <= w28103 and w28104;
w28106 <= not w28103 and not w28104;
w28107 <= not w28105 and not w28106;
w28108 <= w9266 and w25995;
w28109 <= w8353 and w25998;
w28110 <= w8795 and w26001;
w28111 <= not w28109 and not w28110;
w28112 <= not w28108 and w28111;
w28113 <= not w8356 and w28112;
w28114 <= w26023 and w28112;
w28115 <= not w28113 and not w28114;
w28116 <= a(8) and not w28115;
w28117 <= not a(8) and w28115;
w28118 <= not w28116 and not w28117;
w28119 <= w28107 and not w28118;
w28120 <= w28107 and not w28119;
w28121 <= not w28118 and not w28119;
w28122 <= not w28120 and not w28121;
w28123 <= not w27938 and not w28122;
w28124 <= not w27938 and not w28123;
w28125 <= not w28122 and not w28123;
w28126 <= not w28124 and not w28125;
w28127 <= not w27937 and not w28126;
w28128 <= not w27937 and not w28127;
w28129 <= not w28126 and not w28127;
w28130 <= not w28128 and not w28129;
w28131 <= not w27875 and not w27881;
w28132 <= w28130 and w28131;
w28133 <= not w28130 and not w28131;
w28134 <= not w28132 and not w28133;
w28135 <= not w27894 and not w27898;
w28136 <= not a(31) and w32;
w28137 <= not w13373 and not w28136;
w28138 <= w27889 and not w28137;
w28139 <= not w27889 and w28137;
w28140 <= not w28138 and not w28139;
w28141 <= w28135 and not w28140;
w28142 <= not w28135 and w28140;
w28143 <= not w28141 and not w28142;
w28144 <= w11662 and not w28143;
w28145 <= w10990 and w27633;
w28146 <= w11650 and w27899;
w28147 <= not w28145 and not w28146;
w28148 <= not w28144 and w28147;
w28149 <= not w10992 and w28148;
w28150 <= not w27907 and not w27909;
w28151 <= w27899 and not w28143;
w28152 <= not w27899 and w28143;
w28153 <= not w28150 and not w28152;
w28154 <= not w28151 and w28153;
w28155 <= not w28150 and not w28154;
w28156 <= not w28151 and not w28154;
w28157 <= not w28152 and w28156;
w28158 <= not w28155 and not w28157;
w28159 <= w28148 and w28158;
w28160 <= not w28149 and not w28159;
w28161 <= a(2) and not w28160;
w28162 <= not a(2) and w28160;
w28163 <= not w28161 and not w28162;
w28164 <= w28134 and not w28163;
w28165 <= not w28134 and w28163;
w28166 <= not w28164 and not w28165;
w28167 <= not w27926 and w28166;
w28168 <= w27926 and not w28166;
w28169 <= not w28167 and not w28168;
w28170 <= w27923 and w28169;
w28171 <= not w27923 and not w28169;
w28172 <= not w28170 and not w28171;
w28173 <= w6 and w27633;
w28174 <= w9802 and w27108;
w28175 <= w10369 and w27377;
w28176 <= not w28174 and not w28175;
w28177 <= not w28173 and w28176;
w28178 <= w9805 and not w27648;
w28179 <= w28177 and not w28178;
w28180 <= a(5) and not w28179;
w28181 <= not w28179 and not w28180;
w28182 <= a(5) and not w28180;
w28183 <= not w28181 and not w28182;
w28184 <= not w28119 and not w28123;
w28185 <= w7918 and w25998;
w28186 <= w7226 and w22250;
w28187 <= w7567 and w22244;
w28188 <= not w28186 and not w28187;
w28189 <= not w28185 and w28188;
w28190 <= w7229 and not w26539;
w28191 <= w28189 and not w28190;
w28192 <= a(11) and not w28191;
w28193 <= not w28191 and not w28192;
w28194 <= a(11) and not w28192;
w28195 <= not w28193 and not w28194;
w28196 <= not w28092 and not w28096;
w28197 <= w6168 and w22261;
w28198 <= w5598 and w22267;
w28199 <= w5874 and w22264;
w28200 <= not w28198 and not w28199;
w28201 <= not w28197 and w28200;
w28202 <= w5601 and not w24551;
w28203 <= w28201 and not w28202;
w28204 <= a(17) and not w28203;
w28205 <= not w28203 and not w28204;
w28206 <= a(17) and not w28204;
w28207 <= not w28205 and not w28206;
w28208 <= not w28065 and not w28069;
w28209 <= w4629 and w22279;
w28210 <= w4468 and w22285;
w28211 <= w4539 and w22282;
w28212 <= not w28210 and not w28211;
w28213 <= not w28209 and w28212;
w28214 <= w4471 and not w23577;
w28215 <= w28213 and not w28214;
w28216 <= a(23) and not w28215;
w28217 <= not w28215 and not w28216;
w28218 <= a(23) and not w28216;
w28219 <= not w28217 and not w28218;
w28220 <= not w28038 and not w28042;
w28221 <= not w28021 and not w28024;
w28222 <= not w28002 and not w28006;
w28223 <= w1485 and w1628;
w28224 <= not w104 and w28223;
w28225 <= not w163 and w28224;
w28226 <= not w126 and w28225;
w28227 <= not w502 and w28226;
w28228 <= not w260 and w28227;
w28229 <= not w93 and w28228;
w28230 <= w232 and w27457;
w28231 <= w372 and w28230;
w28232 <= w2975 and w28231;
w28233 <= w28229 and w28232;
w28234 <= w14500 and w28233;
w28235 <= w4948 and w28234;
w28236 <= w14982 and w28235;
w28237 <= w442 and w28236;
w28238 <= w913 and w28237;
w28239 <= w162 and w28238;
w28240 <= w2340 and w28239;
w28241 <= w51 and w28240;
w28242 <= not w591 and w28241;
w28243 <= not w181 and w28242;
w28244 <= not w307 and w28243;
w28245 <= not w592 and w28244;
w28246 <= not w647 and w28245;
w28247 <= not w30 and w28246;
w28248 <= not w821 and w28247;
w28249 <= not w363 and w28248;
w28250 <= w2955 and w22306;
w28251 <= w2963 and w22309;
w28252 <= w2958 and w22312;
w28253 <= w10 and w22960;
w28254 <= not w28252 and not w28253;
w28255 <= not w28251 and w28254;
w28256 <= not w28250 and w28255;
w28257 <= not w28249 and not w28256;
w28258 <= not w28249 and not w28257;
w28259 <= not w28256 and not w28257;
w28260 <= not w28258 and not w28259;
w28261 <= not w28222 and not w28260;
w28262 <= not w28222 and not w28261;
w28263 <= not w28260 and not w28261;
w28264 <= not w28262 and not w28263;
w28265 <= w3392 and w22297;
w28266 <= w3477 and w22303;
w28267 <= w3541 and w22300;
w28268 <= not w28266 and not w28267;
w28269 <= not w28265 and w28268;
w28270 <= not w3303 and w28269;
w28271 <= w23255 and w28269;
w28272 <= not w28270 and not w28271;
w28273 <= a(29) and not w28272;
w28274 <= not a(29) and w28272;
w28275 <= not w28273 and not w28274;
w28276 <= not w28264 and not w28275;
w28277 <= w28264 and w28275;
w28278 <= not w28276 and not w28277;
w28279 <= not w28221 and w28278;
w28280 <= w28221 and not w28278;
w28281 <= not w28279 and not w28280;
w28282 <= w3819 and w22288;
w28283 <= w3902 and w22294;
w28284 <= w3981 and w22291;
w28285 <= not w28283 and not w28284;
w28286 <= not w28282 and w28285;
w28287 <= not w3985 and w28286;
w28288 <= w22491 and w28286;
w28289 <= not w28287 and not w28288;
w28290 <= a(26) and not w28289;
w28291 <= not a(26) and w28289;
w28292 <= not w28290 and not w28291;
w28293 <= w28281 and not w28292;
w28294 <= not w28281 and w28292;
w28295 <= not w28293 and not w28294;
w28296 <= not w28220 and w28295;
w28297 <= w28220 and not w28295;
w28298 <= not w28296 and not w28297;
w28299 <= not w28219 and w28298;
w28300 <= not w28219 and not w28299;
w28301 <= w28298 and not w28299;
w28302 <= not w28300 and not w28301;
w28303 <= not w28046 and not w28052;
w28304 <= w28302 and w28303;
w28305 <= not w28302 and not w28303;
w28306 <= not w28304 and not w28305;
w28307 <= w5431 and w22270;
w28308 <= w4870 and w22276;
w28309 <= w5342 and w22273;
w28310 <= not w28308 and not w28309;
w28311 <= not w28307 and w28310;
w28312 <= not w4873 and w28311;
w28313 <= w24102 and w28311;
w28314 <= not w28312 and not w28313;
w28315 <= a(20) and not w28314;
w28316 <= not a(20) and w28314;
w28317 <= not w28315 and not w28316;
w28318 <= w28306 and not w28317;
w28319 <= not w28306 and w28317;
w28320 <= not w28318 and not w28319;
w28321 <= not w28208 and w28320;
w28322 <= w28208 and not w28320;
w28323 <= not w28321 and not w28322;
w28324 <= not w28207 and w28323;
w28325 <= not w28207 and not w28324;
w28326 <= w28323 and not w28324;
w28327 <= not w28325 and not w28326;
w28328 <= not w28073 and not w28079;
w28329 <= w28327 and w28328;
w28330 <= not w28327 and not w28328;
w28331 <= not w28329 and not w28330;
w28332 <= w7036 and w22247;
w28333 <= w6337 and w22258;
w28334 <= w6886 and w22255;
w28335 <= not w28333 and not w28334;
w28336 <= not w28332 and w28335;
w28337 <= not w6332 and w28336;
w28338 <= w25250 and w28336;
w28339 <= not w28337 and not w28338;
w28340 <= a(14) and not w28339;
w28341 <= not a(14) and w28339;
w28342 <= not w28340 and not w28341;
w28343 <= w28331 and not w28342;
w28344 <= not w28331 and w28342;
w28345 <= not w28343 and not w28344;
w28346 <= not w28196 and w28345;
w28347 <= w28196 and not w28345;
w28348 <= not w28346 and not w28347;
w28349 <= not w28195 and w28348;
w28350 <= not w28195 and not w28349;
w28351 <= w28348 and not w28349;
w28352 <= not w28350 and not w28351;
w28353 <= not w28100 and not w28106;
w28354 <= w28352 and w28353;
w28355 <= not w28352 and not w28353;
w28356 <= not w28354 and not w28355;
w28357 <= w9266 and w26825;
w28358 <= w8353 and w26001;
w28359 <= w8795 and w25995;
w28360 <= not w28358 and not w28359;
w28361 <= not w28357 and w28360;
w28362 <= not w8356 and w28361;
w28363 <= w26839 and w28361;
w28364 <= not w28362 and not w28363;
w28365 <= a(8) and not w28364;
w28366 <= not a(8) and w28364;
w28367 <= not w28365 and not w28366;
w28368 <= w28356 and not w28367;
w28369 <= not w28356 and w28367;
w28370 <= not w28368 and not w28369;
w28371 <= not w28184 and w28370;
w28372 <= w28184 and not w28370;
w28373 <= not w28371 and not w28372;
w28374 <= not w28183 and w28373;
w28375 <= not w28183 and not w28374;
w28376 <= w28373 and not w28374;
w28377 <= not w28375 and not w28376;
w28378 <= not w20756 and not w28143;
w28379 <= w10990 and w27899;
w28380 <= not w28378 and not w28379;
w28381 <= w10992 and not w28156;
w28382 <= w28380 and not w28381;
w28383 <= a(2) and not w28382;
w28384 <= a(2) and not w28383;
w28385 <= not w28382 and not w28383;
w28386 <= not w28384 and not w28385;
w28387 <= not w28377 and not w28386;
w28388 <= not w28377 and not w28387;
w28389 <= not w28386 and not w28387;
w28390 <= not w28388 and not w28389;
w28391 <= not w28127 and not w28133;
w28392 <= w28390 and w28391;
w28393 <= not w28390 and not w28391;
w28394 <= not w28392 and not w28393;
w28395 <= not w28164 and not w28167;
w28396 <= not w28394 and w28395;
w28397 <= w28394 and not w28395;
w28398 <= not w28396 and not w28397;
w28399 <= w28170 and w28398;
w28400 <= not w28170 and not w28398;
w28401 <= not w28399 and not w28400;
w28402 <= not w28276 and not w28279;
w28403 <= w10 and w22941;
w28404 <= w2955 and w22303;
w28405 <= w2958 and w22309;
w28406 <= w2963 and w22306;
w28407 <= not w28405 and not w28406;
w28408 <= not w28404 and w28407;
w28409 <= not w28403 and w28408;
w28410 <= w2050 and w2358;
w28411 <= w6669 and w28410;
w28412 <= w13633 and w28411;
w28413 <= w1957 and w28412;
w28414 <= w12879 and w28413;
w28415 <= w1512 and w28414;
w28416 <= w3692 and w28415;
w28417 <= w1819 and w28416;
w28418 <= w1509 and w28417;
w28419 <= w3919 and w28418;
w28420 <= w2418 and w28419;
w28421 <= w1324 and w28420;
w28422 <= not w782 and w28421;
w28423 <= not w554 and w28422;
w28424 <= not w536 and w28423;
w28425 <= not w472 and w28424;
w28426 <= not w92 and w28425;
w28427 <= not w466 and w28426;
w28428 <= not w14966 and not w28143;
w28429 <= a(2) and not w28428;
w28430 <= not a(2) and w28428;
w28431 <= not w28429 and not w28430;
w28432 <= not w28427 and not w28431;
w28433 <= w28427 and w28431;
w28434 <= not w28409 and not w28433;
w28435 <= not w28432 and w28434;
w28436 <= not w28409 and not w28435;
w28437 <= not w28432 and not w28435;
w28438 <= not w28433 and w28437;
w28439 <= not w28436 and not w28438;
w28440 <= not w28257 and not w28261;
w28441 <= w28439 and w28440;
w28442 <= not w28439 and not w28440;
w28443 <= not w28441 and not w28442;
w28444 <= w3392 and w22294;
w28445 <= w3477 and w22300;
w28446 <= w3541 and w22297;
w28447 <= not w28445 and not w28446;
w28448 <= not w28444 and w28447;
w28449 <= not w3303 and w28448;
w28450 <= not w23303 and w28448;
w28451 <= not w28449 and not w28450;
w28452 <= a(29) and not w28451;
w28453 <= not a(29) and w28451;
w28454 <= not w28452 and not w28453;
w28455 <= w28443 and not w28454;
w28456 <= not w28443 and w28454;
w28457 <= not w28455 and not w28456;
w28458 <= not w28402 and w28457;
w28459 <= w28402 and not w28457;
w28460 <= not w28458 and not w28459;
w28461 <= w3819 and w22285;
w28462 <= w3902 and w22291;
w28463 <= w3981 and w22288;
w28464 <= not w28462 and not w28463;
w28465 <= not w28461 and w28464;
w28466 <= w3985 and w23607;
w28467 <= w28465 and not w28466;
w28468 <= a(26) and not w28467;
w28469 <= a(26) and not w28468;
w28470 <= not w28467 and not w28468;
w28471 <= not w28469 and not w28470;
w28472 <= w28460 and not w28471;
w28473 <= w28460 and not w28472;
w28474 <= not w28471 and not w28472;
w28475 <= not w28473 and not w28474;
w28476 <= not w28293 and not w28296;
w28477 <= w28475 and w28476;
w28478 <= not w28475 and not w28476;
w28479 <= not w28477 and not w28478;
w28480 <= w4629 and w22276;
w28481 <= w4468 and w22282;
w28482 <= w4539 and w22279;
w28483 <= not w28481 and not w28482;
w28484 <= not w28480 and w28483;
w28485 <= w4471 and w24077;
w28486 <= w28484 and not w28485;
w28487 <= a(23) and not w28486;
w28488 <= a(23) and not w28487;
w28489 <= not w28486 and not w28487;
w28490 <= not w28488 and not w28489;
w28491 <= w28479 and not w28490;
w28492 <= w28479 and not w28491;
w28493 <= not w28490 and not w28491;
w28494 <= not w28492 and not w28493;
w28495 <= not w28299 and not w28305;
w28496 <= w28494 and w28495;
w28497 <= not w28494 and not w28495;
w28498 <= not w28496 and not w28497;
w28499 <= w5431 and w22267;
w28500 <= w4870 and w22273;
w28501 <= w5342 and w22270;
w28502 <= not w28500 and not w28501;
w28503 <= not w28499 and w28502;
w28504 <= w4873 and w22477;
w28505 <= w28503 and not w28504;
w28506 <= a(20) and not w28505;
w28507 <= a(20) and not w28506;
w28508 <= not w28505 and not w28506;
w28509 <= not w28507 and not w28508;
w28510 <= w28498 and not w28509;
w28511 <= w28498 and not w28510;
w28512 <= not w28509 and not w28510;
w28513 <= not w28511 and not w28512;
w28514 <= not w28318 and not w28321;
w28515 <= w28513 and w28514;
w28516 <= not w28513 and not w28514;
w28517 <= not w28515 and not w28516;
w28518 <= w6168 and w22258;
w28519 <= w5598 and w22264;
w28520 <= w5874 and w22261;
w28521 <= not w28519 and not w28520;
w28522 <= not w28518 and w28521;
w28523 <= w5601 and w24534;
w28524 <= w28522 and not w28523;
w28525 <= a(17) and not w28524;
w28526 <= a(17) and not w28525;
w28527 <= not w28524 and not w28525;
w28528 <= not w28526 and not w28527;
w28529 <= w28517 and not w28528;
w28530 <= w28517 and not w28529;
w28531 <= not w28528 and not w28529;
w28532 <= not w28530 and not w28531;
w28533 <= not w28324 and not w28330;
w28534 <= w28532 and w28533;
w28535 <= not w28532 and not w28533;
w28536 <= not w28534 and not w28535;
w28537 <= w7036 and w22250;
w28538 <= w6337 and w22255;
w28539 <= w6886 and w22247;
w28540 <= not w28538 and not w28539;
w28541 <= not w28537 and w28540;
w28542 <= w6332 and w25229;
w28543 <= w28541 and not w28542;
w28544 <= a(14) and not w28543;
w28545 <= a(14) and not w28544;
w28546 <= not w28543 and not w28544;
w28547 <= not w28545 and not w28546;
w28548 <= w28536 and not w28547;
w28549 <= w28536 and not w28548;
w28550 <= not w28547 and not w28548;
w28551 <= not w28549 and not w28550;
w28552 <= not w28343 and not w28346;
w28553 <= w28551 and w28552;
w28554 <= not w28551 and not w28552;
w28555 <= not w28553 and not w28554;
w28556 <= w7918 and w26001;
w28557 <= w7226 and w22244;
w28558 <= w7567 and w25998;
w28559 <= not w28557 and not w28558;
w28560 <= not w28556 and w28559;
w28561 <= w7229 and not w26559;
w28562 <= w28560 and not w28561;
w28563 <= a(11) and not w28562;
w28564 <= a(11) and not w28563;
w28565 <= not w28562 and not w28563;
w28566 <= not w28564 and not w28565;
w28567 <= w28555 and not w28566;
w28568 <= w28555 and not w28567;
w28569 <= not w28566 and not w28567;
w28570 <= not w28568 and not w28569;
w28571 <= not w28349 and not w28355;
w28572 <= w28570 and w28571;
w28573 <= not w28570 and not w28571;
w28574 <= not w28572 and not w28573;
w28575 <= w9266 and w27108;
w28576 <= w8353 and w25995;
w28577 <= w8795 and w26825;
w28578 <= not w28576 and not w28577;
w28579 <= not w28575 and w28578;
w28580 <= w8356 and w27120;
w28581 <= w28579 and not w28580;
w28582 <= a(8) and not w28581;
w28583 <= a(8) and not w28582;
w28584 <= not w28581 and not w28582;
w28585 <= not w28583 and not w28584;
w28586 <= w28574 and not w28585;
w28587 <= w28574 and not w28586;
w28588 <= not w28585 and not w28586;
w28589 <= not w28587 and not w28588;
w28590 <= not w28368 and not w28371;
w28591 <= w28589 and w28590;
w28592 <= not w28589 and not w28590;
w28593 <= not w28591 and not w28592;
w28594 <= w6 and w27899;
w28595 <= w9802 and w27377;
w28596 <= w10369 and w27633;
w28597 <= not w28595 and not w28596;
w28598 <= not w28594 and w28597;
w28599 <= w9805 and w27911;
w28600 <= w28598 and not w28599;
w28601 <= a(5) and not w28600;
w28602 <= a(5) and not w28601;
w28603 <= not w28600 and not w28601;
w28604 <= not w28602 and not w28603;
w28605 <= w28593 and not w28604;
w28606 <= w28593 and not w28605;
w28607 <= not w28604 and not w28605;
w28608 <= not w28606 and not w28607;
w28609 <= not w28374 and not w28387;
w28610 <= w28608 and w28609;
w28611 <= not w28608 and not w28609;
w28612 <= not w28610 and not w28611;
w28613 <= not w28393 and not w28397;
w28614 <= not w28612 and w28613;
w28615 <= w28612 and not w28613;
w28616 <= not w28614 and not w28615;
w28617 <= w28399 and w28616;
w28618 <= not w28399 and not w28616;
w28619 <= not w28617 and not w28618;
w28620 <= w655 and w15955;
w28621 <= not w236 and w28620;
w28622 <= not w506 and w28621;
w28623 <= not w821 and w28622;
w28624 <= w1282 and w23186;
w28625 <= w1359 and w28624;
w28626 <= w2345 and w28625;
w28627 <= w28623 and w28626;
w28628 <= w16002 and w28627;
w28629 <= w1248 and w28628;
w28630 <= w1717 and w28629;
w28631 <= w804 and w28630;
w28632 <= w914 and w28631;
w28633 <= w334 and w28632;
w28634 <= w2518 and w28633;
w28635 <= w2023 and w28634;
w28636 <= w3098 and w28635;
w28637 <= w214 and w28636;
w28638 <= not w56 and w28637;
w28639 <= not w218 and w28638;
w28640 <= not w601 and w28639;
w28641 <= not w298 and w28640;
w28642 <= not w28431 and not w28641;
w28643 <= w28431 and w28641;
w28644 <= not w28437 and not w28643;
w28645 <= not w28642 and w28644;
w28646 <= not w28437 and not w28645;
w28647 <= not w28642 and not w28645;
w28648 <= not w28643 and w28647;
w28649 <= not w28646 and not w28648;
w28650 <= w10 and not w22928;
w28651 <= w2955 and w22300;
w28652 <= w2958 and w22306;
w28653 <= w2963 and w22303;
w28654 <= not w28652 and not w28653;
w28655 <= not w28651 and w28654;
w28656 <= not w28650 and w28655;
w28657 <= not w28649 and not w28656;
w28658 <= not w28649 and not w28657;
w28659 <= not w28656 and not w28657;
w28660 <= not w28658 and not w28659;
w28661 <= not w28442 and not w28455;
w28662 <= w28660 and w28661;
w28663 <= not w28660 and not w28661;
w28664 <= not w28662 and not w28663;
w28665 <= w3392 and w22291;
w28666 <= w3477 and w22297;
w28667 <= w3541 and w22294;
w28668 <= not w28666 and not w28667;
w28669 <= not w28665 and w28668;
w28670 <= w3303 and not w23280;
w28671 <= w28669 and not w28670;
w28672 <= a(29) and not w28671;
w28673 <= a(29) and not w28672;
w28674 <= not w28671 and not w28672;
w28675 <= not w28673 and not w28674;
w28676 <= w28664 and not w28675;
w28677 <= w28664 and not w28676;
w28678 <= not w28675 and not w28676;
w28679 <= not w28677 and not w28678;
w28680 <= w3819 and w22282;
w28681 <= w3902 and w22288;
w28682 <= w3981 and w22285;
w28683 <= not w28681 and not w28682;
w28684 <= not w28680 and w28683;
w28685 <= w3985 and not w23594;
w28686 <= w28684 and not w28685;
w28687 <= a(26) and not w28686;
w28688 <= a(26) and not w28687;
w28689 <= not w28686 and not w28687;
w28690 <= not w28688 and not w28689;
w28691 <= not w28679 and not w28690;
w28692 <= not w28679 and not w28691;
w28693 <= not w28690 and not w28691;
w28694 <= not w28692 and not w28693;
w28695 <= not w28458 and not w28472;
w28696 <= w28694 and w28695;
w28697 <= not w28694 and not w28695;
w28698 <= not w28696 and not w28697;
w28699 <= w4629 and w22273;
w28700 <= w4468 and w22279;
w28701 <= w4539 and w22276;
w28702 <= not w28700 and not w28701;
w28703 <= not w28699 and w28702;
w28704 <= w4471 and not w24123;
w28705 <= w28703 and not w28704;
w28706 <= a(23) and not w28705;
w28707 <= a(23) and not w28706;
w28708 <= not w28705 and not w28706;
w28709 <= not w28707 and not w28708;
w28710 <= w28698 and not w28709;
w28711 <= w28698 and not w28710;
w28712 <= not w28709 and not w28710;
w28713 <= not w28711 and not w28712;
w28714 <= not w28478 and not w28491;
w28715 <= w28713 and w28714;
w28716 <= not w28713 and not w28714;
w28717 <= not w28715 and not w28716;
w28718 <= w5431 and w22264;
w28719 <= w4870 and w22270;
w28720 <= w5342 and w22267;
w28721 <= not w28719 and not w28720;
w28722 <= not w28718 and w28721;
w28723 <= w4873 and not w24568;
w28724 <= w28722 and not w28723;
w28725 <= a(20) and not w28724;
w28726 <= a(20) and not w28725;
w28727 <= not w28724 and not w28725;
w28728 <= not w28726 and not w28727;
w28729 <= w28717 and not w28728;
w28730 <= w28717 and not w28729;
w28731 <= not w28728 and not w28729;
w28732 <= not w28730 and not w28731;
w28733 <= not w28497 and not w28510;
w28734 <= w28732 and w28733;
w28735 <= not w28732 and not w28733;
w28736 <= not w28734 and not w28735;
w28737 <= w6168 and w22255;
w28738 <= w5598 and w22261;
w28739 <= w5874 and w22258;
w28740 <= not w28738 and not w28739;
w28741 <= not w28737 and w28740;
w28742 <= w5601 and not w25205;
w28743 <= w28741 and not w28742;
w28744 <= a(17) and not w28743;
w28745 <= a(17) and not w28744;
w28746 <= not w28743 and not w28744;
w28747 <= not w28745 and not w28746;
w28748 <= w28736 and not w28747;
w28749 <= w28736 and not w28748;
w28750 <= not w28747 and not w28748;
w28751 <= not w28749 and not w28750;
w28752 <= not w28516 and not w28529;
w28753 <= w28751 and w28752;
w28754 <= not w28751 and not w28752;
w28755 <= not w28753 and not w28754;
w28756 <= w7036 and w22244;
w28757 <= w6337 and w22247;
w28758 <= w6886 and w22250;
w28759 <= not w28757 and not w28758;
w28760 <= not w28756 and w28759;
w28761 <= w6332 and not w22464;
w28762 <= w28760 and not w28761;
w28763 <= a(14) and not w28762;
w28764 <= a(14) and not w28763;
w28765 <= not w28762 and not w28763;
w28766 <= not w28764 and not w28765;
w28767 <= w28755 and not w28766;
w28768 <= w28755 and not w28767;
w28769 <= not w28766 and not w28767;
w28770 <= not w28768 and not w28769;
w28771 <= not w28535 and not w28548;
w28772 <= w28770 and w28771;
w28773 <= not w28770 and not w28771;
w28774 <= not w28772 and not w28773;
w28775 <= w7918 and w25995;
w28776 <= w7226 and w25998;
w28777 <= w7567 and w26001;
w28778 <= not w28776 and not w28777;
w28779 <= not w28775 and w28778;
w28780 <= w7229 and not w26023;
w28781 <= w28779 and not w28780;
w28782 <= a(11) and not w28781;
w28783 <= a(11) and not w28782;
w28784 <= not w28781 and not w28782;
w28785 <= not w28783 and not w28784;
w28786 <= w28774 and not w28785;
w28787 <= w28774 and not w28786;
w28788 <= not w28785 and not w28786;
w28789 <= not w28787 and not w28788;
w28790 <= not w28554 and not w28567;
w28791 <= w28789 and w28790;
w28792 <= not w28789 and not w28790;
w28793 <= not w28791 and not w28792;
w28794 <= w9266 and w27377;
w28795 <= w8353 and w26825;
w28796 <= w8795 and w27108;
w28797 <= not w28795 and not w28796;
w28798 <= not w28794 and w28797;
w28799 <= w8356 and w27390;
w28800 <= w28798 and not w28799;
w28801 <= a(8) and not w28800;
w28802 <= a(8) and not w28801;
w28803 <= not w28800 and not w28801;
w28804 <= not w28802 and not w28803;
w28805 <= w28793 and not w28804;
w28806 <= w28793 and not w28805;
w28807 <= not w28804 and not w28805;
w28808 <= not w28806 and not w28807;
w28809 <= not w28573 and not w28586;
w28810 <= w28808 and w28809;
w28811 <= not w28808 and not w28809;
w28812 <= not w28810 and not w28811;
w28813 <= w6 and not w28143;
w28814 <= w9802 and w27633;
w28815 <= w10369 and w27899;
w28816 <= not w28814 and not w28815;
w28817 <= not w28813 and w28816;
w28818 <= w9805 and not w28158;
w28819 <= w28817 and not w28818;
w28820 <= a(5) and not w28819;
w28821 <= a(5) and not w28820;
w28822 <= not w28819 and not w28820;
w28823 <= not w28821 and not w28822;
w28824 <= w28812 and not w28823;
w28825 <= w28812 and not w28824;
w28826 <= not w28823 and not w28824;
w28827 <= not w28825 and not w28826;
w28828 <= not w28592 and not w28605;
w28829 <= w28827 and w28828;
w28830 <= not w28827 and not w28828;
w28831 <= not w28829 and not w28830;
w28832 <= not w28611 and not w28615;
w28833 <= not w28831 and w28832;
w28834 <= w28831 and not w28832;
w28835 <= not w28833 and not w28834;
w28836 <= w28617 and w28835;
w28837 <= not w28617 and not w28835;
w28838 <= not w28836 and not w28837;
w28839 <= w2359 and w15221;
w28840 <= w2639 and w28839;
w28841 <= w1038 and w28840;
w28842 <= w3620 and w28841;
w28843 <= w5134 and w28842;
w28844 <= w705 and w28843;
w28845 <= w350 and w28844;
w28846 <= w1117 and w28845;
w28847 <= w2378 and w28846;
w28848 <= w872 and w28847;
w28849 <= w2102 and w28848;
w28850 <= not w211 and w28849;
w28851 <= not w946 and w28850;
w28852 <= not w190 and w28851;
w28853 <= not w85 and w28852;
w28854 <= not w230 and w28853;
w28855 <= not w28431 and not w28854;
w28856 <= w28431 and w28854;
w28857 <= not w28647 and not w28856;
w28858 <= not w28855 and w28857;
w28859 <= not w28647 and not w28858;
w28860 <= not w28855 and not w28858;
w28861 <= not w28856 and w28860;
w28862 <= not w28859 and not w28861;
w28863 <= w10 and not w23255;
w28864 <= w2955 and w22297;
w28865 <= w2958 and w22303;
w28866 <= w2963 and w22300;
w28867 <= not w28865 and not w28866;
w28868 <= not w28864 and w28867;
w28869 <= not w28863 and w28868;
w28870 <= not w28862 and not w28869;
w28871 <= not w28862 and not w28870;
w28872 <= not w28869 and not w28870;
w28873 <= not w28871 and not w28872;
w28874 <= not w28657 and not w28663;
w28875 <= w28873 and w28874;
w28876 <= not w28873 and not w28874;
w28877 <= not w28875 and not w28876;
w28878 <= w3392 and w22288;
w28879 <= w3477 and w22294;
w28880 <= w3541 and w22291;
w28881 <= not w28879 and not w28880;
w28882 <= not w28878 and w28881;
w28883 <= w3303 and not w22491;
w28884 <= w28882 and not w28883;
w28885 <= a(29) and not w28884;
w28886 <= a(29) and not w28885;
w28887 <= not w28884 and not w28885;
w28888 <= not w28886 and not w28887;
w28889 <= w28877 and not w28888;
w28890 <= w28877 and not w28889;
w28891 <= not w28888 and not w28889;
w28892 <= not w28890 and not w28891;
w28893 <= w3819 and w22279;
w28894 <= w3902 and w22285;
w28895 <= w3981 and w22282;
w28896 <= not w28894 and not w28895;
w28897 <= not w28893 and w28896;
w28898 <= w3985 and not w23577;
w28899 <= w28897 and not w28898;
w28900 <= a(26) and not w28899;
w28901 <= a(26) and not w28900;
w28902 <= not w28899 and not w28900;
w28903 <= not w28901 and not w28902;
w28904 <= not w28892 and not w28903;
w28905 <= not w28892 and not w28904;
w28906 <= not w28903 and not w28904;
w28907 <= not w28905 and not w28906;
w28908 <= not w28676 and not w28691;
w28909 <= w28907 and w28908;
w28910 <= not w28907 and not w28908;
w28911 <= not w28909 and not w28910;
w28912 <= w4629 and w22270;
w28913 <= w4468 and w22276;
w28914 <= w4539 and w22273;
w28915 <= not w28913 and not w28914;
w28916 <= not w28912 and w28915;
w28917 <= w4471 and not w24102;
w28918 <= w28916 and not w28917;
w28919 <= a(23) and not w28918;
w28920 <= a(23) and not w28919;
w28921 <= not w28918 and not w28919;
w28922 <= not w28920 and not w28921;
w28923 <= w28911 and not w28922;
w28924 <= w28911 and not w28923;
w28925 <= not w28922 and not w28923;
w28926 <= not w28924 and not w28925;
w28927 <= not w28697 and not w28710;
w28928 <= w28926 and w28927;
w28929 <= not w28926 and not w28927;
w28930 <= not w28928 and not w28929;
w28931 <= w5431 and w22261;
w28932 <= w4870 and w22267;
w28933 <= w5342 and w22264;
w28934 <= not w28932 and not w28933;
w28935 <= not w28931 and w28934;
w28936 <= w4873 and not w24551;
w28937 <= w28935 and not w28936;
w28938 <= a(20) and not w28937;
w28939 <= a(20) and not w28938;
w28940 <= not w28937 and not w28938;
w28941 <= not w28939 and not w28940;
w28942 <= w28930 and not w28941;
w28943 <= w28930 and not w28942;
w28944 <= not w28941 and not w28942;
w28945 <= not w28943 and not w28944;
w28946 <= not w28716 and not w28729;
w28947 <= w28945 and w28946;
w28948 <= not w28945 and not w28946;
w28949 <= not w28947 and not w28948;
w28950 <= w6168 and w22247;
w28951 <= w5598 and w22258;
w28952 <= w5874 and w22255;
w28953 <= not w28951 and not w28952;
w28954 <= not w28950 and w28953;
w28955 <= w5601 and not w25250;
w28956 <= w28954 and not w28955;
w28957 <= a(17) and not w28956;
w28958 <= a(17) and not w28957;
w28959 <= not w28956 and not w28957;
w28960 <= not w28958 and not w28959;
w28961 <= w28949 and not w28960;
w28962 <= w28949 and not w28961;
w28963 <= not w28960 and not w28961;
w28964 <= not w28962 and not w28963;
w28965 <= not w28735 and not w28748;
w28966 <= w28964 and w28965;
w28967 <= not w28964 and not w28965;
w28968 <= not w28966 and not w28967;
w28969 <= w7036 and w25998;
w28970 <= w6337 and w22250;
w28971 <= w6886 and w22244;
w28972 <= not w28970 and not w28971;
w28973 <= not w28969 and w28972;
w28974 <= w6332 and not w26539;
w28975 <= w28973 and not w28974;
w28976 <= a(14) and not w28975;
w28977 <= a(14) and not w28976;
w28978 <= not w28975 and not w28976;
w28979 <= not w28977 and not w28978;
w28980 <= w28968 and not w28979;
w28981 <= w28968 and not w28980;
w28982 <= not w28979 and not w28980;
w28983 <= not w28981 and not w28982;
w28984 <= not w28754 and not w28767;
w28985 <= w28983 and w28984;
w28986 <= not w28983 and not w28984;
w28987 <= not w28985 and not w28986;
w28988 <= w7918 and w26825;
w28989 <= w7226 and w26001;
w28990 <= w7567 and w25995;
w28991 <= not w28989 and not w28990;
w28992 <= not w28988 and w28991;
w28993 <= w7229 and not w26839;
w28994 <= w28992 and not w28993;
w28995 <= a(11) and not w28994;
w28996 <= a(11) and not w28995;
w28997 <= not w28994 and not w28995;
w28998 <= not w28996 and not w28997;
w28999 <= w28987 and not w28998;
w29000 <= w28987 and not w28999;
w29001 <= not w28998 and not w28999;
w29002 <= not w29000 and not w29001;
w29003 <= not w28773 and not w28786;
w29004 <= w29002 and w29003;
w29005 <= not w29002 and not w29003;
w29006 <= not w29004 and not w29005;
w29007 <= w9266 and w27633;
w29008 <= w8353 and w27108;
w29009 <= w8795 and w27377;
w29010 <= not w29008 and not w29009;
w29011 <= not w29007 and w29010;
w29012 <= w8356 and not w27648;
w29013 <= w29011 and not w29012;
w29014 <= a(8) and not w29013;
w29015 <= a(8) and not w29014;
w29016 <= not w29013 and not w29014;
w29017 <= not w29015 and not w29016;
w29018 <= w29006 and not w29017;
w29019 <= w29006 and not w29018;
w29020 <= not w29017 and not w29018;
w29021 <= not w29019 and not w29020;
w29022 <= not w28792 and not w28805;
w29023 <= not w15011 and not w28143;
w29024 <= w9802 and w27899;
w29025 <= not w29023 and not w29024;
w29026 <= not w9805 and w29025;
w29027 <= w28156 and w29025;
w29028 <= not w29026 and not w29027;
w29029 <= a(5) and not w29028;
w29030 <= not a(5) and w29028;
w29031 <= not w29029 and not w29030;
w29032 <= not w29022 and not w29031;
w29033 <= w29022 and w29031;
w29034 <= not w29032 and not w29033;
w29035 <= not w29021 and w29034;
w29036 <= not w29021 and not w29035;
w29037 <= w29034 and not w29035;
w29038 <= not w29036 and not w29037;
w29039 <= not w28811 and not w28824;
w29040 <= w29038 and w29039;
w29041 <= not w29038 and not w29039;
w29042 <= not w29040 and not w29041;
w29043 <= not w28830 and not w28834;
w29044 <= not w29042 and w29043;
w29045 <= w29042 and not w29043;
w29046 <= not w29044 and not w29045;
w29047 <= w28836 and w29046;
w29048 <= not w28836 and not w29046;
w29049 <= not w29047 and not w29048;
w29050 <= not w29041 and not w29045;
w29051 <= not w29032 and not w29035;
w29052 <= not w28870 and not w28876;
w29053 <= w1794 and w4270;
w29054 <= w1008 and w29053;
w29055 <= w4292 and w29054;
w29056 <= w895 and w29055;
w29057 <= w461 and w29056;
w29058 <= w13761 and w29057;
w29059 <= w2992 and w29058;
w29060 <= w2402 and w29059;
w29061 <= w3821 and w29060;
w29062 <= w1696 and w29061;
w29063 <= w22683 and w29062;
w29064 <= not w681 and w29063;
w29065 <= not w215 and w29064;
w29066 <= not w54 and w29065;
w29067 <= not w293 and w29066;
w29068 <= w28431 and w29067;
w29069 <= not w28431 and not w29067;
w29070 <= not w29068 and not w29069;
w29071 <= not w15013 and not w28143;
w29072 <= not a(5) and w29071;
w29073 <= a(5) and not w29071;
w29074 <= not w29070 and not w29073;
w29075 <= not w29072 and w29074;
w29076 <= not w29070 and not w29075;
w29077 <= not w29073 and not w29075;
w29078 <= not w29072 and w29077;
w29079 <= not w29076 and not w29078;
w29080 <= not w28860 and w29079;
w29081 <= w28860 and not w29079;
w29082 <= not w29080 and not w29081;
w29083 <= w10 and w23303;
w29084 <= w2955 and w22294;
w29085 <= w2958 and w22300;
w29086 <= w2963 and w22297;
w29087 <= not w29085 and not w29086;
w29088 <= not w29084 and w29087;
w29089 <= not w29083 and w29088;
w29090 <= not w29082 and not w29089;
w29091 <= w29082 and w29089;
w29092 <= not w29090 and not w29091;
w29093 <= w29052 and not w29092;
w29094 <= not w29052 and w29092;
w29095 <= not w29093 and not w29094;
w29096 <= w3392 and w22285;
w29097 <= w3477 and w22291;
w29098 <= w3541 and w22288;
w29099 <= not w29097 and not w29098;
w29100 <= not w29096 and w29099;
w29101 <= w3303 and w23607;
w29102 <= w29100 and not w29101;
w29103 <= a(29) and not w29102;
w29104 <= a(29) and not w29103;
w29105 <= not w29102 and not w29103;
w29106 <= not w29104 and not w29105;
w29107 <= w29095 and not w29106;
w29108 <= w29095 and not w29107;
w29109 <= not w29106 and not w29107;
w29110 <= not w29108 and not w29109;
w29111 <= w3819 and w22276;
w29112 <= w3902 and w22282;
w29113 <= w3981 and w22279;
w29114 <= not w29112 and not w29113;
w29115 <= not w29111 and w29114;
w29116 <= w3985 and w24077;
w29117 <= w29115 and not w29116;
w29118 <= a(26) and not w29117;
w29119 <= a(26) and not w29118;
w29120 <= not w29117 and not w29118;
w29121 <= not w29119 and not w29120;
w29122 <= not w29110 and not w29121;
w29123 <= not w29110 and not w29122;
w29124 <= not w29121 and not w29122;
w29125 <= not w29123 and not w29124;
w29126 <= not w28889 and not w28904;
w29127 <= w29125 and w29126;
w29128 <= not w29125 and not w29126;
w29129 <= not w29127 and not w29128;
w29130 <= w4629 and w22267;
w29131 <= w4468 and w22273;
w29132 <= w4539 and w22270;
w29133 <= not w29131 and not w29132;
w29134 <= not w29130 and w29133;
w29135 <= w4471 and w22477;
w29136 <= w29134 and not w29135;
w29137 <= a(23) and not w29136;
w29138 <= a(23) and not w29137;
w29139 <= not w29136 and not w29137;
w29140 <= not w29138 and not w29139;
w29141 <= w29129 and not w29140;
w29142 <= w29129 and not w29141;
w29143 <= not w29140 and not w29141;
w29144 <= not w29142 and not w29143;
w29145 <= not w28910 and not w28923;
w29146 <= w29144 and w29145;
w29147 <= not w29144 and not w29145;
w29148 <= not w29146 and not w29147;
w29149 <= w5431 and w22258;
w29150 <= w4870 and w22264;
w29151 <= w5342 and w22261;
w29152 <= not w29150 and not w29151;
w29153 <= not w29149 and w29152;
w29154 <= w4873 and w24534;
w29155 <= w29153 and not w29154;
w29156 <= a(20) and not w29155;
w29157 <= a(20) and not w29156;
w29158 <= not w29155 and not w29156;
w29159 <= not w29157 and not w29158;
w29160 <= w29148 and not w29159;
w29161 <= w29148 and not w29160;
w29162 <= not w29159 and not w29160;
w29163 <= not w29161 and not w29162;
w29164 <= not w28929 and not w28942;
w29165 <= w29163 and w29164;
w29166 <= not w29163 and not w29164;
w29167 <= not w29165 and not w29166;
w29168 <= w6168 and w22250;
w29169 <= w5598 and w22255;
w29170 <= w5874 and w22247;
w29171 <= not w29169 and not w29170;
w29172 <= not w29168 and w29171;
w29173 <= w5601 and w25229;
w29174 <= w29172 and not w29173;
w29175 <= a(17) and not w29174;
w29176 <= a(17) and not w29175;
w29177 <= not w29174 and not w29175;
w29178 <= not w29176 and not w29177;
w29179 <= w29167 and not w29178;
w29180 <= w29167 and not w29179;
w29181 <= not w29178 and not w29179;
w29182 <= not w29180 and not w29181;
w29183 <= not w28948 and not w28961;
w29184 <= w29182 and w29183;
w29185 <= not w29182 and not w29183;
w29186 <= not w29184 and not w29185;
w29187 <= not w28967 and not w28980;
w29188 <= w7036 and w26001;
w29189 <= w6337 and w22244;
w29190 <= w6886 and w25998;
w29191 <= not w29189 and not w29190;
w29192 <= not w29188 and w29191;
w29193 <= w6332 and not w26559;
w29194 <= w29192 and not w29193;
w29195 <= a(14) and not w29194;
w29196 <= a(14) and not w29195;
w29197 <= not w29194 and not w29195;
w29198 <= not w29196 and not w29197;
w29199 <= not w29187 and not w29198;
w29200 <= not w29187 and not w29199;
w29201 <= not w29198 and not w29199;
w29202 <= not w29200 and not w29201;
w29203 <= not w29186 and w29202;
w29204 <= w29186 and not w29202;
w29205 <= not w29203 and not w29204;
w29206 <= w7918 and w27108;
w29207 <= w7226 and w25995;
w29208 <= w7567 and w26825;
w29209 <= not w29207 and not w29208;
w29210 <= not w29206 and w29209;
w29211 <= w7229 and w27120;
w29212 <= w29210 and not w29211;
w29213 <= a(11) and not w29212;
w29214 <= a(11) and not w29213;
w29215 <= not w29212 and not w29213;
w29216 <= not w29214 and not w29215;
w29217 <= w29205 and not w29216;
w29218 <= w29205 and not w29217;
w29219 <= not w29216 and not w29217;
w29220 <= not w29218 and not w29219;
w29221 <= not w28986 and not w28999;
w29222 <= w29220 and w29221;
w29223 <= not w29220 and not w29221;
w29224 <= not w29222 and not w29223;
w29225 <= not w29005 and not w29018;
w29226 <= w9266 and w27899;
w29227 <= w8353 and w27377;
w29228 <= w8795 and w27633;
w29229 <= not w29227 and not w29228;
w29230 <= not w29226 and w29229;
w29231 <= w8356 and w27911;
w29232 <= w29230 and not w29231;
w29233 <= a(8) and not w29232;
w29234 <= a(8) and not w29233;
w29235 <= not w29232 and not w29233;
w29236 <= not w29234 and not w29235;
w29237 <= not w29225 and not w29236;
w29238 <= not w29225 and not w29237;
w29239 <= not w29236 and not w29237;
w29240 <= not w29238 and not w29239;
w29241 <= not w29224 and w29240;
w29242 <= w29224 and not w29240;
w29243 <= not w29241 and not w29242;
w29244 <= not w29051 and w29243;
w29245 <= w29051 and not w29243;
w29246 <= not w29244 and not w29245;
w29247 <= not w29050 and w29246;
w29248 <= w29050 and not w29246;
w29249 <= not w29247 and not w29248;
w29250 <= not w29047 and not w29249;
w29251 <= w29047 and w29249;
w29252 <= not w29250 and not w29251;
w29253 <= not w29094 and not w29107;
w29254 <= w10 and not w23280;
w29255 <= w2955 and w22291;
w29256 <= w2958 and w22297;
w29257 <= w2963 and w22294;
w29258 <= not w29256 and not w29257;
w29259 <= not w29255 and w29258;
w29260 <= not w29254 and w29259;
w29261 <= w1259 and w5991;
w29262 <= w1141 and w29261;
w29263 <= w1281 and w29262;
w29264 <= w6640 and w29263;
w29265 <= w589 and w29264;
w29266 <= w3405 and w29265;
w29267 <= w804 and w29266;
w29268 <= w1076 and w29267;
w29269 <= not w164 and w29268;
w29270 <= not w56 and w29269;
w29271 <= not w183 and w29270;
w29272 <= not w141 and w29271;
w29273 <= w1667 and w2198;
w29274 <= w3095 and w29273;
w29275 <= w6706 and w29274;
w29276 <= w29272 and w29275;
w29277 <= w1313 and w29276;
w29278 <= w2613 and w29277;
w29279 <= w535 and w29278;
w29280 <= w423 and w29279;
w29281 <= w944 and w29280;
w29282 <= w1760 and w29281;
w29283 <= w1457 and w29282;
w29284 <= not w946 and w29283;
w29285 <= not w1181 and w29284;
w29286 <= not w210 and w29285;
w29287 <= not w292 and w29286;
w29288 <= not w100 and w29287;
w29289 <= not w428 and w29288;
w29290 <= not w590 and w29289;
w29291 <= w28431 and not w29067;
w29292 <= not w29075 and not w29291;
w29293 <= w29290 and not w29292;
w29294 <= not w29290 and w29292;
w29295 <= not w29293 and not w29294;
w29296 <= not w29260 and w29295;
w29297 <= not w29260 and not w29296;
w29298 <= w29295 and not w29296;
w29299 <= not w29297 and not w29298;
w29300 <= not w28860 and not w29079;
w29301 <= not w29090 and not w29300;
w29302 <= w29299 and w29301;
w29303 <= not w29299 and not w29301;
w29304 <= not w29302 and not w29303;
w29305 <= w3392 and w22282;
w29306 <= w3477 and w22288;
w29307 <= w3541 and w22285;
w29308 <= not w29306 and not w29307;
w29309 <= not w29305 and w29308;
w29310 <= not w3303 and w29309;
w29311 <= w23594 and w29309;
w29312 <= not w29310 and not w29311;
w29313 <= a(29) and not w29312;
w29314 <= not a(29) and w29312;
w29315 <= not w29313 and not w29314;
w29316 <= w29304 and not w29315;
w29317 <= not w29304 and w29315;
w29318 <= not w29316 and not w29317;
w29319 <= not w29253 and w29318;
w29320 <= w29253 and not w29318;
w29321 <= not w29319 and not w29320;
w29322 <= w3819 and w22273;
w29323 <= w3902 and w22279;
w29324 <= w3981 and w22276;
w29325 <= not w29323 and not w29324;
w29326 <= not w29322 and w29325;
w29327 <= w3985 and not w24123;
w29328 <= w29326 and not w29327;
w29329 <= a(26) and not w29328;
w29330 <= a(26) and not w29329;
w29331 <= not w29328 and not w29329;
w29332 <= not w29330 and not w29331;
w29333 <= w29321 and not w29332;
w29334 <= w29321 and not w29333;
w29335 <= not w29332 and not w29333;
w29336 <= not w29334 and not w29335;
w29337 <= not w29122 and not w29128;
w29338 <= w29336 and w29337;
w29339 <= not w29336 and not w29337;
w29340 <= not w29338 and not w29339;
w29341 <= w4629 and w22264;
w29342 <= w4468 and w22270;
w29343 <= w4539 and w22267;
w29344 <= not w29342 and not w29343;
w29345 <= not w29341 and w29344;
w29346 <= w4471 and not w24568;
w29347 <= w29345 and not w29346;
w29348 <= a(23) and not w29347;
w29349 <= a(23) and not w29348;
w29350 <= not w29347 and not w29348;
w29351 <= not w29349 and not w29350;
w29352 <= w29340 and not w29351;
w29353 <= w29340 and not w29352;
w29354 <= not w29351 and not w29352;
w29355 <= not w29353 and not w29354;
w29356 <= not w29141 and not w29147;
w29357 <= w29355 and w29356;
w29358 <= not w29355 and not w29356;
w29359 <= not w29357 and not w29358;
w29360 <= w5431 and w22255;
w29361 <= w4870 and w22261;
w29362 <= w5342 and w22258;
w29363 <= not w29361 and not w29362;
w29364 <= not w29360 and w29363;
w29365 <= w4873 and not w25205;
w29366 <= w29364 and not w29365;
w29367 <= a(20) and not w29366;
w29368 <= a(20) and not w29367;
w29369 <= not w29366 and not w29367;
w29370 <= not w29368 and not w29369;
w29371 <= w29359 and not w29370;
w29372 <= w29359 and not w29371;
w29373 <= not w29370 and not w29371;
w29374 <= not w29372 and not w29373;
w29375 <= not w29160 and not w29166;
w29376 <= w29374 and w29375;
w29377 <= not w29374 and not w29375;
w29378 <= not w29376 and not w29377;
w29379 <= w6168 and w22244;
w29380 <= w5598 and w22247;
w29381 <= w5874 and w22250;
w29382 <= not w29380 and not w29381;
w29383 <= not w29379 and w29382;
w29384 <= w5601 and not w22464;
w29385 <= w29383 and not w29384;
w29386 <= a(17) and not w29385;
w29387 <= a(17) and not w29386;
w29388 <= not w29385 and not w29386;
w29389 <= not w29387 and not w29388;
w29390 <= w29378 and not w29389;
w29391 <= w29378 and not w29390;
w29392 <= not w29389 and not w29390;
w29393 <= not w29391 and not w29392;
w29394 <= not w29179 and not w29185;
w29395 <= w29393 and w29394;
w29396 <= not w29393 and not w29394;
w29397 <= not w29395 and not w29396;
w29398 <= w7036 and w25995;
w29399 <= w6337 and w25998;
w29400 <= w6886 and w26001;
w29401 <= not w29399 and not w29400;
w29402 <= not w29398 and w29401;
w29403 <= w6332 and not w26023;
w29404 <= w29402 and not w29403;
w29405 <= a(14) and not w29404;
w29406 <= a(14) and not w29405;
w29407 <= not w29404 and not w29405;
w29408 <= not w29406 and not w29407;
w29409 <= w29397 and not w29408;
w29410 <= w29397 and not w29409;
w29411 <= not w29408 and not w29409;
w29412 <= not w29410 and not w29411;
w29413 <= not w29199 and not w29204;
w29414 <= not w29412 and not w29413;
w29415 <= not w29412 and not w29414;
w29416 <= not w29413 and not w29414;
w29417 <= not w29415 and not w29416;
w29418 <= w7918 and w27377;
w29419 <= w7226 and w26825;
w29420 <= w7567 and w27108;
w29421 <= not w29419 and not w29420;
w29422 <= not w29418 and w29421;
w29423 <= w7229 and w27390;
w29424 <= w29422 and not w29423;
w29425 <= a(11) and not w29424;
w29426 <= a(11) and not w29425;
w29427 <= not w29424 and not w29425;
w29428 <= not w29426 and not w29427;
w29429 <= not w29417 and not w29428;
w29430 <= not w29417 and not w29429;
w29431 <= not w29428 and not w29429;
w29432 <= not w29430 and not w29431;
w29433 <= not w29217 and not w29223;
w29434 <= w29432 and w29433;
w29435 <= not w29432 and not w29433;
w29436 <= not w29434 and not w29435;
w29437 <= w9266 and not w28143;
w29438 <= w8353 and w27633;
w29439 <= w8795 and w27899;
w29440 <= not w29438 and not w29439;
w29441 <= not w29437 and w29440;
w29442 <= w8356 and not w28158;
w29443 <= w29441 and not w29442;
w29444 <= a(8) and not w29443;
w29445 <= a(8) and not w29444;
w29446 <= not w29443 and not w29444;
w29447 <= not w29445 and not w29446;
w29448 <= w29436 and not w29447;
w29449 <= w29436 and not w29448;
w29450 <= not w29447 and not w29448;
w29451 <= not w29449 and not w29450;
w29452 <= not w29237 and not w29242;
w29453 <= not w29451 and not w29452;
w29454 <= not w29451 and not w29453;
w29455 <= not w29452 and not w29453;
w29456 <= not w29454 and not w29455;
w29457 <= not w29244 and not w29247;
w29458 <= w29456 and w29457;
w29459 <= not w29456 and not w29457;
w29460 <= not w29458 and not w29459;
w29461 <= not w29251 and w29460;
w29462 <= w29251 and not w29460;
w29463 <= not w29461 and not w29462;
w29464 <= w29251 and w29460;
w29465 <= not w29293 and not w29296;
w29466 <= not w110 and not w190;
w29467 <= not w234 and w29466;
w29468 <= not w240 and w29467;
w29469 <= not w427 and w29468;
w29470 <= not w100 and w29469;
w29471 <= not w527 and w29470;
w29472 <= not w607 and w29471;
w29473 <= not w205 and w29472;
w29474 <= w2377 and w12647;
w29475 <= w875 and w29474;
w29476 <= w4230 and w29475;
w29477 <= w2341 and w29476;
w29478 <= w981 and w29477;
w29479 <= w2352 and w29478;
w29480 <= w820 and w29479;
w29481 <= not w224 and w29480;
w29482 <= not w90 and w29481;
w29483 <= not w99 and w29482;
w29484 <= not w126 and w29483;
w29485 <= not w180 and w29484;
w29486 <= w12846 and w13743;
w29487 <= w6483 and w29486;
w29488 <= w29485 and w29487;
w29489 <= w29473 and w29488;
w29490 <= w3000 and w29489;
w29491 <= w12331 and w29490;
w29492 <= not w129 and w29491;
w29493 <= not w189 and w29492;
w29494 <= not w370 and w29493;
w29495 <= not w178 and w29494;
w29496 <= not w401 and w29495;
w29497 <= not w472 and w29496;
w29498 <= not w267 and w29497;
w29499 <= not w260 and w29498;
w29500 <= not w29290 and w29499;
w29501 <= w29290 and not w29499;
w29502 <= not w29465 and not w29501;
w29503 <= not w29500 and w29502;
w29504 <= not w29465 and not w29503;
w29505 <= not w29501 and not w29503;
w29506 <= not w29500 and w29505;
w29507 <= not w29504 and not w29506;
w29508 <= w10 and not w22491;
w29509 <= w2955 and w22288;
w29510 <= w2958 and w22294;
w29511 <= w2963 and w22291;
w29512 <= not w29510 and not w29511;
w29513 <= not w29509 and w29512;
w29514 <= not w29508 and w29513;
w29515 <= not w29507 and not w29514;
w29516 <= not w29507 and not w29515;
w29517 <= not w29514 and not w29515;
w29518 <= not w29516 and not w29517;
w29519 <= not w29303 and not w29316;
w29520 <= w29518 and w29519;
w29521 <= not w29518 and not w29519;
w29522 <= not w29520 and not w29521;
w29523 <= w3392 and w22279;
w29524 <= w3477 and w22285;
w29525 <= w3541 and w22282;
w29526 <= not w29524 and not w29525;
w29527 <= not w29523 and w29526;
w29528 <= w3303 and not w23577;
w29529 <= w29527 and not w29528;
w29530 <= a(29) and not w29529;
w29531 <= a(29) and not w29530;
w29532 <= not w29529 and not w29530;
w29533 <= not w29531 and not w29532;
w29534 <= w29522 and not w29533;
w29535 <= w29522 and not w29534;
w29536 <= not w29533 and not w29534;
w29537 <= not w29535 and not w29536;
w29538 <= w3819 and w22270;
w29539 <= w3902 and w22276;
w29540 <= w3981 and w22273;
w29541 <= not w29539 and not w29540;
w29542 <= not w29538 and w29541;
w29543 <= w3985 and not w24102;
w29544 <= w29542 and not w29543;
w29545 <= a(26) and not w29544;
w29546 <= a(26) and not w29545;
w29547 <= not w29544 and not w29545;
w29548 <= not w29546 and not w29547;
w29549 <= not w29537 and not w29548;
w29550 <= not w29537 and not w29549;
w29551 <= not w29548 and not w29549;
w29552 <= not w29550 and not w29551;
w29553 <= not w29319 and not w29333;
w29554 <= w29552 and w29553;
w29555 <= not w29552 and not w29553;
w29556 <= not w29554 and not w29555;
w29557 <= w4629 and w22261;
w29558 <= w4468 and w22267;
w29559 <= w4539 and w22264;
w29560 <= not w29558 and not w29559;
w29561 <= not w29557 and w29560;
w29562 <= w4471 and not w24551;
w29563 <= w29561 and not w29562;
w29564 <= a(23) and not w29563;
w29565 <= a(23) and not w29564;
w29566 <= not w29563 and not w29564;
w29567 <= not w29565 and not w29566;
w29568 <= w29556 and not w29567;
w29569 <= w29556 and not w29568;
w29570 <= not w29567 and not w29568;
w29571 <= not w29569 and not w29570;
w29572 <= not w29339 and not w29352;
w29573 <= w29571 and w29572;
w29574 <= not w29571 and not w29572;
w29575 <= not w29573 and not w29574;
w29576 <= w5431 and w22247;
w29577 <= w4870 and w22258;
w29578 <= w5342 and w22255;
w29579 <= not w29577 and not w29578;
w29580 <= not w29576 and w29579;
w29581 <= w4873 and not w25250;
w29582 <= w29580 and not w29581;
w29583 <= a(20) and not w29582;
w29584 <= a(20) and not w29583;
w29585 <= not w29582 and not w29583;
w29586 <= not w29584 and not w29585;
w29587 <= w29575 and not w29586;
w29588 <= w29575 and not w29587;
w29589 <= not w29586 and not w29587;
w29590 <= not w29588 and not w29589;
w29591 <= not w29358 and not w29371;
w29592 <= w29590 and w29591;
w29593 <= not w29590 and not w29591;
w29594 <= not w29592 and not w29593;
w29595 <= w6168 and w25998;
w29596 <= w5598 and w22250;
w29597 <= w5874 and w22244;
w29598 <= not w29596 and not w29597;
w29599 <= not w29595 and w29598;
w29600 <= w5601 and not w26539;
w29601 <= w29599 and not w29600;
w29602 <= a(17) and not w29601;
w29603 <= a(17) and not w29602;
w29604 <= not w29601 and not w29602;
w29605 <= not w29603 and not w29604;
w29606 <= w29594 and not w29605;
w29607 <= w29594 and not w29606;
w29608 <= not w29605 and not w29606;
w29609 <= not w29607 and not w29608;
w29610 <= not w29377 and not w29390;
w29611 <= w29609 and w29610;
w29612 <= not w29609 and not w29610;
w29613 <= not w29611 and not w29612;
w29614 <= w7036 and w26825;
w29615 <= w6337 and w26001;
w29616 <= w6886 and w25995;
w29617 <= not w29615 and not w29616;
w29618 <= not w29614 and w29617;
w29619 <= w6332 and not w26839;
w29620 <= w29618 and not w29619;
w29621 <= a(14) and not w29620;
w29622 <= a(14) and not w29621;
w29623 <= not w29620 and not w29621;
w29624 <= not w29622 and not w29623;
w29625 <= w29613 and not w29624;
w29626 <= w29613 and not w29625;
w29627 <= not w29624 and not w29625;
w29628 <= not w29626 and not w29627;
w29629 <= not w29396 and not w29409;
w29630 <= w29628 and w29629;
w29631 <= not w29628 and not w29629;
w29632 <= not w29630 and not w29631;
w29633 <= w7918 and w27633;
w29634 <= w7226 and w27108;
w29635 <= w7567 and w27377;
w29636 <= not w29634 and not w29635;
w29637 <= not w29633 and w29636;
w29638 <= w7229 and not w27648;
w29639 <= w29637 and not w29638;
w29640 <= a(11) and not w29639;
w29641 <= a(11) and not w29640;
w29642 <= not w29639 and not w29640;
w29643 <= not w29641 and not w29642;
w29644 <= w29632 and not w29643;
w29645 <= w29632 and not w29644;
w29646 <= not w29643 and not w29644;
w29647 <= not w29645 and not w29646;
w29648 <= not w29414 and not w29429;
w29649 <= not w14525 and not w28143;
w29650 <= w8353 and w27899;
w29651 <= not w29649 and not w29650;
w29652 <= not w8356 and w29651;
w29653 <= w28156 and w29651;
w29654 <= not w29652 and not w29653;
w29655 <= a(8) and not w29654;
w29656 <= not a(8) and w29654;
w29657 <= not w29655 and not w29656;
w29658 <= not w29648 and not w29657;
w29659 <= w29648 and w29657;
w29660 <= not w29658 and not w29659;
w29661 <= not w29647 and w29660;
w29662 <= not w29647 and not w29661;
w29663 <= w29660 and not w29661;
w29664 <= not w29662 and not w29663;
w29665 <= not w29435 and not w29448;
w29666 <= w29664 and w29665;
w29667 <= not w29664 and not w29665;
w29668 <= not w29666 and not w29667;
w29669 <= not w29453 and not w29459;
w29670 <= not w29668 and w29669;
w29671 <= w29668 and not w29669;
w29672 <= not w29670 and not w29671;
w29673 <= w29464 and w29672;
w29674 <= not w29464 and not w29672;
w29675 <= not w29673 and not w29674;
w29676 <= not w29667 and not w29671;
w29677 <= not w29658 and not w29661;
w29678 <= w10 and w23607;
w29679 <= w2955 and w22285;
w29680 <= w2958 and w22291;
w29681 <= w2963 and w22288;
w29682 <= not w29680 and not w29681;
w29683 <= not w29679 and w29682;
w29684 <= not w29678 and w29683;
w29685 <= not w14527 and not w28143;
w29686 <= a(8) and not w29685;
w29687 <= not a(8) and w29685;
w29688 <= not w29686 and not w29687;
w29689 <= w895 and w3409;
w29690 <= w1357 and w29689;
w29691 <= w235 and w29690;
w29692 <= w13708 and w29691;
w29693 <= w1941 and w29692;
w29694 <= w1510 and w29693;
w29695 <= w2632 and w29694;
w29696 <= w170 and w29695;
w29697 <= w2893 and w29696;
w29698 <= w2419 and w29697;
w29699 <= w2105 and w29698;
w29700 <= w91 and w29699;
w29701 <= not w648 and w29700;
w29702 <= not w303 and w29701;
w29703 <= w29290 and w29702;
w29704 <= not w29290 and not w29702;
w29705 <= not w29703 and not w29704;
w29706 <= w29688 and w29705;
w29707 <= not w29688 and not w29705;
w29708 <= not w29706 and not w29707;
w29709 <= not w29505 and w29708;
w29710 <= w29505 and not w29708;
w29711 <= not w29709 and not w29710;
w29712 <= not w29684 and w29711;
w29713 <= w29711 and not w29712;
w29714 <= not w29684 and not w29712;
w29715 <= not w29713 and not w29714;
w29716 <= w3392 and w22276;
w29717 <= w3477 and w22282;
w29718 <= w3541 and w22279;
w29719 <= not w29717 and not w29718;
w29720 <= not w29716 and w29719;
w29721 <= w3303 and w24077;
w29722 <= w29720 and not w29721;
w29723 <= a(29) and not w29722;
w29724 <= a(29) and not w29723;
w29725 <= not w29722 and not w29723;
w29726 <= not w29724 and not w29725;
w29727 <= not w29715 and not w29726;
w29728 <= not w29715 and not w29727;
w29729 <= not w29726 and not w29727;
w29730 <= not w29728 and not w29729;
w29731 <= not w29515 and not w29521;
w29732 <= w29730 and w29731;
w29733 <= not w29730 and not w29731;
w29734 <= not w29732 and not w29733;
w29735 <= w3819 and w22267;
w29736 <= w3902 and w22273;
w29737 <= w3981 and w22270;
w29738 <= not w29736 and not w29737;
w29739 <= not w29735 and w29738;
w29740 <= w3985 and w22477;
w29741 <= w29739 and not w29740;
w29742 <= a(26) and not w29741;
w29743 <= a(26) and not w29742;
w29744 <= not w29741 and not w29742;
w29745 <= not w29743 and not w29744;
w29746 <= w29734 and not w29745;
w29747 <= w29734 and not w29746;
w29748 <= not w29745 and not w29746;
w29749 <= not w29747 and not w29748;
w29750 <= not w29534 and not w29549;
w29751 <= w29749 and w29750;
w29752 <= not w29749 and not w29750;
w29753 <= not w29751 and not w29752;
w29754 <= w4629 and w22258;
w29755 <= w4468 and w22264;
w29756 <= w4539 and w22261;
w29757 <= not w29755 and not w29756;
w29758 <= not w29754 and w29757;
w29759 <= w4471 and w24534;
w29760 <= w29758 and not w29759;
w29761 <= a(23) and not w29760;
w29762 <= a(23) and not w29761;
w29763 <= not w29760 and not w29761;
w29764 <= not w29762 and not w29763;
w29765 <= w29753 and not w29764;
w29766 <= w29753 and not w29765;
w29767 <= not w29764 and not w29765;
w29768 <= not w29766 and not w29767;
w29769 <= not w29555 and not w29568;
w29770 <= w29768 and w29769;
w29771 <= not w29768 and not w29769;
w29772 <= not w29770 and not w29771;
w29773 <= w5431 and w22250;
w29774 <= w4870 and w22255;
w29775 <= w5342 and w22247;
w29776 <= not w29774 and not w29775;
w29777 <= not w29773 and w29776;
w29778 <= w4873 and w25229;
w29779 <= w29777 and not w29778;
w29780 <= a(20) and not w29779;
w29781 <= a(20) and not w29780;
w29782 <= not w29779 and not w29780;
w29783 <= not w29781 and not w29782;
w29784 <= w29772 and not w29783;
w29785 <= w29772 and not w29784;
w29786 <= not w29783 and not w29784;
w29787 <= not w29785 and not w29786;
w29788 <= not w29574 and not w29587;
w29789 <= w29787 and w29788;
w29790 <= not w29787 and not w29788;
w29791 <= not w29789 and not w29790;
w29792 <= not w29593 and not w29606;
w29793 <= w6168 and w26001;
w29794 <= w5598 and w22244;
w29795 <= w5874 and w25998;
w29796 <= not w29794 and not w29795;
w29797 <= not w29793 and w29796;
w29798 <= w5601 and not w26559;
w29799 <= w29797 and not w29798;
w29800 <= a(17) and not w29799;
w29801 <= a(17) and not w29800;
w29802 <= not w29799 and not w29800;
w29803 <= not w29801 and not w29802;
w29804 <= not w29792 and not w29803;
w29805 <= not w29792 and not w29804;
w29806 <= not w29803 and not w29804;
w29807 <= not w29805 and not w29806;
w29808 <= not w29791 and w29807;
w29809 <= w29791 and not w29807;
w29810 <= not w29808 and not w29809;
w29811 <= w7036 and w27108;
w29812 <= w6337 and w25995;
w29813 <= w6886 and w26825;
w29814 <= not w29812 and not w29813;
w29815 <= not w29811 and w29814;
w29816 <= w6332 and w27120;
w29817 <= w29815 and not w29816;
w29818 <= a(14) and not w29817;
w29819 <= a(14) and not w29818;
w29820 <= not w29817 and not w29818;
w29821 <= not w29819 and not w29820;
w29822 <= w29810 and not w29821;
w29823 <= w29810 and not w29822;
w29824 <= not w29821 and not w29822;
w29825 <= not w29823 and not w29824;
w29826 <= not w29612 and not w29625;
w29827 <= w29825 and w29826;
w29828 <= not w29825 and not w29826;
w29829 <= not w29827 and not w29828;
w29830 <= not w29631 and not w29644;
w29831 <= w7918 and w27899;
w29832 <= w7226 and w27377;
w29833 <= w7567 and w27633;
w29834 <= not w29832 and not w29833;
w29835 <= not w29831 and w29834;
w29836 <= w7229 and w27911;
w29837 <= w29835 and not w29836;
w29838 <= a(11) and not w29837;
w29839 <= a(11) and not w29838;
w29840 <= not w29837 and not w29838;
w29841 <= not w29839 and not w29840;
w29842 <= not w29830 and not w29841;
w29843 <= not w29830 and not w29842;
w29844 <= not w29841 and not w29842;
w29845 <= not w29843 and not w29844;
w29846 <= not w29829 and w29845;
w29847 <= w29829 and not w29845;
w29848 <= not w29846 and not w29847;
w29849 <= not w29677 and w29848;
w29850 <= w29677 and not w29848;
w29851 <= not w29849 and not w29850;
w29852 <= not w29676 and w29851;
w29853 <= w29676 and not w29851;
w29854 <= not w29852 and not w29853;
w29855 <= not w29673 and not w29854;
w29856 <= w29673 and w29854;
w29857 <= not w29855 and not w29856;
w29858 <= not w29727 and not w29733;
w29859 <= w10 and not w23594;
w29860 <= w2955 and w22282;
w29861 <= w2958 and w22288;
w29862 <= w2963 and w22285;
w29863 <= not w29861 and not w29862;
w29864 <= not w29860 and w29863;
w29865 <= not w29859 and w29864;
w29866 <= not w29704 and not w29706;
w29867 <= w897 and w1425;
w29868 <= w15789 and w29867;
w29869 <= w14342 and w29868;
w29870 <= w4702 and w29869;
w29871 <= w4721 and w29870;
w29872 <= w1654 and w29871;
w29873 <= w3494 and w29872;
w29874 <= w2570 and w29873;
w29875 <= not w177 and w29874;
w29876 <= not w85 and w29875;
w29877 <= not w292 and w29876;
w29878 <= not w221 and w29877;
w29879 <= not w915 and w29878;
w29880 <= not w945 and w29879;
w29881 <= not w205 and w29880;
w29882 <= not w29866 and w29881;
w29883 <= w29866 and not w29881;
w29884 <= not w29882 and not w29883;
w29885 <= not w29865 and w29884;
w29886 <= not w29865 and not w29885;
w29887 <= w29884 and not w29885;
w29888 <= not w29886 and not w29887;
w29889 <= not w29709 and not w29712;
w29890 <= w29888 and w29889;
w29891 <= not w29888 and not w29889;
w29892 <= not w29890 and not w29891;
w29893 <= w3392 and w22273;
w29894 <= w3477 and w22279;
w29895 <= w3541 and w22276;
w29896 <= not w29894 and not w29895;
w29897 <= not w29893 and w29896;
w29898 <= not w3303 and w29897;
w29899 <= w24123 and w29897;
w29900 <= not w29898 and not w29899;
w29901 <= a(29) and not w29900;
w29902 <= not a(29) and w29900;
w29903 <= not w29901 and not w29902;
w29904 <= w29892 and not w29903;
w29905 <= not w29892 and w29903;
w29906 <= not w29904 and not w29905;
w29907 <= not w29858 and w29906;
w29908 <= w29858 and not w29906;
w29909 <= not w29907 and not w29908;
w29910 <= w3819 and w22264;
w29911 <= w3902 and w22270;
w29912 <= w3981 and w22267;
w29913 <= not w29911 and not w29912;
w29914 <= not w29910 and w29913;
w29915 <= w3985 and not w24568;
w29916 <= w29914 and not w29915;
w29917 <= a(26) and not w29916;
w29918 <= a(26) and not w29917;
w29919 <= not w29916 and not w29917;
w29920 <= not w29918 and not w29919;
w29921 <= w29909 and not w29920;
w29922 <= w29909 and not w29921;
w29923 <= not w29920 and not w29921;
w29924 <= not w29922 and not w29923;
w29925 <= not w29746 and not w29752;
w29926 <= w29924 and w29925;
w29927 <= not w29924 and not w29925;
w29928 <= not w29926 and not w29927;
w29929 <= w4629 and w22255;
w29930 <= w4468 and w22261;
w29931 <= w4539 and w22258;
w29932 <= not w29930 and not w29931;
w29933 <= not w29929 and w29932;
w29934 <= w4471 and not w25205;
w29935 <= w29933 and not w29934;
w29936 <= a(23) and not w29935;
w29937 <= a(23) and not w29936;
w29938 <= not w29935 and not w29936;
w29939 <= not w29937 and not w29938;
w29940 <= w29928 and not w29939;
w29941 <= w29928 and not w29940;
w29942 <= not w29939 and not w29940;
w29943 <= not w29941 and not w29942;
w29944 <= not w29765 and not w29771;
w29945 <= w29943 and w29944;
w29946 <= not w29943 and not w29944;
w29947 <= not w29945 and not w29946;
w29948 <= w5431 and w22244;
w29949 <= w4870 and w22247;
w29950 <= w5342 and w22250;
w29951 <= not w29949 and not w29950;
w29952 <= not w29948 and w29951;
w29953 <= w4873 and not w22464;
w29954 <= w29952 and not w29953;
w29955 <= a(20) and not w29954;
w29956 <= a(20) and not w29955;
w29957 <= not w29954 and not w29955;
w29958 <= not w29956 and not w29957;
w29959 <= w29947 and not w29958;
w29960 <= w29947 and not w29959;
w29961 <= not w29958 and not w29959;
w29962 <= not w29960 and not w29961;
w29963 <= not w29784 and not w29790;
w29964 <= w29962 and w29963;
w29965 <= not w29962 and not w29963;
w29966 <= not w29964 and not w29965;
w29967 <= w6168 and w25995;
w29968 <= w5598 and w25998;
w29969 <= w5874 and w26001;
w29970 <= not w29968 and not w29969;
w29971 <= not w29967 and w29970;
w29972 <= w5601 and not w26023;
w29973 <= w29971 and not w29972;
w29974 <= a(17) and not w29973;
w29975 <= a(17) and not w29974;
w29976 <= not w29973 and not w29974;
w29977 <= not w29975 and not w29976;
w29978 <= w29966 and not w29977;
w29979 <= w29966 and not w29978;
w29980 <= not w29977 and not w29978;
w29981 <= not w29979 and not w29980;
w29982 <= not w29804 and not w29809;
w29983 <= not w29981 and not w29982;
w29984 <= not w29981 and not w29983;
w29985 <= not w29982 and not w29983;
w29986 <= not w29984 and not w29985;
w29987 <= w7036 and w27377;
w29988 <= w6337 and w26825;
w29989 <= w6886 and w27108;
w29990 <= not w29988 and not w29989;
w29991 <= not w29987 and w29990;
w29992 <= w6332 and w27390;
w29993 <= w29991 and not w29992;
w29994 <= a(14) and not w29993;
w29995 <= a(14) and not w29994;
w29996 <= not w29993 and not w29994;
w29997 <= not w29995 and not w29996;
w29998 <= not w29986 and not w29997;
w29999 <= not w29986 and not w29998;
w30000 <= not w29997 and not w29998;
w30001 <= not w29999 and not w30000;
w30002 <= not w29822 and not w29828;
w30003 <= w30001 and w30002;
w30004 <= not w30001 and not w30002;
w30005 <= not w30003 and not w30004;
w30006 <= w7918 and not w28143;
w30007 <= w7226 and w27633;
w30008 <= w7567 and w27899;
w30009 <= not w30007 and not w30008;
w30010 <= not w30006 and w30009;
w30011 <= w7229 and not w28158;
w30012 <= w30010 and not w30011;
w30013 <= a(11) and not w30012;
w30014 <= a(11) and not w30013;
w30015 <= not w30012 and not w30013;
w30016 <= not w30014 and not w30015;
w30017 <= w30005 and not w30016;
w30018 <= w30005 and not w30017;
w30019 <= not w30016 and not w30017;
w30020 <= not w30018 and not w30019;
w30021 <= not w29842 and not w29847;
w30022 <= not w30020 and not w30021;
w30023 <= not w30020 and not w30022;
w30024 <= not w30021 and not w30022;
w30025 <= not w30023 and not w30024;
w30026 <= not w29849 and not w29852;
w30027 <= w30025 and w30026;
w30028 <= not w30025 and not w30026;
w30029 <= not w30027 and not w30028;
w30030 <= w29856 and not w30029;
w30031 <= not w29856 and w30029;
w30032 <= not w30030 and not w30031;
w30033 <= not w29891 and not w29904;
w30034 <= not w29882 and not w29885;
w30035 <= w2640 and w2746;
w30036 <= w1942 and w30035;
w30037 <= w947 and w30036;
w30038 <= w812 and w30037;
w30039 <= w13703 and w30038;
w30040 <= w15247 and w30039;
w30041 <= w5221 and w30040;
w30042 <= w2586 and w30041;
w30043 <= w226 and w30042;
w30044 <= w1265 and w30043;
w30045 <= w29272 and w30044;
w30046 <= w666 and w30045;
w30047 <= w1182 and w30046;
w30048 <= not w361 and w30047;
w30049 <= not w227 and w30048;
w30050 <= not w37 and w30049;
w30051 <= not w357 and w30050;
w30052 <= not w466 and w30051;
w30053 <= not w29881 and w30052;
w30054 <= w29881 and not w30052;
w30055 <= not w30034 and not w30054;
w30056 <= not w30053 and w30055;
w30057 <= not w30034 and not w30056;
w30058 <= not w30054 and not w30056;
w30059 <= not w30053 and w30058;
w30060 <= not w30057 and not w30059;
w30061 <= w10 and not w23577;
w30062 <= w2955 and w22279;
w30063 <= w2958 and w22285;
w30064 <= w2963 and w22282;
w30065 <= not w30063 and not w30064;
w30066 <= not w30062 and w30065;
w30067 <= not w30061 and w30066;
w30068 <= not w30060 and not w30067;
w30069 <= not w30060 and not w30068;
w30070 <= not w30067 and not w30068;
w30071 <= not w30069 and not w30070;
w30072 <= w3392 and w22270;
w30073 <= w3477 and w22276;
w30074 <= w3541 and w22273;
w30075 <= not w30073 and not w30074;
w30076 <= not w30072 and w30075;
w30077 <= not w3303 and w30076;
w30078 <= w24102 and w30076;
w30079 <= not w30077 and not w30078;
w30080 <= a(29) and not w30079;
w30081 <= not a(29) and w30079;
w30082 <= not w30080 and not w30081;
w30083 <= not w30071 and not w30082;
w30084 <= w30071 and w30082;
w30085 <= not w30083 and not w30084;
w30086 <= not w30033 and w30085;
w30087 <= w30033 and not w30085;
w30088 <= not w30086 and not w30087;
w30089 <= w3819 and w22261;
w30090 <= w3902 and w22267;
w30091 <= w3981 and w22264;
w30092 <= not w30090 and not w30091;
w30093 <= not w30089 and w30092;
w30094 <= w3985 and not w24551;
w30095 <= w30093 and not w30094;
w30096 <= a(26) and not w30095;
w30097 <= a(26) and not w30096;
w30098 <= not w30095 and not w30096;
w30099 <= not w30097 and not w30098;
w30100 <= w30088 and not w30099;
w30101 <= w30088 and not w30100;
w30102 <= not w30099 and not w30100;
w30103 <= not w30101 and not w30102;
w30104 <= not w29907 and not w29921;
w30105 <= w30103 and w30104;
w30106 <= not w30103 and not w30104;
w30107 <= not w30105 and not w30106;
w30108 <= w4629 and w22247;
w30109 <= w4468 and w22258;
w30110 <= w4539 and w22255;
w30111 <= not w30109 and not w30110;
w30112 <= not w30108 and w30111;
w30113 <= w4471 and not w25250;
w30114 <= w30112 and not w30113;
w30115 <= a(23) and not w30114;
w30116 <= a(23) and not w30115;
w30117 <= not w30114 and not w30115;
w30118 <= not w30116 and not w30117;
w30119 <= w30107 and not w30118;
w30120 <= w30107 and not w30119;
w30121 <= not w30118 and not w30119;
w30122 <= not w30120 and not w30121;
w30123 <= not w29927 and not w29940;
w30124 <= w30122 and w30123;
w30125 <= not w30122 and not w30123;
w30126 <= not w30124 and not w30125;
w30127 <= w5431 and w25998;
w30128 <= w4870 and w22250;
w30129 <= w5342 and w22244;
w30130 <= not w30128 and not w30129;
w30131 <= not w30127 and w30130;
w30132 <= w4873 and not w26539;
w30133 <= w30131 and not w30132;
w30134 <= a(20) and not w30133;
w30135 <= a(20) and not w30134;
w30136 <= not w30133 and not w30134;
w30137 <= not w30135 and not w30136;
w30138 <= w30126 and not w30137;
w30139 <= w30126 and not w30138;
w30140 <= not w30137 and not w30138;
w30141 <= not w30139 and not w30140;
w30142 <= not w29946 and not w29959;
w30143 <= w30141 and w30142;
w30144 <= not w30141 and not w30142;
w30145 <= not w30143 and not w30144;
w30146 <= w6168 and w26825;
w30147 <= w5598 and w26001;
w30148 <= w5874 and w25995;
w30149 <= not w30147 and not w30148;
w30150 <= not w30146 and w30149;
w30151 <= w5601 and not w26839;
w30152 <= w30150 and not w30151;
w30153 <= a(17) and not w30152;
w30154 <= a(17) and not w30153;
w30155 <= not w30152 and not w30153;
w30156 <= not w30154 and not w30155;
w30157 <= w30145 and not w30156;
w30158 <= w30145 and not w30157;
w30159 <= not w30156 and not w30157;
w30160 <= not w30158 and not w30159;
w30161 <= not w29965 and not w29978;
w30162 <= w30160 and w30161;
w30163 <= not w30160 and not w30161;
w30164 <= not w30162 and not w30163;
w30165 <= w7036 and w27633;
w30166 <= w6337 and w27108;
w30167 <= w6886 and w27377;
w30168 <= not w30166 and not w30167;
w30169 <= not w30165 and w30168;
w30170 <= w6332 and not w27648;
w30171 <= w30169 and not w30170;
w30172 <= a(14) and not w30171;
w30173 <= a(14) and not w30172;
w30174 <= not w30171 and not w30172;
w30175 <= not w30173 and not w30174;
w30176 <= w30164 and not w30175;
w30177 <= w30164 and not w30176;
w30178 <= not w30175 and not w30176;
w30179 <= not w30177 and not w30178;
w30180 <= not w29983 and not w29998;
w30181 <= not w14359 and not w28143;
w30182 <= w7226 and w27899;
w30183 <= not w30181 and not w30182;
w30184 <= not w7229 and w30183;
w30185 <= w28156 and w30183;
w30186 <= not w30184 and not w30185;
w30187 <= a(11) and not w30186;
w30188 <= not a(11) and w30186;
w30189 <= not w30187 and not w30188;
w30190 <= not w30180 and not w30189;
w30191 <= w30180 and w30189;
w30192 <= not w30190 and not w30191;
w30193 <= not w30179 and w30192;
w30194 <= not w30179 and not w30193;
w30195 <= w30192 and not w30193;
w30196 <= not w30194 and not w30195;
w30197 <= not w30004 and not w30017;
w30198 <= w30196 and w30197;
w30199 <= not w30196 and not w30197;
w30200 <= not w30198 and not w30199;
w30201 <= not w30022 and not w30028;
w30202 <= not w30200 and w30201;
w30203 <= w30200 and not w30201;
w30204 <= not w30202 and not w30203;
w30205 <= w29856 and w30029;
w30206 <= w30204 and w30205;
w30207 <= not w30204 and not w30205;
w30208 <= not w30206 and not w30207;
w30209 <= not w30199 and not w30203;
w30210 <= not w30190 and not w30193;
w30211 <= not w30068 and not w30083;
w30212 <= w10 and w24077;
w30213 <= w2955 and w22276;
w30214 <= w2958 and w22282;
w30215 <= w2963 and w22279;
w30216 <= not w30214 and not w30215;
w30217 <= not w30213 and w30216;
w30218 <= not w30212 and w30217;
w30219 <= not w14361 and not w28143;
w30220 <= a(11) and not w30219;
w30221 <= not a(11) and w30219;
w30222 <= not w30220 and not w30221;
w30223 <= w610 and w2109;
w30224 <= w4973 and w30223;
w30225 <= w2743 and w30224;
w30226 <= w4954 and w30225;
w30227 <= w1342 and w30226;
w30228 <= w3445 and w30227;
w30229 <= w176 and w30228;
w30230 <= w1370 and w30229;
w30231 <= w1511 and w30230;
w30232 <= w1187 and w30231;
w30233 <= w3821 and w30232;
w30234 <= w525 and w30233;
w30235 <= not w177 and w30234;
w30236 <= not w370 and w30235;
w30237 <= not w467 and w30236;
w30238 <= not w298 and w30237;
w30239 <= w29881 and w30238;
w30240 <= not w29881 and not w30238;
w30241 <= not w30239 and not w30240;
w30242 <= w30222 and w30241;
w30243 <= not w30222 and not w30241;
w30244 <= not w30242 and not w30243;
w30245 <= not w30218 and w30244;
w30246 <= w30244 and not w30245;
w30247 <= not w30218 and not w30245;
w30248 <= not w30246 and not w30247;
w30249 <= not w30058 and not w30248;
w30250 <= not w30248 and not w30249;
w30251 <= not w30058 and not w30249;
w30252 <= not w30250 and not w30251;
w30253 <= not w30211 and not w30252;
w30254 <= not w30211 and not w30253;
w30255 <= not w30252 and not w30253;
w30256 <= not w30254 and not w30255;
w30257 <= w3392 and w22267;
w30258 <= w3477 and w22273;
w30259 <= w3541 and w22270;
w30260 <= not w30258 and not w30259;
w30261 <= not w30257 and w30260;
w30262 <= w3303 and w22477;
w30263 <= w30261 and not w30262;
w30264 <= a(29) and not w30263;
w30265 <= a(29) and not w30264;
w30266 <= not w30263 and not w30264;
w30267 <= not w30265 and not w30266;
w30268 <= not w30256 and not w30267;
w30269 <= not w30256 and not w30268;
w30270 <= not w30267 and not w30268;
w30271 <= not w30269 and not w30270;
w30272 <= w3819 and w22258;
w30273 <= w3902 and w22264;
w30274 <= w3981 and w22261;
w30275 <= not w30273 and not w30274;
w30276 <= not w30272 and w30275;
w30277 <= w3985 and w24534;
w30278 <= w30276 and not w30277;
w30279 <= a(26) and not w30278;
w30280 <= a(26) and not w30279;
w30281 <= not w30278 and not w30279;
w30282 <= not w30280 and not w30281;
w30283 <= not w30271 and not w30282;
w30284 <= not w30271 and not w30283;
w30285 <= not w30282 and not w30283;
w30286 <= not w30284 and not w30285;
w30287 <= not w30086 and not w30100;
w30288 <= w30286 and w30287;
w30289 <= not w30286 and not w30287;
w30290 <= not w30288 and not w30289;
w30291 <= w4629 and w22250;
w30292 <= w4468 and w22255;
w30293 <= w4539 and w22247;
w30294 <= not w30292 and not w30293;
w30295 <= not w30291 and w30294;
w30296 <= w4471 and w25229;
w30297 <= w30295 and not w30296;
w30298 <= a(23) and not w30297;
w30299 <= a(23) and not w30298;
w30300 <= not w30297 and not w30298;
w30301 <= not w30299 and not w30300;
w30302 <= w30290 and not w30301;
w30303 <= w30290 and not w30302;
w30304 <= not w30301 and not w30302;
w30305 <= not w30303 and not w30304;
w30306 <= not w30106 and not w30119;
w30307 <= w30305 and w30306;
w30308 <= not w30305 and not w30306;
w30309 <= not w30307 and not w30308;
w30310 <= not w30125 and not w30138;
w30311 <= w5431 and w26001;
w30312 <= w4870 and w22244;
w30313 <= w5342 and w25998;
w30314 <= not w30312 and not w30313;
w30315 <= not w30311 and w30314;
w30316 <= w4873 and not w26559;
w30317 <= w30315 and not w30316;
w30318 <= a(20) and not w30317;
w30319 <= a(20) and not w30318;
w30320 <= not w30317 and not w30318;
w30321 <= not w30319 and not w30320;
w30322 <= not w30310 and not w30321;
w30323 <= not w30310 and not w30322;
w30324 <= not w30321 and not w30322;
w30325 <= not w30323 and not w30324;
w30326 <= not w30309 and w30325;
w30327 <= w30309 and not w30325;
w30328 <= not w30326 and not w30327;
w30329 <= w6168 and w27108;
w30330 <= w5598 and w25995;
w30331 <= w5874 and w26825;
w30332 <= not w30330 and not w30331;
w30333 <= not w30329 and w30332;
w30334 <= w5601 and w27120;
w30335 <= w30333 and not w30334;
w30336 <= a(17) and not w30335;
w30337 <= a(17) and not w30336;
w30338 <= not w30335 and not w30336;
w30339 <= not w30337 and not w30338;
w30340 <= w30328 and not w30339;
w30341 <= w30328 and not w30340;
w30342 <= not w30339 and not w30340;
w30343 <= not w30341 and not w30342;
w30344 <= not w30144 and not w30157;
w30345 <= w30343 and w30344;
w30346 <= not w30343 and not w30344;
w30347 <= not w30345 and not w30346;
w30348 <= not w30163 and not w30176;
w30349 <= w7036 and w27899;
w30350 <= w6337 and w27377;
w30351 <= w6886 and w27633;
w30352 <= not w30350 and not w30351;
w30353 <= not w30349 and w30352;
w30354 <= w6332 and w27911;
w30355 <= w30353 and not w30354;
w30356 <= a(14) and not w30355;
w30357 <= a(14) and not w30356;
w30358 <= not w30355 and not w30356;
w30359 <= not w30357 and not w30358;
w30360 <= not w30348 and not w30359;
w30361 <= not w30348 and not w30360;
w30362 <= not w30359 and not w30360;
w30363 <= not w30361 and not w30362;
w30364 <= not w30347 and w30363;
w30365 <= w30347 and not w30363;
w30366 <= not w30364 and not w30365;
w30367 <= not w30210 and w30366;
w30368 <= w30210 and not w30366;
w30369 <= not w30367 and not w30368;
w30370 <= not w30209 and w30369;
w30371 <= w30209 and not w30369;
w30372 <= not w30370 and not w30371;
w30373 <= not w30206 and not w30372;
w30374 <= w30206 and w30372;
w30375 <= not w30373 and not w30374;
w30376 <= not w30253 and not w30268;
w30377 <= w10 and not w24123;
w30378 <= w2955 and w22273;
w30379 <= w2958 and w22279;
w30380 <= w2963 and w22276;
w30381 <= not w30379 and not w30380;
w30382 <= not w30378 and w30381;
w30383 <= not w30377 and w30382;
w30384 <= not w30240 and not w30242;
w30385 <= w1434 and w1994;
w30386 <= w713 and w30385;
w30387 <= w3063 and w30386;
w30388 <= w12912 and w30387;
w30389 <= w27724 and w30388;
w30390 <= w13393 and w30389;
w30391 <= w15259 and w30390;
w30392 <= w28229 and w30391;
w30393 <= w1315 and w30392;
w30394 <= w745 and w30393;
w30395 <= not w404 and w30394;
w30396 <= not w681 and w30395;
w30397 <= not w1037 and w30396;
w30398 <= not w331 and w30397;
w30399 <= not w405 and w30398;
w30400 <= not w30384 and w30399;
w30401 <= w30384 and not w30399;
w30402 <= not w30400 and not w30401;
w30403 <= not w30383 and w30402;
w30404 <= not w30383 and not w30403;
w30405 <= w30402 and not w30403;
w30406 <= not w30404 and not w30405;
w30407 <= not w30245 and not w30249;
w30408 <= w30406 and w30407;
w30409 <= not w30406 and not w30407;
w30410 <= not w30408 and not w30409;
w30411 <= w3392 and w22264;
w30412 <= w3477 and w22270;
w30413 <= w3541 and w22267;
w30414 <= not w30412 and not w30413;
w30415 <= not w30411 and w30414;
w30416 <= not w3303 and w30415;
w30417 <= w24568 and w30415;
w30418 <= not w30416 and not w30417;
w30419 <= a(29) and not w30418;
w30420 <= not a(29) and w30418;
w30421 <= not w30419 and not w30420;
w30422 <= w30410 and not w30421;
w30423 <= not w30410 and w30421;
w30424 <= not w30422 and not w30423;
w30425 <= not w30376 and w30424;
w30426 <= w30376 and not w30424;
w30427 <= not w30425 and not w30426;
w30428 <= w3819 and w22255;
w30429 <= w3902 and w22261;
w30430 <= w3981 and w22258;
w30431 <= not w30429 and not w30430;
w30432 <= not w30428 and w30431;
w30433 <= w3985 and not w25205;
w30434 <= w30432 and not w30433;
w30435 <= a(26) and not w30434;
w30436 <= a(26) and not w30435;
w30437 <= not w30434 and not w30435;
w30438 <= not w30436 and not w30437;
w30439 <= w30427 and not w30438;
w30440 <= w30427 and not w30439;
w30441 <= not w30438 and not w30439;
w30442 <= not w30440 and not w30441;
w30443 <= not w30283 and not w30289;
w30444 <= w30442 and w30443;
w30445 <= not w30442 and not w30443;
w30446 <= not w30444 and not w30445;
w30447 <= w4629 and w22244;
w30448 <= w4468 and w22247;
w30449 <= w4539 and w22250;
w30450 <= not w30448 and not w30449;
w30451 <= not w30447 and w30450;
w30452 <= w4471 and not w22464;
w30453 <= w30451 and not w30452;
w30454 <= a(23) and not w30453;
w30455 <= a(23) and not w30454;
w30456 <= not w30453 and not w30454;
w30457 <= not w30455 and not w30456;
w30458 <= w30446 and not w30457;
w30459 <= w30446 and not w30458;
w30460 <= not w30457 and not w30458;
w30461 <= not w30459 and not w30460;
w30462 <= not w30302 and not w30308;
w30463 <= w30461 and w30462;
w30464 <= not w30461 and not w30462;
w30465 <= not w30463 and not w30464;
w30466 <= w5431 and w25995;
w30467 <= w4870 and w25998;
w30468 <= w5342 and w26001;
w30469 <= not w30467 and not w30468;
w30470 <= not w30466 and w30469;
w30471 <= w4873 and not w26023;
w30472 <= w30470 and not w30471;
w30473 <= a(20) and not w30472;
w30474 <= a(20) and not w30473;
w30475 <= not w30472 and not w30473;
w30476 <= not w30474 and not w30475;
w30477 <= w30465 and not w30476;
w30478 <= w30465 and not w30477;
w30479 <= not w30476 and not w30477;
w30480 <= not w30478 and not w30479;
w30481 <= not w30322 and not w30327;
w30482 <= not w30480 and not w30481;
w30483 <= not w30480 and not w30482;
w30484 <= not w30481 and not w30482;
w30485 <= not w30483 and not w30484;
w30486 <= w6168 and w27377;
w30487 <= w5598 and w26825;
w30488 <= w5874 and w27108;
w30489 <= not w30487 and not w30488;
w30490 <= not w30486 and w30489;
w30491 <= w5601 and w27390;
w30492 <= w30490 and not w30491;
w30493 <= a(17) and not w30492;
w30494 <= a(17) and not w30493;
w30495 <= not w30492 and not w30493;
w30496 <= not w30494 and not w30495;
w30497 <= not w30485 and not w30496;
w30498 <= not w30485 and not w30497;
w30499 <= not w30496 and not w30497;
w30500 <= not w30498 and not w30499;
w30501 <= not w30340 and not w30346;
w30502 <= w30500 and w30501;
w30503 <= not w30500 and not w30501;
w30504 <= not w30502 and not w30503;
w30505 <= w7036 and not w28143;
w30506 <= w6337 and w27633;
w30507 <= w6886 and w27899;
w30508 <= not w30506 and not w30507;
w30509 <= not w30505 and w30508;
w30510 <= w6332 and not w28158;
w30511 <= w30509 and not w30510;
w30512 <= a(14) and not w30511;
w30513 <= a(14) and not w30512;
w30514 <= not w30511 and not w30512;
w30515 <= not w30513 and not w30514;
w30516 <= w30504 and not w30515;
w30517 <= w30504 and not w30516;
w30518 <= not w30515 and not w30516;
w30519 <= not w30517 and not w30518;
w30520 <= not w30360 and not w30365;
w30521 <= not w30519 and not w30520;
w30522 <= not w30519 and not w30521;
w30523 <= not w30520 and not w30521;
w30524 <= not w30522 and not w30523;
w30525 <= not w30367 and not w30370;
w30526 <= w30524 and w30525;
w30527 <= not w30524 and not w30525;
w30528 <= not w30526 and not w30527;
w30529 <= not w30374 and w30528;
w30530 <= w30374 and not w30528;
w30531 <= not w30529 and not w30530;
w30532 <= w30374 and w30528;
w30533 <= w10 and not w24102;
w30534 <= w2955 and w22270;
w30535 <= w2958 and w22276;
w30536 <= w2963 and w22273;
w30537 <= not w30535 and not w30536;
w30538 <= not w30534 and w30537;
w30539 <= not w30533 and w30538;
w30540 <= w629 and w2111;
w30541 <= w6019 and w30540;
w30542 <= w3043 and w30541;
w30543 <= w12645 and w30542;
w30544 <= w13058 and w30543;
w30545 <= w3321 and w30544;
w30546 <= w2435 and w30545;
w30547 <= w5144 and w30546;
w30548 <= w2674 and w30547;
w30549 <= not w493 and w30548;
w30550 <= not w1037 and w30549;
w30551 <= not w90 and w30550;
w30552 <= not w183 and w30551;
w30553 <= not w292 and w30552;
w30554 <= not w140 and w30553;
w30555 <= not w371 and w30554;
w30556 <= not w16 and w30555;
w30557 <= not w30399 and w30556;
w30558 <= w30399 and not w30556;
w30559 <= not w30539 and not w30558;
w30560 <= not w30557 and w30559;
w30561 <= not w30539 and not w30560;
w30562 <= not w30558 and not w30560;
w30563 <= not w30557 and w30562;
w30564 <= not w30561 and not w30563;
w30565 <= not w30400 and not w30403;
w30566 <= w30564 and w30565;
w30567 <= not w30564 and not w30565;
w30568 <= not w30566 and not w30567;
w30569 <= not w30409 and not w30422;
w30570 <= not w30568 and w30569;
w30571 <= w30568 and not w30569;
w30572 <= not w30570 and not w30571;
w30573 <= w3392 and w22261;
w30574 <= w3477 and w22267;
w30575 <= w3541 and w22264;
w30576 <= not w30574 and not w30575;
w30577 <= not w30573 and w30576;
w30578 <= w3303 and not w24551;
w30579 <= w30577 and not w30578;
w30580 <= a(29) and not w30579;
w30581 <= a(29) and not w30580;
w30582 <= not w30579 and not w30580;
w30583 <= not w30581 and not w30582;
w30584 <= w30572 and not w30583;
w30585 <= w30572 and not w30584;
w30586 <= not w30583 and not w30584;
w30587 <= not w30585 and not w30586;
w30588 <= w3819 and w22247;
w30589 <= w3902 and w22258;
w30590 <= w3981 and w22255;
w30591 <= not w30589 and not w30590;
w30592 <= not w30588 and w30591;
w30593 <= w3985 and not w25250;
w30594 <= w30592 and not w30593;
w30595 <= a(26) and not w30594;
w30596 <= a(26) and not w30595;
w30597 <= not w30594 and not w30595;
w30598 <= not w30596 and not w30597;
w30599 <= not w30587 and not w30598;
w30600 <= not w30587 and not w30599;
w30601 <= not w30598 and not w30599;
w30602 <= not w30600 and not w30601;
w30603 <= not w30425 and not w30439;
w30604 <= w30602 and w30603;
w30605 <= not w30602 and not w30603;
w30606 <= not w30604 and not w30605;
w30607 <= w4629 and w25998;
w30608 <= w4468 and w22250;
w30609 <= w4539 and w22244;
w30610 <= not w30608 and not w30609;
w30611 <= not w30607 and w30610;
w30612 <= w4471 and not w26539;
w30613 <= w30611 and not w30612;
w30614 <= a(23) and not w30613;
w30615 <= a(23) and not w30614;
w30616 <= not w30613 and not w30614;
w30617 <= not w30615 and not w30616;
w30618 <= w30606 and not w30617;
w30619 <= w30606 and not w30618;
w30620 <= not w30617 and not w30618;
w30621 <= not w30619 and not w30620;
w30622 <= not w30445 and not w30458;
w30623 <= w30621 and w30622;
w30624 <= not w30621 and not w30622;
w30625 <= not w30623 and not w30624;
w30626 <= w5431 and w26825;
w30627 <= w4870 and w26001;
w30628 <= w5342 and w25995;
w30629 <= not w30627 and not w30628;
w30630 <= not w30626 and w30629;
w30631 <= w4873 and not w26839;
w30632 <= w30630 and not w30631;
w30633 <= a(20) and not w30632;
w30634 <= a(20) and not w30633;
w30635 <= not w30632 and not w30633;
w30636 <= not w30634 and not w30635;
w30637 <= w30625 and not w30636;
w30638 <= w30625 and not w30637;
w30639 <= not w30636 and not w30637;
w30640 <= not w30638 and not w30639;
w30641 <= not w30464 and not w30477;
w30642 <= w30640 and w30641;
w30643 <= not w30640 and not w30641;
w30644 <= not w30642 and not w30643;
w30645 <= w6168 and w27633;
w30646 <= w5598 and w27108;
w30647 <= w5874 and w27377;
w30648 <= not w30646 and not w30647;
w30649 <= not w30645 and w30648;
w30650 <= w5601 and not w27648;
w30651 <= w30649 and not w30650;
w30652 <= a(17) and not w30651;
w30653 <= a(17) and not w30652;
w30654 <= not w30651 and not w30652;
w30655 <= not w30653 and not w30654;
w30656 <= w30644 and not w30655;
w30657 <= w30644 and not w30656;
w30658 <= not w30655 and not w30656;
w30659 <= not w30657 and not w30658;
w30660 <= not w30482 and not w30497;
w30661 <= not w13780 and not w28143;
w30662 <= w6337 and w27899;
w30663 <= not w30661 and not w30662;
w30664 <= not w6332 and w30663;
w30665 <= w28156 and w30663;
w30666 <= not w30664 and not w30665;
w30667 <= a(14) and not w30666;
w30668 <= not a(14) and w30666;
w30669 <= not w30667 and not w30668;
w30670 <= not w30660 and not w30669;
w30671 <= w30660 and w30669;
w30672 <= not w30670 and not w30671;
w30673 <= not w30659 and w30672;
w30674 <= not w30659 and not w30673;
w30675 <= w30672 and not w30673;
w30676 <= not w30674 and not w30675;
w30677 <= not w30503 and not w30516;
w30678 <= w30676 and w30677;
w30679 <= not w30676 and not w30677;
w30680 <= not w30678 and not w30679;
w30681 <= not w30521 and not w30527;
w30682 <= not w30680 and w30681;
w30683 <= w30680 and not w30681;
w30684 <= not w30682 and not w30683;
w30685 <= w30532 and w30684;
w30686 <= not w30532 and not w30684;
w30687 <= not w30685 and not w30686;
w30688 <= not w30679 and not w30683;
w30689 <= not w30670 and not w30673;
w30690 <= w10 and w22477;
w30691 <= w2955 and w22267;
w30692 <= w2958 and w22273;
w30693 <= w2963 and w22270;
w30694 <= not w30692 and not w30693;
w30695 <= not w30691 and w30694;
w30696 <= not w30690 and w30695;
w30697 <= not w13782 and not w28143;
w30698 <= a(14) and not w30697;
w30699 <= not a(14) and w30697;
w30700 <= not w30698 and not w30699;
w30701 <= w2472 and w2980;
w30702 <= w14417 and w30701;
w30703 <= w1829 and w30702;
w30704 <= w14137 and w30703;
w30705 <= w6649 and w30704;
w30706 <= w1226 and w30705;
w30707 <= w911 and w30706;
w30708 <= w1074 and w30707;
w30709 <= w2154 and w30708;
w30710 <= not w292 and w30709;
w30711 <= not w261 and w30710;
w30712 <= not w387 and w30711;
w30713 <= w30399 and w30712;
w30714 <= not w30399 and not w30712;
w30715 <= not w30713 and not w30714;
w30716 <= w30700 and w30715;
w30717 <= not w30700 and not w30715;
w30718 <= not w30716 and not w30717;
w30719 <= not w30562 and w30718;
w30720 <= w30562 and not w30718;
w30721 <= not w30719 and not w30720;
w30722 <= not w30696 and w30721;
w30723 <= w30721 and not w30722;
w30724 <= not w30696 and not w30722;
w30725 <= not w30723 and not w30724;
w30726 <= w3392 and w22258;
w30727 <= w3477 and w22264;
w30728 <= w3541 and w22261;
w30729 <= not w30727 and not w30728;
w30730 <= not w30726 and w30729;
w30731 <= w3303 and w24534;
w30732 <= w30730 and not w30731;
w30733 <= a(29) and not w30732;
w30734 <= a(29) and not w30733;
w30735 <= not w30732 and not w30733;
w30736 <= not w30734 and not w30735;
w30737 <= not w30725 and not w30736;
w30738 <= not w30725 and not w30737;
w30739 <= not w30736 and not w30737;
w30740 <= not w30738 and not w30739;
w30741 <= not w30567 and not w30571;
w30742 <= w30740 and w30741;
w30743 <= not w30740 and not w30741;
w30744 <= not w30742 and not w30743;
w30745 <= w3819 and w22250;
w30746 <= w3902 and w22255;
w30747 <= w3981 and w22247;
w30748 <= not w30746 and not w30747;
w30749 <= not w30745 and w30748;
w30750 <= w3985 and w25229;
w30751 <= w30749 and not w30750;
w30752 <= a(26) and not w30751;
w30753 <= a(26) and not w30752;
w30754 <= not w30751 and not w30752;
w30755 <= not w30753 and not w30754;
w30756 <= w30744 and not w30755;
w30757 <= w30744 and not w30756;
w30758 <= not w30755 and not w30756;
w30759 <= not w30757 and not w30758;
w30760 <= not w30584 and not w30599;
w30761 <= w30759 and w30760;
w30762 <= not w30759 and not w30760;
w30763 <= not w30761 and not w30762;
w30764 <= not w30605 and not w30618;
w30765 <= w4629 and w26001;
w30766 <= w4468 and w22244;
w30767 <= w4539 and w25998;
w30768 <= not w30766 and not w30767;
w30769 <= not w30765 and w30768;
w30770 <= w4471 and not w26559;
w30771 <= w30769 and not w30770;
w30772 <= a(23) and not w30771;
w30773 <= a(23) and not w30772;
w30774 <= not w30771 and not w30772;
w30775 <= not w30773 and not w30774;
w30776 <= not w30764 and not w30775;
w30777 <= not w30764 and not w30776;
w30778 <= not w30775 and not w30776;
w30779 <= not w30777 and not w30778;
w30780 <= not w30763 and w30779;
w30781 <= w30763 and not w30779;
w30782 <= not w30780 and not w30781;
w30783 <= w5431 and w27108;
w30784 <= w4870 and w25995;
w30785 <= w5342 and w26825;
w30786 <= not w30784 and not w30785;
w30787 <= not w30783 and w30786;
w30788 <= w4873 and w27120;
w30789 <= w30787 and not w30788;
w30790 <= a(20) and not w30789;
w30791 <= a(20) and not w30790;
w30792 <= not w30789 and not w30790;
w30793 <= not w30791 and not w30792;
w30794 <= w30782 and not w30793;
w30795 <= w30782 and not w30794;
w30796 <= not w30793 and not w30794;
w30797 <= not w30795 and not w30796;
w30798 <= not w30624 and not w30637;
w30799 <= w30797 and w30798;
w30800 <= not w30797 and not w30798;
w30801 <= not w30799 and not w30800;
w30802 <= not w30643 and not w30656;
w30803 <= w6168 and w27899;
w30804 <= w5598 and w27377;
w30805 <= w5874 and w27633;
w30806 <= not w30804 and not w30805;
w30807 <= not w30803 and w30806;
w30808 <= w5601 and w27911;
w30809 <= w30807 and not w30808;
w30810 <= a(17) and not w30809;
w30811 <= a(17) and not w30810;
w30812 <= not w30809 and not w30810;
w30813 <= not w30811 and not w30812;
w30814 <= not w30802 and not w30813;
w30815 <= not w30802 and not w30814;
w30816 <= not w30813 and not w30814;
w30817 <= not w30815 and not w30816;
w30818 <= not w30801 and w30817;
w30819 <= w30801 and not w30817;
w30820 <= not w30818 and not w30819;
w30821 <= not w30689 and w30820;
w30822 <= w30689 and not w30820;
w30823 <= not w30821 and not w30822;
w30824 <= not w30688 and w30823;
w30825 <= w30688 and not w30823;
w30826 <= not w30824 and not w30825;
w30827 <= not w30685 and not w30826;
w30828 <= w30685 and w30826;
w30829 <= not w30827 and not w30828;
w30830 <= not w30737 and not w30743;
w30831 <= w10 and not w24568;
w30832 <= w2955 and w22264;
w30833 <= w2958 and w22270;
w30834 <= w2963 and w22267;
w30835 <= not w30833 and not w30834;
w30836 <= not w30832 and w30835;
w30837 <= not w30831 and w30836;
w30838 <= not w30714 and not w30716;
w30839 <= w1304 and w3328;
w30840 <= w2296 and w30839;
w30841 <= w14460 and w30840;
w30842 <= w4969 and w30841;
w30843 <= w5708 and w30842;
w30844 <= w912 and w30843;
w30845 <= w426 and w30844;
w30846 <= w1118 and w30845;
w30847 <= w2281 and w30846;
w30848 <= w2632 and w30847;
w30849 <= w406 and w30848;
w30850 <= w1717 and w30849;
w30851 <= not w159 and w30850;
w30852 <= not w81 and w30851;
w30853 <= not w96 and w30852;
w30854 <= not w293 and w30853;
w30855 <= not w30838 and w30854;
w30856 <= w30838 and not w30854;
w30857 <= not w30855 and not w30856;
w30858 <= not w30837 and w30857;
w30859 <= not w30837 and not w30858;
w30860 <= w30857 and not w30858;
w30861 <= not w30859 and not w30860;
w30862 <= not w30719 and not w30722;
w30863 <= w30861 and w30862;
w30864 <= not w30861 and not w30862;
w30865 <= not w30863 and not w30864;
w30866 <= w3392 and w22255;
w30867 <= w3477 and w22261;
w30868 <= w3541 and w22258;
w30869 <= not w30867 and not w30868;
w30870 <= not w30866 and w30869;
w30871 <= not w3303 and w30870;
w30872 <= w25205 and w30870;
w30873 <= not w30871 and not w30872;
w30874 <= a(29) and not w30873;
w30875 <= not a(29) and w30873;
w30876 <= not w30874 and not w30875;
w30877 <= w30865 and not w30876;
w30878 <= not w30865 and w30876;
w30879 <= not w30877 and not w30878;
w30880 <= not w30830 and w30879;
w30881 <= w30830 and not w30879;
w30882 <= not w30880 and not w30881;
w30883 <= w3819 and w22244;
w30884 <= w3902 and w22247;
w30885 <= w3981 and w22250;
w30886 <= not w30884 and not w30885;
w30887 <= not w30883 and w30886;
w30888 <= w3985 and not w22464;
w30889 <= w30887 and not w30888;
w30890 <= a(26) and not w30889;
w30891 <= a(26) and not w30890;
w30892 <= not w30889 and not w30890;
w30893 <= not w30891 and not w30892;
w30894 <= w30882 and not w30893;
w30895 <= w30882 and not w30894;
w30896 <= not w30893 and not w30894;
w30897 <= not w30895 and not w30896;
w30898 <= not w30756 and not w30762;
w30899 <= w30897 and w30898;
w30900 <= not w30897 and not w30898;
w30901 <= not w30899 and not w30900;
w30902 <= w4629 and w25995;
w30903 <= w4468 and w25998;
w30904 <= w4539 and w26001;
w30905 <= not w30903 and not w30904;
w30906 <= not w30902 and w30905;
w30907 <= w4471 and not w26023;
w30908 <= w30906 and not w30907;
w30909 <= a(23) and not w30908;
w30910 <= a(23) and not w30909;
w30911 <= not w30908 and not w30909;
w30912 <= not w30910 and not w30911;
w30913 <= w30901 and not w30912;
w30914 <= w30901 and not w30913;
w30915 <= not w30912 and not w30913;
w30916 <= not w30914 and not w30915;
w30917 <= not w30776 and not w30781;
w30918 <= not w30916 and not w30917;
w30919 <= not w30916 and not w30918;
w30920 <= not w30917 and not w30918;
w30921 <= not w30919 and not w30920;
w30922 <= w5431 and w27377;
w30923 <= w4870 and w26825;
w30924 <= w5342 and w27108;
w30925 <= not w30923 and not w30924;
w30926 <= not w30922 and w30925;
w30927 <= w4873 and w27390;
w30928 <= w30926 and not w30927;
w30929 <= a(20) and not w30928;
w30930 <= a(20) and not w30929;
w30931 <= not w30928 and not w30929;
w30932 <= not w30930 and not w30931;
w30933 <= not w30921 and not w30932;
w30934 <= not w30921 and not w30933;
w30935 <= not w30932 and not w30933;
w30936 <= not w30934 and not w30935;
w30937 <= not w30794 and not w30800;
w30938 <= w30936 and w30937;
w30939 <= not w30936 and not w30937;
w30940 <= not w30938 and not w30939;
w30941 <= w6168 and not w28143;
w30942 <= w5598 and w27633;
w30943 <= w5874 and w27899;
w30944 <= not w30942 and not w30943;
w30945 <= not w30941 and w30944;
w30946 <= w5601 and not w28158;
w30947 <= w30945 and not w30946;
w30948 <= a(17) and not w30947;
w30949 <= a(17) and not w30948;
w30950 <= not w30947 and not w30948;
w30951 <= not w30949 and not w30950;
w30952 <= w30940 and not w30951;
w30953 <= w30940 and not w30952;
w30954 <= not w30951 and not w30952;
w30955 <= not w30953 and not w30954;
w30956 <= not w30814 and not w30819;
w30957 <= not w30955 and not w30956;
w30958 <= not w30955 and not w30957;
w30959 <= not w30956 and not w30957;
w30960 <= not w30958 and not w30959;
w30961 <= not w30821 and not w30824;
w30962 <= w30960 and w30961;
w30963 <= not w30960 and not w30961;
w30964 <= not w30962 and not w30963;
w30965 <= w30828 and not w30964;
w30966 <= not w30828 and w30964;
w30967 <= not w30965 and not w30966;
w30968 <= not w30864 and not w30877;
w30969 <= not w30855 and not w30858;
w30970 <= not w177 and w1188;
w30971 <= not w70 and w30970;
w30972 <= w311 and w1961;
w30973 <= w30971 and w30972;
w30974 <= w2198 and w30973;
w30975 <= w5123 and w30974;
w30976 <= w13182 and w30975;
w30977 <= w1035 and w30976;
w30978 <= w2441 and w30977;
w30979 <= w1716 and w30978;
w30980 <= w3674 and w30979;
w30981 <= w1315 and w30980;
w30982 <= not w1241 and w30981;
w30983 <= not w227 and w30982;
w30984 <= not w175 and w30983;
w30985 <= not w160 and w30984;
w30986 <= not w460 and w30985;
w30987 <= not w424 and w30986;
w30988 <= w30854 and not w30987;
w30989 <= not w30854 and w30987;
w30990 <= not w30969 and not w30989;
w30991 <= not w30988 and w30990;
w30992 <= not w30969 and not w30991;
w30993 <= not w30989 and not w30991;
w30994 <= not w30988 and w30993;
w30995 <= not w30992 and not w30994;
w30996 <= w10 and not w24551;
w30997 <= w2955 and w22261;
w30998 <= w2958 and w22267;
w30999 <= w2963 and w22264;
w31000 <= not w30998 and not w30999;
w31001 <= not w30997 and w31000;
w31002 <= not w30996 and w31001;
w31003 <= not w30995 and not w31002;
w31004 <= not w30995 and not w31003;
w31005 <= not w31002 and not w31003;
w31006 <= not w31004 and not w31005;
w31007 <= w3392 and w22247;
w31008 <= w3477 and w22258;
w31009 <= w3541 and w22255;
w31010 <= not w31008 and not w31009;
w31011 <= not w31007 and w31010;
w31012 <= not w3303 and w31011;
w31013 <= w25250 and w31011;
w31014 <= not w31012 and not w31013;
w31015 <= a(29) and not w31014;
w31016 <= not a(29) and w31014;
w31017 <= not w31015 and not w31016;
w31018 <= not w31006 and not w31017;
w31019 <= w31006 and w31017;
w31020 <= not w31018 and not w31019;
w31021 <= not w30968 and w31020;
w31022 <= w30968 and not w31020;
w31023 <= not w31021 and not w31022;
w31024 <= w3819 and w25998;
w31025 <= w3902 and w22250;
w31026 <= w3981 and w22244;
w31027 <= not w31025 and not w31026;
w31028 <= not w31024 and w31027;
w31029 <= w3985 and not w26539;
w31030 <= w31028 and not w31029;
w31031 <= a(26) and not w31030;
w31032 <= a(26) and not w31031;
w31033 <= not w31030 and not w31031;
w31034 <= not w31032 and not w31033;
w31035 <= w31023 and not w31034;
w31036 <= w31023 and not w31035;
w31037 <= not w31034 and not w31035;
w31038 <= not w31036 and not w31037;
w31039 <= not w30880 and not w30894;
w31040 <= w31038 and w31039;
w31041 <= not w31038 and not w31039;
w31042 <= not w31040 and not w31041;
w31043 <= w4629 and w26825;
w31044 <= w4468 and w26001;
w31045 <= w4539 and w25995;
w31046 <= not w31044 and not w31045;
w31047 <= not w31043 and w31046;
w31048 <= w4471 and not w26839;
w31049 <= w31047 and not w31048;
w31050 <= a(23) and not w31049;
w31051 <= a(23) and not w31050;
w31052 <= not w31049 and not w31050;
w31053 <= not w31051 and not w31052;
w31054 <= w31042 and not w31053;
w31055 <= w31042 and not w31054;
w31056 <= not w31053 and not w31054;
w31057 <= not w31055 and not w31056;
w31058 <= not w30900 and not w30913;
w31059 <= w31057 and w31058;
w31060 <= not w31057 and not w31058;
w31061 <= not w31059 and not w31060;
w31062 <= w5431 and w27633;
w31063 <= w4870 and w27108;
w31064 <= w5342 and w27377;
w31065 <= not w31063 and not w31064;
w31066 <= not w31062 and w31065;
w31067 <= w4873 and not w27648;
w31068 <= w31066 and not w31067;
w31069 <= a(20) and not w31068;
w31070 <= a(20) and not w31069;
w31071 <= not w31068 and not w31069;
w31072 <= not w31070 and not w31071;
w31073 <= w31061 and not w31072;
w31074 <= w31061 and not w31073;
w31075 <= not w31072 and not w31073;
w31076 <= not w31074 and not w31075;
w31077 <= not w30918 and not w30933;
w31078 <= not w13652 and not w28143;
w31079 <= w5598 and w27899;
w31080 <= not w31078 and not w31079;
w31081 <= not w5601 and w31080;
w31082 <= w28156 and w31080;
w31083 <= not w31081 and not w31082;
w31084 <= a(17) and not w31083;
w31085 <= not a(17) and w31083;
w31086 <= not w31084 and not w31085;
w31087 <= not w31077 and not w31086;
w31088 <= w31077 and w31086;
w31089 <= not w31087 and not w31088;
w31090 <= not w31076 and w31089;
w31091 <= not w31076 and not w31090;
w31092 <= w31089 and not w31090;
w31093 <= not w31091 and not w31092;
w31094 <= not w30939 and not w30952;
w31095 <= w31093 and w31094;
w31096 <= not w31093 and not w31094;
w31097 <= not w31095 and not w31096;
w31098 <= not w30957 and not w30963;
w31099 <= not w31097 and w31098;
w31100 <= w31097 and not w31098;
w31101 <= not w31099 and not w31100;
w31102 <= w30828 and w30964;
w31103 <= w31101 and w31102;
w31104 <= not w31101 and not w31102;
w31105 <= not w31103 and not w31104;
w31106 <= not w31096 and not w31100;
w31107 <= not w31087 and not w31090;
w31108 <= not w31041 and not w31054;
w31109 <= not w31021 and not w31035;
w31110 <= w3819 and w26001;
w31111 <= w3902 and w22244;
w31112 <= w3981 and w25998;
w31113 <= not w31111 and not w31112;
w31114 <= not w31110 and w31113;
w31115 <= w3985 and not w26559;
w31116 <= w31114 and not w31115;
w31117 <= a(26) and not w31116;
w31118 <= a(26) and not w31117;
w31119 <= not w31116 and not w31117;
w31120 <= not w31118 and not w31119;
w31121 <= not w31109 and not w31120;
w31122 <= not w31109 and not w31121;
w31123 <= not w31120 and not w31121;
w31124 <= not w31122 and not w31123;
w31125 <= not w31003 and not w31018;
w31126 <= w10 and w24534;
w31127 <= w2955 and w22258;
w31128 <= w2958 and w22264;
w31129 <= w2963 and w22261;
w31130 <= not w31128 and not w31129;
w31131 <= not w31127 and w31130;
w31132 <= not w31126 and w31131;
w31133 <= not w13654 and not w28143;
w31134 <= a(17) and not w31133;
w31135 <= not a(17) and w31133;
w31136 <= not w31134 and not w31135;
w31137 <= w1078 and w23976;
w31138 <= w2654 and w31137;
w31139 <= w4720 and w31138;
w31140 <= w3217 and w31139;
w31141 <= w12859 and w31140;
w31142 <= w817 and w31141;
w31143 <= w383 and w31142;
w31144 <= w214 and w31143;
w31145 <= not w164 and w31144;
w31146 <= not w270 and w31145;
w31147 <= not w234 and w31146;
w31148 <= not w460 and w31147;
w31149 <= not w706 and w31148;
w31150 <= w30987 and w31149;
w31151 <= not w30987 and not w31149;
w31152 <= not w31150 and not w31151;
w31153 <= w31136 and w31152;
w31154 <= not w31136 and not w31152;
w31155 <= not w31153 and not w31154;
w31156 <= not w31132 and w31155;
w31157 <= w31155 and not w31156;
w31158 <= not w31132 and not w31156;
w31159 <= not w31157 and not w31158;
w31160 <= not w30993 and not w31159;
w31161 <= not w31159 and not w31160;
w31162 <= not w30993 and not w31160;
w31163 <= not w31161 and not w31162;
w31164 <= not w31125 and not w31163;
w31165 <= not w31125 and not w31164;
w31166 <= not w31163 and not w31164;
w31167 <= not w31165 and not w31166;
w31168 <= w3392 and w22250;
w31169 <= w3477 and w22255;
w31170 <= w3541 and w22247;
w31171 <= not w31169 and not w31170;
w31172 <= not w31168 and w31171;
w31173 <= w3303 and w25229;
w31174 <= w31172 and not w31173;
w31175 <= a(29) and not w31174;
w31176 <= a(29) and not w31175;
w31177 <= not w31174 and not w31175;
w31178 <= not w31176 and not w31177;
w31179 <= not w31167 and not w31178;
w31180 <= not w31167 and not w31179;
w31181 <= not w31178 and not w31179;
w31182 <= not w31180 and not w31181;
w31183 <= not w31124 and w31182;
w31184 <= w31124 and not w31182;
w31185 <= not w31183 and not w31184;
w31186 <= w4629 and w27108;
w31187 <= w4468 and w25995;
w31188 <= w4539 and w26825;
w31189 <= not w31187 and not w31188;
w31190 <= not w31186 and w31189;
w31191 <= w4471 and w27120;
w31192 <= w31190 and not w31191;
w31193 <= a(23) and not w31192;
w31194 <= a(23) and not w31193;
w31195 <= not w31192 and not w31193;
w31196 <= not w31194 and not w31195;
w31197 <= not w31185 and not w31196;
w31198 <= w31185 and w31196;
w31199 <= not w31197 and not w31198;
w31200 <= w31108 and not w31199;
w31201 <= not w31108 and w31199;
w31202 <= not w31200 and not w31201;
w31203 <= not w31060 and not w31073;
w31204 <= w5431 and w27899;
w31205 <= w4870 and w27377;
w31206 <= w5342 and w27633;
w31207 <= not w31205 and not w31206;
w31208 <= not w31204 and w31207;
w31209 <= w4873 and w27911;
w31210 <= w31208 and not w31209;
w31211 <= a(20) and not w31210;
w31212 <= a(20) and not w31211;
w31213 <= not w31210 and not w31211;
w31214 <= not w31212 and not w31213;
w31215 <= not w31203 and not w31214;
w31216 <= not w31203 and not w31215;
w31217 <= not w31214 and not w31215;
w31218 <= not w31216 and not w31217;
w31219 <= not w31202 and w31218;
w31220 <= w31202 and not w31218;
w31221 <= not w31219 and not w31220;
w31222 <= not w31107 and w31221;
w31223 <= w31107 and not w31221;
w31224 <= not w31222 and not w31223;
w31225 <= not w31106 and w31224;
w31226 <= w31106 and not w31224;
w31227 <= not w31225 and not w31226;
w31228 <= not w31103 and not w31227;
w31229 <= w31103 and w31227;
w31230 <= not w31228 and not w31229;
w31231 <= not w31164 and not w31179;
w31232 <= w10 and not w25205;
w31233 <= w2955 and w22255;
w31234 <= w2958 and w22261;
w31235 <= w2963 and w22258;
w31236 <= not w31234 and not w31235;
w31237 <= not w31233 and w31236;
w31238 <= not w31232 and w31237;
w31239 <= not w31151 and not w31153;
w31240 <= w567 and w12949;
w31241 <= w2591 and w31240;
w31242 <= w6449 and w31241;
w31243 <= w2478 and w31242;
w31244 <= w3432 and w31243;
w31245 <= w29485 and w31244;
w31246 <= w358 and w31245;
w31247 <= w353 and w31246;
w31248 <= w4036 and w31247;
w31249 <= not w265 and w31248;
w31250 <= not w264 and w31249;
w31251 <= not w215 and w31250;
w31252 <= not w138 and w31251;
w31253 <= not w554 and w31252;
w31254 <= not w471 and w31253;
w31255 <= not w31239 and w31254;
w31256 <= w31239 and not w31254;
w31257 <= not w31255 and not w31256;
w31258 <= not w31238 and w31257;
w31259 <= not w31238 and not w31258;
w31260 <= w31257 and not w31258;
w31261 <= not w31259 and not w31260;
w31262 <= not w31156 and not w31160;
w31263 <= w31261 and w31262;
w31264 <= not w31261 and not w31262;
w31265 <= not w31263 and not w31264;
w31266 <= w3392 and w22244;
w31267 <= w3477 and w22247;
w31268 <= w3541 and w22250;
w31269 <= not w31267 and not w31268;
w31270 <= not w31266 and w31269;
w31271 <= not w3303 and w31270;
w31272 <= w22464 and w31270;
w31273 <= not w31271 and not w31272;
w31274 <= a(29) and not w31273;
w31275 <= not a(29) and w31273;
w31276 <= not w31274 and not w31275;
w31277 <= w31265 and not w31276;
w31278 <= not w31265 and w31276;
w31279 <= not w31277 and not w31278;
w31280 <= not w31231 and w31279;
w31281 <= w31231 and not w31279;
w31282 <= not w31280 and not w31281;
w31283 <= w3819 and w25995;
w31284 <= w3902 and w25998;
w31285 <= w3981 and w26001;
w31286 <= not w31284 and not w31285;
w31287 <= not w31283 and w31286;
w31288 <= w3985 and not w26023;
w31289 <= w31287 and not w31288;
w31290 <= a(26) and not w31289;
w31291 <= a(26) and not w31290;
w31292 <= not w31289 and not w31290;
w31293 <= not w31291 and not w31292;
w31294 <= w31282 and not w31293;
w31295 <= w31282 and not w31294;
w31296 <= not w31293 and not w31294;
w31297 <= not w31295 and not w31296;
w31298 <= not w31124 and not w31182;
w31299 <= not w31121 and not w31298;
w31300 <= not w31297 and not w31299;
w31301 <= not w31297 and not w31300;
w31302 <= not w31299 and not w31300;
w31303 <= not w31301 and not w31302;
w31304 <= w4629 and w27377;
w31305 <= w4468 and w26825;
w31306 <= w4539 and w27108;
w31307 <= not w31305 and not w31306;
w31308 <= not w31304 and w31307;
w31309 <= w4471 and w27390;
w31310 <= w31308 and not w31309;
w31311 <= a(23) and not w31310;
w31312 <= a(23) and not w31311;
w31313 <= not w31310 and not w31311;
w31314 <= not w31312 and not w31313;
w31315 <= not w31303 and not w31314;
w31316 <= not w31303 and not w31315;
w31317 <= not w31314 and not w31315;
w31318 <= not w31316 and not w31317;
w31319 <= not w31197 and not w31201;
w31320 <= w31318 and w31319;
w31321 <= not w31318 and not w31319;
w31322 <= not w31320 and not w31321;
w31323 <= w5431 and not w28143;
w31324 <= w4870 and w27633;
w31325 <= w5342 and w27899;
w31326 <= not w31324 and not w31325;
w31327 <= not w31323 and w31326;
w31328 <= w4873 and not w28158;
w31329 <= w31327 and not w31328;
w31330 <= a(20) and not w31329;
w31331 <= a(20) and not w31330;
w31332 <= not w31329 and not w31330;
w31333 <= not w31331 and not w31332;
w31334 <= w31322 and not w31333;
w31335 <= w31322 and not w31334;
w31336 <= not w31333 and not w31334;
w31337 <= not w31335 and not w31336;
w31338 <= not w31215 and not w31220;
w31339 <= not w31337 and not w31338;
w31340 <= not w31337 and not w31339;
w31341 <= not w31338 and not w31339;
w31342 <= not w31340 and not w31341;
w31343 <= not w31222 and not w31225;
w31344 <= w31342 and w31343;
w31345 <= not w31342 and not w31343;
w31346 <= not w31344 and not w31345;
w31347 <= not w31229 and w31346;
w31348 <= w31229 and not w31346;
w31349 <= not w31347 and not w31348;
w31350 <= w31229 and w31346;
w31351 <= w10 and not w25250;
w31352 <= w2955 and w22247;
w31353 <= w2958 and w22258;
w31354 <= w2963 and w22255;
w31355 <= not w31353 and not w31354;
w31356 <= not w31352 and w31355;
w31357 <= not w31351 and w31356;
w31358 <= w12876 and w30971;
w31359 <= w4301 and w31358;
w31360 <= w6496 and w31359;
w31361 <= w3194 and w31360;
w31362 <= w2586 and w31361;
w31363 <= w2618 and w31362;
w31364 <= w165 and w31363;
w31365 <= w423 and w31364;
w31366 <= w28623 and w31365;
w31367 <= not w537 and w31366;
w31368 <= not w1036 and w31367;
w31369 <= not w77 and w31368;
w31370 <= not w60 and w31369;
w31371 <= not w31254 and w31370;
w31372 <= w31254 and not w31370;
w31373 <= not w31357 and not w31372;
w31374 <= not w31371 and w31373;
w31375 <= not w31357 and not w31374;
w31376 <= not w31372 and not w31374;
w31377 <= not w31371 and w31376;
w31378 <= not w31375 and not w31377;
w31379 <= not w31255 and not w31258;
w31380 <= w31378 and w31379;
w31381 <= not w31378 and not w31379;
w31382 <= not w31380 and not w31381;
w31383 <= not w31264 and not w31277;
w31384 <= not w31382 and w31383;
w31385 <= w31382 and not w31383;
w31386 <= not w31384 and not w31385;
w31387 <= w3392 and w25998;
w31388 <= w3477 and w22250;
w31389 <= w3541 and w22244;
w31390 <= not w31388 and not w31389;
w31391 <= not w31387 and w31390;
w31392 <= w3303 and not w26539;
w31393 <= w31391 and not w31392;
w31394 <= a(29) and not w31393;
w31395 <= a(29) and not w31394;
w31396 <= not w31393 and not w31394;
w31397 <= not w31395 and not w31396;
w31398 <= w31386 and not w31397;
w31399 <= w31386 and not w31398;
w31400 <= not w31397 and not w31398;
w31401 <= not w31399 and not w31400;
w31402 <= w3819 and w26825;
w31403 <= w3902 and w26001;
w31404 <= w3981 and w25995;
w31405 <= not w31403 and not w31404;
w31406 <= not w31402 and w31405;
w31407 <= w3985 and not w26839;
w31408 <= w31406 and not w31407;
w31409 <= a(26) and not w31408;
w31410 <= a(26) and not w31409;
w31411 <= not w31408 and not w31409;
w31412 <= not w31410 and not w31411;
w31413 <= not w31401 and not w31412;
w31414 <= not w31401 and not w31413;
w31415 <= not w31412 and not w31413;
w31416 <= not w31414 and not w31415;
w31417 <= not w31280 and not w31294;
w31418 <= w31416 and w31417;
w31419 <= not w31416 and not w31417;
w31420 <= not w31418 and not w31419;
w31421 <= w4629 and w27633;
w31422 <= w4468 and w27108;
w31423 <= w4539 and w27377;
w31424 <= not w31422 and not w31423;
w31425 <= not w31421 and w31424;
w31426 <= w4471 and not w27648;
w31427 <= w31425 and not w31426;
w31428 <= a(23) and not w31427;
w31429 <= a(23) and not w31428;
w31430 <= not w31427 and not w31428;
w31431 <= not w31429 and not w31430;
w31432 <= w31420 and not w31431;
w31433 <= w31420 and not w31432;
w31434 <= not w31431 and not w31432;
w31435 <= not w31433 and not w31434;
w31436 <= not w31300 and not w31315;
w31437 <= not w13374 and not w28143;
w31438 <= w4870 and w27899;
w31439 <= not w31437 and not w31438;
w31440 <= not w4873 and w31439;
w31441 <= w28156 and w31439;
w31442 <= not w31440 and not w31441;
w31443 <= a(20) and not w31442;
w31444 <= not a(20) and w31442;
w31445 <= not w31443 and not w31444;
w31446 <= not w31436 and not w31445;
w31447 <= w31436 and w31445;
w31448 <= not w31446 and not w31447;
w31449 <= not w31435 and w31448;
w31450 <= not w31435 and not w31449;
w31451 <= w31448 and not w31449;
w31452 <= not w31450 and not w31451;
w31453 <= not w31321 and not w31334;
w31454 <= w31452 and w31453;
w31455 <= not w31452 and not w31453;
w31456 <= not w31454 and not w31455;
w31457 <= not w31339 and not w31345;
w31458 <= not w31456 and w31457;
w31459 <= w31456 and not w31457;
w31460 <= not w31458 and not w31459;
w31461 <= w31350 and w31460;
w31462 <= not w31350 and not w31460;
w31463 <= not w31461 and not w31462;
w31464 <= not w31455 and not w31459;
w31465 <= not w31446 and not w31449;
w31466 <= w10 and w25229;
w31467 <= w2955 and w22250;
w31468 <= w2958 and w22255;
w31469 <= w2963 and w22247;
w31470 <= not w31468 and not w31469;
w31471 <= not w31467 and w31470;
w31472 <= not w31466 and w31471;
w31473 <= not w13376 and not w28143;
w31474 <= a(20) and not w31473;
w31475 <= not a(20) and w31473;
w31476 <= not w31474 and not w31475;
w31477 <= w2688 and w3305;
w31478 <= w465 and w31477;
w31479 <= w14985 and w31478;
w31480 <= w15888 and w31479;
w31481 <= w4228 and w31480;
w31482 <= w943 and w31481;
w31483 <= w740 and w31482;
w31484 <= w474 and w31483;
w31485 <= w2441 and w31484;
w31486 <= w550 and w31485;
w31487 <= w1509 and w31486;
w31488 <= not w493 and w31487;
w31489 <= not w355 and w31488;
w31490 <= not w124 and w31489;
w31491 <= not w651 and w31490;
w31492 <= not w387 and w31491;
w31493 <= not w136 and w31492;
w31494 <= w31254 and w31493;
w31495 <= not w31254 and not w31493;
w31496 <= not w31494 and not w31495;
w31497 <= w31476 and w31496;
w31498 <= not w31476 and not w31496;
w31499 <= not w31497 and not w31498;
w31500 <= not w31376 and w31499;
w31501 <= w31376 and not w31499;
w31502 <= not w31500 and not w31501;
w31503 <= not w31472 and w31502;
w31504 <= w31502 and not w31503;
w31505 <= not w31472 and not w31503;
w31506 <= not w31504 and not w31505;
w31507 <= not w31381 and not w31385;
w31508 <= w31506 and w31507;
w31509 <= not w31506 and not w31507;
w31510 <= not w31508 and not w31509;
w31511 <= w3392 and w26001;
w31512 <= w3477 and w22244;
w31513 <= w3541 and w25998;
w31514 <= not w31512 and not w31513;
w31515 <= not w31511 and w31514;
w31516 <= w3303 and not w26559;
w31517 <= w31515 and not w31516;
w31518 <= a(29) and not w31517;
w31519 <= a(29) and not w31518;
w31520 <= not w31517 and not w31518;
w31521 <= not w31519 and not w31520;
w31522 <= w31510 and not w31521;
w31523 <= w31510 and not w31522;
w31524 <= not w31521 and not w31522;
w31525 <= not w31523 and not w31524;
w31526 <= w3819 and w27108;
w31527 <= w3902 and w25995;
w31528 <= w3981 and w26825;
w31529 <= not w31527 and not w31528;
w31530 <= not w31526 and w31529;
w31531 <= w3985 and w27120;
w31532 <= w31530 and not w31531;
w31533 <= a(26) and not w31532;
w31534 <= a(26) and not w31533;
w31535 <= not w31532 and not w31533;
w31536 <= not w31534 and not w31535;
w31537 <= not w31525 and not w31536;
w31538 <= not w31525 and not w31537;
w31539 <= not w31536 and not w31537;
w31540 <= not w31538 and not w31539;
w31541 <= not w31398 and not w31413;
w31542 <= w31540 and w31541;
w31543 <= not w31540 and not w31541;
w31544 <= not w31542 and not w31543;
w31545 <= not w31419 and not w31432;
w31546 <= w4629 and w27899;
w31547 <= w4468 and w27377;
w31548 <= w4539 and w27633;
w31549 <= not w31547 and not w31548;
w31550 <= not w31546 and w31549;
w31551 <= w4471 and w27911;
w31552 <= w31550 and not w31551;
w31553 <= a(23) and not w31552;
w31554 <= a(23) and not w31553;
w31555 <= not w31552 and not w31553;
w31556 <= not w31554 and not w31555;
w31557 <= not w31545 and not w31556;
w31558 <= not w31545 and not w31557;
w31559 <= not w31556 and not w31557;
w31560 <= not w31558 and not w31559;
w31561 <= not w31544 and w31560;
w31562 <= w31544 and not w31560;
w31563 <= not w31561 and not w31562;
w31564 <= not w31465 and w31563;
w31565 <= w31465 and not w31563;
w31566 <= not w31564 and not w31565;
w31567 <= not w31464 and w31566;
w31568 <= w31464 and not w31566;
w31569 <= not w31567 and not w31568;
w31570 <= not w31461 and not w31569;
w31571 <= w31461 and w31569;
w31572 <= not w31570 and not w31571;
w31573 <= not w31509 and not w31522;
w31574 <= w10 and not w22464;
w31575 <= w2955 and w22244;
w31576 <= w2958 and w22247;
w31577 <= w2963 and w22250;
w31578 <= not w31576 and not w31577;
w31579 <= not w31575 and w31578;
w31580 <= not w31574 and w31579;
w31581 <= not w31495 and not w31497;
w31582 <= w1675 and w4763;
w31583 <= w1539 and w31582;
w31584 <= w1575 and w31583;
w31585 <= w14469 and w31584;
w31586 <= w964 and w31585;
w31587 <= w3217 and w31586;
w31588 <= w1614 and w31587;
w31589 <= w2974 and w31588;
w31590 <= w15990 and w31589;
w31591 <= w1187 and w31590;
w31592 <= not w1181 and w31591;
w31593 <= not w537 and w31592;
w31594 <= not w80 and w31593;
w31595 <= not w233 and w31594;
w31596 <= not w157 and w31595;
w31597 <= not w31581 and w31596;
w31598 <= w31581 and not w31596;
w31599 <= not w31597 and not w31598;
w31600 <= not w31580 and w31599;
w31601 <= not w31580 and not w31600;
w31602 <= w31599 and not w31600;
w31603 <= not w31601 and not w31602;
w31604 <= not w31500 and not w31503;
w31605 <= w31603 and w31604;
w31606 <= not w31603 and not w31604;
w31607 <= not w31605 and not w31606;
w31608 <= w3392 and w25995;
w31609 <= w3477 and w25998;
w31610 <= w3541 and w26001;
w31611 <= not w31609 and not w31610;
w31612 <= not w31608 and w31611;
w31613 <= not w3303 and w31612;
w31614 <= w26023 and w31612;
w31615 <= not w31613 and not w31614;
w31616 <= a(29) and not w31615;
w31617 <= not a(29) and w31615;
w31618 <= not w31616 and not w31617;
w31619 <= w31607 and not w31618;
w31620 <= not w31607 and w31618;
w31621 <= not w31619 and not w31620;
w31622 <= not w31573 and w31621;
w31623 <= w31573 and not w31621;
w31624 <= not w31622 and not w31623;
w31625 <= w3819 and w27377;
w31626 <= w3902 and w26825;
w31627 <= w3981 and w27108;
w31628 <= not w31626 and not w31627;
w31629 <= not w31625 and w31628;
w31630 <= w3985 and w27390;
w31631 <= w31629 and not w31630;
w31632 <= a(26) and not w31631;
w31633 <= a(26) and not w31632;
w31634 <= not w31631 and not w31632;
w31635 <= not w31633 and not w31634;
w31636 <= w31624 and not w31635;
w31637 <= w31624 and not w31636;
w31638 <= not w31635 and not w31636;
w31639 <= not w31637 and not w31638;
w31640 <= not w31537 and not w31543;
w31641 <= w31639 and w31640;
w31642 <= not w31639 and not w31640;
w31643 <= not w31641 and not w31642;
w31644 <= w4629 and not w28143;
w31645 <= w4468 and w27633;
w31646 <= w4539 and w27899;
w31647 <= not w31645 and not w31646;
w31648 <= not w31644 and w31647;
w31649 <= w4471 and not w28158;
w31650 <= w31648 and not w31649;
w31651 <= a(23) and not w31650;
w31652 <= a(23) and not w31651;
w31653 <= not w31650 and not w31651;
w31654 <= not w31652 and not w31653;
w31655 <= w31643 and not w31654;
w31656 <= w31643 and not w31655;
w31657 <= not w31654 and not w31655;
w31658 <= not w31656 and not w31657;
w31659 <= not w31557 and not w31562;
w31660 <= not w31658 and not w31659;
w31661 <= not w31658 and not w31660;
w31662 <= not w31659 and not w31660;
w31663 <= not w31661 and not w31662;
w31664 <= not w31564 and not w31567;
w31665 <= w31663 and w31664;
w31666 <= not w31663 and not w31664;
w31667 <= not w31665 and not w31666;
w31668 <= w31571 and not w31667;
w31669 <= not w31571 and w31667;
w31670 <= not w31668 and not w31669;
w31671 <= not w31597 and not w31600;
w31672 <= w3394 and w12951;
w31673 <= w1005 and w31672;
w31674 <= w15817 and w31673;
w31675 <= w25798 and w31674;
w31676 <= w4167 and w31675;
w31677 <= w2586 and w31676;
w31678 <= w29473 and w31677;
w31679 <= w220 and w31678;
w31680 <= w1187 and w31679;
w31681 <= w655 and w31680;
w31682 <= w22697 and w31681;
w31683 <= not w269 and w31682;
w31684 <= not w168 and w31683;
w31685 <= not w237 and w31684;
w31686 <= not w649 and w31685;
w31687 <= w31596 and not w31686;
w31688 <= not w31596 and w31686;
w31689 <= not w31671 and not w31688;
w31690 <= not w31687 and w31689;
w31691 <= not w31671 and not w31690;
w31692 <= not w31688 and not w31690;
w31693 <= not w31687 and w31692;
w31694 <= not w31691 and not w31693;
w31695 <= w10 and not w26539;
w31696 <= w2955 and w25998;
w31697 <= w2958 and w22250;
w31698 <= w2963 and w22244;
w31699 <= not w31697 and not w31698;
w31700 <= not w31696 and w31699;
w31701 <= not w31695 and w31700;
w31702 <= not w31694 and not w31701;
w31703 <= not w31694 and not w31702;
w31704 <= not w31701 and not w31702;
w31705 <= not w31703 and not w31704;
w31706 <= not w31606 and not w31619;
w31707 <= w31705 and w31706;
w31708 <= not w31705 and not w31706;
w31709 <= not w31707 and not w31708;
w31710 <= w3392 and w26825;
w31711 <= w3477 and w26001;
w31712 <= w3541 and w25995;
w31713 <= not w31711 and not w31712;
w31714 <= not w31710 and w31713;
w31715 <= w3303 and not w26839;
w31716 <= w31714 and not w31715;
w31717 <= a(29) and not w31716;
w31718 <= a(29) and not w31717;
w31719 <= not w31716 and not w31717;
w31720 <= not w31718 and not w31719;
w31721 <= w31709 and not w31720;
w31722 <= w31709 and not w31721;
w31723 <= not w31720 and not w31721;
w31724 <= not w31722 and not w31723;
w31725 <= w3819 and w27633;
w31726 <= w3902 and w27108;
w31727 <= w3981 and w27377;
w31728 <= not w31726 and not w31727;
w31729 <= not w31725 and w31728;
w31730 <= w3985 and not w27648;
w31731 <= w31729 and not w31730;
w31732 <= a(26) and not w31731;
w31733 <= a(26) and not w31732;
w31734 <= not w31731 and not w31732;
w31735 <= not w31733 and not w31734;
w31736 <= not w31724 and not w31735;
w31737 <= not w31724 and not w31736;
w31738 <= not w31735 and not w31736;
w31739 <= not w31737 and not w31738;
w31740 <= not w31622 and not w31636;
w31741 <= not w13873 and not w28143;
w31742 <= w4468 and w27899;
w31743 <= not w31741 and not w31742;
w31744 <= not w4471 and w31743;
w31745 <= w28156 and w31743;
w31746 <= not w31744 and not w31745;
w31747 <= a(23) and not w31746;
w31748 <= not a(23) and w31746;
w31749 <= not w31747 and not w31748;
w31750 <= not w31740 and not w31749;
w31751 <= w31740 and w31749;
w31752 <= not w31750 and not w31751;
w31753 <= not w31739 and w31752;
w31754 <= not w31739 and not w31753;
w31755 <= w31752 and not w31753;
w31756 <= not w31754 and not w31755;
w31757 <= not w31642 and not w31655;
w31758 <= w31756 and w31757;
w31759 <= not w31756 and not w31757;
w31760 <= not w31758 and not w31759;
w31761 <= not w31660 and not w31666;
w31762 <= not w31760 and w31761;
w31763 <= w31760 and not w31761;
w31764 <= not w31762 and not w31763;
w31765 <= w31571 and w31667;
w31766 <= w31764 and w31765;
w31767 <= not w31764 and not w31765;
w31768 <= not w31766 and not w31767;
w31769 <= not w31759 and not w31763;
w31770 <= not w31750 and not w31753;
w31771 <= not w31721 and not w31736;
w31772 <= w3819 and w27899;
w31773 <= w3902 and w27377;
w31774 <= w3981 and w27633;
w31775 <= not w31773 and not w31774;
w31776 <= not w31772 and w31775;
w31777 <= w3985 and w27911;
w31778 <= w31776 and not w31777;
w31779 <= a(26) and not w31778;
w31780 <= a(26) and not w31779;
w31781 <= not w31778 and not w31779;
w31782 <= not w31780 and not w31781;
w31783 <= not w31771 and not w31782;
w31784 <= not w31771 and not w31783;
w31785 <= not w31782 and not w31783;
w31786 <= not w31784 and not w31785;
w31787 <= w10 and not w26559;
w31788 <= w2955 and w26001;
w31789 <= w2958 and w22244;
w31790 <= w2963 and w25998;
w31791 <= not w31789 and not w31790;
w31792 <= not w31788 and w31791;
w31793 <= not w31787 and w31792;
w31794 <= not w22183 and not w28143;
w31795 <= a(23) and not w31794;
w31796 <= not a(23) and w31794;
w31797 <= not w31795 and not w31796;
w31798 <= w4734 and w13096;
w31799 <= w1090 and w31798;
w31800 <= w3938 and w31799;
w31801 <= w3801 and w31800;
w31802 <= w223 and w31801;
w31803 <= w872 and w31802;
w31804 <= w1413 and w31803;
w31805 <= w128 and w31804;
w31806 <= not w444 and w31805;
w31807 <= not w946 and w31806;
w31808 <= not w163 and w31807;
w31809 <= not w760 and w31808;
w31810 <= not w503 and w31809;
w31811 <= not w454 and w31810;
w31812 <= w31686 and w31811;
w31813 <= not w31686 and not w31811;
w31814 <= not w31812 and not w31813;
w31815 <= w31797 and w31814;
w31816 <= not w31797 and not w31814;
w31817 <= not w31815 and not w31816;
w31818 <= not w31692 and w31817;
w31819 <= w31692 and not w31817;
w31820 <= not w31818 and not w31819;
w31821 <= not w31793 and w31820;
w31822 <= w31820 and not w31821;
w31823 <= not w31793 and not w31821;
w31824 <= not w31822 and not w31823;
w31825 <= not w31702 and not w31708;
w31826 <= w31824 and w31825;
w31827 <= not w31824 and not w31825;
w31828 <= not w31826 and not w31827;
w31829 <= w3392 and w27108;
w31830 <= w3477 and w25995;
w31831 <= w3541 and w26825;
w31832 <= not w31830 and not w31831;
w31833 <= not w31829 and w31832;
w31834 <= w3303 and w27120;
w31835 <= w31833 and not w31834;
w31836 <= a(29) and not w31835;
w31837 <= a(29) and not w31836;
w31838 <= not w31835 and not w31836;
w31839 <= not w31837 and not w31838;
w31840 <= w31828 and not w31839;
w31841 <= w31828 and not w31840;
w31842 <= not w31839 and not w31840;
w31843 <= not w31841 and not w31842;
w31844 <= not w31786 and w31843;
w31845 <= w31786 and not w31843;
w31846 <= not w31844 and not w31845;
w31847 <= not w31770 and not w31846;
w31848 <= w31770 and w31846;
w31849 <= not w31847 and not w31848;
w31850 <= not w31769 and w31849;
w31851 <= w31769 and not w31849;
w31852 <= not w31850 and not w31851;
w31853 <= not w31766 and not w31852;
w31854 <= w31766 and w31852;
w31855 <= not w31853 and not w31854;
w31856 <= not w31827 and not w31840;
w31857 <= w10 and not w26023;
w31858 <= w2955 and w25995;
w31859 <= w2958 and w25998;
w31860 <= w2963 and w26001;
w31861 <= not w31859 and not w31860;
w31862 <= not w31858 and w31861;
w31863 <= not w31857 and w31862;
w31864 <= not w31813 and not w31815;
w31865 <= w1673 and w14947;
w31866 <= w3373 and w31865;
w31867 <= w6545 and w31866;
w31868 <= w25951 and w31867;
w31869 <= w15815 and w31868;
w31870 <= w3874 and w31869;
w31871 <= w3932 and w31870;
w31872 <= w1118 and w31871;
w31873 <= w1466 and w31872;
w31874 <= w1301 and w31873;
w31875 <= w1718 and w31874;
w31876 <= w35 and w31875;
w31877 <= not w355 and w31876;
w31878 <= not w401 and w31877;
w31879 <= not w233 and w31878;
w31880 <= not w186 and w31879;
w31881 <= not w31864 and w31880;
w31882 <= w31864 and not w31880;
w31883 <= not w31881 and not w31882;
w31884 <= not w31863 and w31883;
w31885 <= not w31863 and not w31884;
w31886 <= w31883 and not w31884;
w31887 <= not w31885 and not w31886;
w31888 <= not w31818 and not w31821;
w31889 <= w31887 and w31888;
w31890 <= not w31887 and not w31888;
w31891 <= not w31889 and not w31890;
w31892 <= w3392 and w27377;
w31893 <= w3477 and w26825;
w31894 <= w3541 and w27108;
w31895 <= not w31893 and not w31894;
w31896 <= not w31892 and w31895;
w31897 <= not w3303 and w31896;
w31898 <= not w27390 and w31896;
w31899 <= not w31897 and not w31898;
w31900 <= a(29) and not w31899;
w31901 <= not a(29) and w31899;
w31902 <= not w31900 and not w31901;
w31903 <= w31891 and not w31902;
w31904 <= not w31891 and w31902;
w31905 <= not w31903 and not w31904;
w31906 <= not w31856 and w31905;
w31907 <= w31856 and not w31905;
w31908 <= not w31906 and not w31907;
w31909 <= w3819 and not w28143;
w31910 <= w3902 and w27633;
w31911 <= w3981 and w27899;
w31912 <= not w31910 and not w31911;
w31913 <= not w31909 and w31912;
w31914 <= w3985 and not w28158;
w31915 <= w31913 and not w31914;
w31916 <= a(26) and not w31915;
w31917 <= a(26) and not w31916;
w31918 <= not w31915 and not w31916;
w31919 <= not w31917 and not w31918;
w31920 <= w31908 and not w31919;
w31921 <= w31908 and not w31920;
w31922 <= not w31919 and not w31920;
w31923 <= not w31921 and not w31922;
w31924 <= not w31786 and not w31843;
w31925 <= not w31783 and not w31924;
w31926 <= not w31923 and not w31925;
w31927 <= not w31923 and not w31926;
w31928 <= not w31925 and not w31926;
w31929 <= not w31927 and not w31928;
w31930 <= not w31847 and not w31850;
w31931 <= w31929 and w31930;
w31932 <= not w31929 and not w31930;
w31933 <= not w31931 and not w31932;
w31934 <= not w31854 and w31933;
w31935 <= w31854 and not w31933;
w31936 <= not w31934 and not w31935;
w31937 <= w31854 and w31933;
w31938 <= not w31926 and not w31932;
w31939 <= not w31906 and not w31920;
w31940 <= not w31881 and not w31884;
w31941 <= w3944 and w13010;
w31942 <= w3783 and w31941;
w31943 <= w3774 and w31942;
w31944 <= w2208 and w31943;
w31945 <= w25951 and w31944;
w31946 <= w3919 and w31945;
w31947 <= not w760 and w31946;
w31948 <= not w31880 and w31947;
w31949 <= w31880 and not w31947;
w31950 <= not w31940 and not w31949;
w31951 <= not w31948 and w31950;
w31952 <= not w31940 and not w31951;
w31953 <= not w31949 and not w31951;
w31954 <= not w31948 and w31953;
w31955 <= not w31952 and not w31954;
w31956 <= w10 and not w26839;
w31957 <= w2955 and w26825;
w31958 <= w2958 and w26001;
w31959 <= w2963 and w25995;
w31960 <= not w31958 and not w31959;
w31961 <= not w31957 and w31960;
w31962 <= not w31956 and w31961;
w31963 <= not w31955 and not w31962;
w31964 <= not w31955 and not w31963;
w31965 <= not w31962 and not w31963;
w31966 <= not w31964 and not w31965;
w31967 <= not w31890 and not w31903;
w31968 <= w31966 and w31967;
w31969 <= not w31966 and not w31967;
w31970 <= not w31968 and not w31969;
w31971 <= not w25892 and not w28143;
w31972 <= w3902 and w27899;
w31973 <= not w31971 and not w31972;
w31974 <= w3985 and not w28156;
w31975 <= w31973 and not w31974;
w31976 <= a(26) and not w31975;
w31977 <= not w31975 and not w31976;
w31978 <= a(26) and not w31976;
w31979 <= not w31977 and not w31978;
w31980 <= w3392 and w27633;
w31981 <= w3477 and w27108;
w31982 <= w3541 and w27377;
w31983 <= not w31981 and not w31982;
w31984 <= not w31980 and w31983;
w31985 <= w3303 and not w27648;
w31986 <= w31984 and not w31985;
w31987 <= a(29) and not w31986;
w31988 <= a(29) and not w31987;
w31989 <= not w31986 and not w31987;
w31990 <= not w31988 and not w31989;
w31991 <= not w31979 and not w31990;
w31992 <= not w31979 and not w31991;
w31993 <= not w31990 and not w31991;
w31994 <= not w31992 and not w31993;
w31995 <= not w31970 and w31994;
w31996 <= w31970 and not w31994;
w31997 <= not w31995 and not w31996;
w31998 <= not w31939 and w31997;
w31999 <= w31939 and not w31997;
w32000 <= not w31998 and not w31999;
w32001 <= not w31938 and w32000;
w32002 <= w31938 and not w32000;
w32003 <= not w32001 and not w32002;
w32004 <= not w31937 and not w32003;
w32005 <= w31937 and w32003;
w32006 <= not w32004 and not w32005;
w32007 <= not w31998 and not w32001;
w32008 <= w3392 and w27899;
w32009 <= w3477 and w27377;
w32010 <= w3541 and w27633;
w32011 <= not w32009 and not w32010;
w32012 <= not w32008 and w32011;
w32013 <= w3303 and w27911;
w32014 <= w32012 and not w32013;
w32015 <= not w31963 and not w31969;
w32016 <= a(29) and not w32015;
w32017 <= not a(29) and w32015;
w32018 <= not w32016 and not w32017;
w32019 <= w32014 and w32018;
w32020 <= not w32014 and not w32018;
w32021 <= not w32019 and not w32020;
w32022 <= w10 and w27120;
w32023 <= w2955 and w27108;
w32024 <= w2958 and w25995;
w32025 <= w2963 and w26825;
w32026 <= not w32024 and not w32025;
w32027 <= not w32023 and w32026;
w32028 <= not w32022 and w32027;
w32029 <= w31953 and not w32028;
w32030 <= not w31953 and w32028;
w32031 <= not w32029 and not w32030;
w32032 <= w32021 and not w32031;
w32033 <= not w32021 and w32031;
w32034 <= not w32032 and not w32033;
w32035 <= not w31991 and not w31996;
w32036 <= w3809 and w4446;
w32037 <= not w536 and w32036;
w32038 <= a(26) and not w32037;
w32039 <= not a(26) and w32037;
w32040 <= not w32038 and not w32039;
w32041 <= not w25945 and not w28143;
w32042 <= w31880 and not w32041;
w32043 <= not w31880 and w32041;
w32044 <= not w32042 and not w32043;
w32045 <= w32040 and w32044;
w32046 <= not w32040 and not w32044;
w32047 <= not w32045 and not w32046;
w32048 <= w32035 and not w32047;
w32049 <= not w32035 and w32047;
w32050 <= not w32048 and not w32049;
w32051 <= w32034 and w32050;
w32052 <= not w32034 and not w32050;
w32053 <= not w32051 and not w32052;
w32054 <= not w32007 and not w32053;
w32055 <= w32007 and w32053;
w32056 <= not w32054 and not w32055;
w32057 <= w32005 and w32056;
w32058 <= not w32005 and not w32056;
w32059 <= not w32057 and not w32058;
one <= '1';
result(0) <= not w26856;-- level 360
result(1) <= w27134;-- level 362
result(2) <= w27404;-- level 364
result(3) <= w27662;-- level 366
result(4) <= w27925;-- level 368
result(5) <= w28172;-- level 370
result(6) <= w28401;-- level 372
result(7) <= w28619;-- level 393
result(8) <= w28838;-- level 398
result(9) <= w29049;-- level 400
result(10) <= w29252;-- level 402
result(11) <= not w29463;-- level 404
result(12) <= w29675;-- level 406
result(13) <= w29857;-- level 408
result(14) <= not w30032;-- level 410
result(15) <= w30208;-- level 412
result(16) <= w30375;-- level 414
result(17) <= not w30531;-- level 416
result(18) <= w30687;-- level 418
result(19) <= w30829;-- level 420
result(20) <= not w30967;-- level 422
result(21) <= w31105;-- level 424
result(22) <= w31230;-- level 426
result(23) <= not w31349;-- level 428
result(24) <= w31463;-- level 430
result(25) <= w31572;-- level 432
result(26) <= not w31670;-- level 434
result(27) <= w31768;-- level 436
result(28) <= w31855;-- level 438
result(29) <= not w31936;-- level 440
result(30) <= w32006;-- level 442
result(31) <= not w32059;-- level 444
end Behavioral;