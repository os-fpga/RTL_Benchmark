-------------------------------------------------------------------------------
--
-- GCpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: gcpad_ctrl-c.vhd,v 1.1 2004-10-07 21:23:10 arniml Exp $
--
-------------------------------------------------------------------------------

configuration gcpad_ctrl_rtl_c0 of gcpad_ctrl is

  for rtl
  end for;

end gcpad_ctrl_rtl_c0;
