module AF_IO_H (
	inout		PAD,
	input		DIN,
	output		DOUT,
	input		OE,
	input		PUD,
	input		PE,
	input		DS0,
	input		DS1
	);
endmodule
