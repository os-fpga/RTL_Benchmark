
class apb_env_config extends uvm_object;
	`uvm_object_utils(apb_env_config)

function new(string name);
	super.new(name);
endfunction
