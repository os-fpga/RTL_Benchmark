module top ( 
    \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] , \B[8] ,
    \B[9] , \B[10] ,
    \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2]   );
  input  \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] ,
    \B[8] , \B[9] , \B[10] ;
  output \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2] ;
  wire n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
    n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
    n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
    n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
    n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n274, n275,
    n276, n277;
  assign n19 = ~\B[1]  & \B[4] ;
  assign n20 = ~\B[4]  & ~\B[8] ;
  assign n21 = ~n19 & ~n20;
  assign n22 = \B[0]  & ~n21;
  assign n23 = \B[1]  & \B[4] ;
  assign n24 = ~\B[0]  & n23;
  assign n25 = ~n22 & ~n24;
  assign n26 = ~\B[6]  & ~n25;
  assign n27 = ~\B[7]  & n26;
  assign n28 = \B[4]  & \B[8] ;
  assign n29 = ~n27 & ~n28;
  assign n30 = ~\B[5]  & ~n29;
  assign n31 = ~\B[4]  & \B[7] ;
  assign n32 = \B[1]  & ~\B[2] ;
  assign n33 = \B[5]  & ~\B[7] ;
  assign n34 = n32 & n33;
  assign n35 = ~n31 & ~n34;
  assign n36 = \B[3]  & ~n35;
  assign n37 = \B[4]  & \B[7] ;
  assign n38 = ~\B[3]  & n37;
  assign n39 = ~n36 & ~n38;
  assign n40 = ~\B[8]  & ~n39;
  assign n41 = \B[5]  & \B[8] ;
  assign n42 = ~\B[4]  & n41;
  assign n43 = ~n40 & ~n42;
  assign n44 = ~n30 & n43;
  assign n45 = ~\B[9]  & ~n44;
  assign n46 = \B[4]  & ~\B[8] ;
  assign n47 = ~\B[3]  & n46;
  assign n48 = ~\B[4]  & ~\B[7] ;
  assign n49 = ~n47 & ~n48;
  assign n50 = ~\B[2]  & ~n49;
  assign n51 = \B[1]  & n50;
  assign n52 = ~\B[1]  & \B[2] ;
  assign n53 = ~\B[7]  & ~\B[8] ;
  assign n54 = n52 & n53;
  assign n55 = ~\B[9]  & ~n54;
  assign n56 = ~n51 & n55;
  assign n57 = ~\B[6]  & ~n56;
  assign n58 = \B[5]  & n57;
  assign n59 = \B[6]  & \B[9] ;
  assign n60 = ~\B[5]  & n59;
  assign n61 = ~n58 & ~n60;
  assign n62 = ~n45 & n61;
  assign n63 = ~\B[10]  & ~n62;
  assign n64 = ~\B[2]  & \B[3] ;
  assign n65 = \B[2]  & ~\B[3] ;
  assign n66 = ~n64 & ~n65;
  assign n67 = ~\B[9]  & ~n66;
  assign n68 = ~\B[8]  & n67;
  assign n69 = ~\B[10]  & ~n68;
  assign n70 = ~\B[7]  & ~n69;
  assign n71 = \B[9]  & \B[10] ;
  assign n72 = \B[8]  & n71;
  assign n73 = ~n70 & ~n72;
  assign n74 = \B[6]  & ~n73;
  assign n75 = ~\B[6]  & \B[10] ;
  assign n76 = \B[7]  & n75;
  assign n77 = ~n74 & ~n76;
  assign \M[0]  = n63 | ~n77;
  assign n79 = ~\B[4]  & ~\B[9] ;
  assign n80 = ~\B[2]  & ~\B[7] ;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~\B[1]  & ~n81;
  assign n83 = \B[1]  & \B[2] ;
  assign n84 = \B[0]  & n83;
  assign n85 = ~\B[0]  & ~\B[2] ;
  assign n86 = ~n84 & ~n85;
  assign n87 = ~\B[7]  & ~n86;
  assign n88 = \B[4]  & n87;
  assign n89 = \B[8]  & ~\B[9] ;
  assign n90 = ~n88 & ~n89;
  assign n91 = ~n82 & n90;
  assign n92 = ~\B[6]  & ~n91;
  assign n93 = \B[3]  & \B[4] ;
  assign n94 = \B[7]  & ~n93;
  assign n95 = ~\B[9]  & n94;
  assign n96 = ~\B[8]  & n95;
  assign n97 = ~\B[7]  & \B[9] ;
  assign n98 = ~n96 & ~n97;
  assign n99 = ~n92 & n98;
  assign n100 = ~\B[5]  & ~n99;
  assign n101 = ~\B[8]  & ~\B[9] ;
  assign n102 = \B[4]  & n101;
  assign n103 = ~\B[6]  & ~\B[7] ;
  assign n104 = ~\B[4]  & n103;
  assign n105 = ~n102 & ~n104;
  assign n106 = \B[2]  & ~n105;
  assign n107 = \B[1]  & n106;
  assign n108 = \B[7]  & ~\B[9] ;
  assign n109 = n46 & n108;
  assign n110 = ~n107 & ~n109;
  assign n111 = \B[3]  & ~n110;
  assign n112 = \B[4]  & n89;
  assign n113 = \B[7]  & \B[9] ;
  assign n114 = ~n112 & ~n113;
  assign n115 = \B[6]  & ~n114;
  assign n116 = ~n111 & ~n115;
  assign n117 = \B[5]  & ~n116;
  assign n118 = ~\B[4]  & n89;
  assign n119 = ~n97 & ~n118;
  assign n120 = ~\B[6]  & ~n119;
  assign n121 = ~n117 & ~n120;
  assign n122 = ~n100 & n121;
  assign n123 = ~\B[10]  & ~n122;
  assign n124 = \B[6]  & ~\B[9] ;
  assign n125 = ~\B[4]  & n124;
  assign n126 = \B[5]  & ~\B[6] ;
  assign n127 = ~\B[3]  & n126;
  assign n128 = ~n125 & ~n127;
  assign n129 = ~\B[2]  & ~n128;
  assign n130 = ~\B[1]  & n126;
  assign n131 = ~n125 & ~n130;
  assign n132 = ~\B[3]  & ~n131;
  assign n133 = \B[2]  & \B[3] ;
  assign n134 = \B[4]  & n124;
  assign n135 = n133 & n134;
  assign n136 = ~\B[10]  & ~n135;
  assign n137 = ~n132 & n136;
  assign n138 = ~n129 & n137;
  assign n139 = ~\B[7]  & ~n138;
  assign n140 = ~n75 & ~n139;
  assign n141 = ~\B[8]  & ~n140;
  assign n142 = \B[6]  & \B[10] ;
  assign n143 = \B[7]  & n142;
  assign n144 = n89 & n143;
  assign n145 = ~n141 & ~n144;
  assign \M[1]  = ~n123 & n145;
  assign n147 = \B[4]  & ~\B[6] ;
  assign n148 = \B[0]  & ~\B[3] ;
  assign n149 = n147 & n148;
  assign n150 = ~\B[4]  & \B[5] ;
  assign n151 = \B[3]  & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = \B[1]  & ~n152;
  assign n154 = ~\B[4]  & ~\B[6] ;
  assign n155 = \B[0]  & \B[1] ;
  assign n156 = \B[4]  & ~n155;
  assign n157 = \B[3]  & n156;
  assign n158 = ~n154 & ~n157;
  assign n159 = ~\B[5]  & ~n158;
  assign n160 = ~n153 & ~n159;
  assign n161 = \B[2]  & ~n160;
  assign n162 = \B[3]  & ~\B[6] ;
  assign n163 = ~\B[2]  & n162;
  assign n164 = ~\B[3]  & \B[5] ;
  assign n165 = ~n163 & ~n164;
  assign n166 = \B[4]  & ~n165;
  assign n167 = ~n161 & ~n166;
  assign n168 = ~\B[7]  & ~n167;
  assign n169 = ~\B[5]  & \B[6] ;
  assign n170 = \B[2]  & n169;
  assign n171 = ~n130 & ~n170;
  assign n172 = \B[4]  & ~n171;
  assign n173 = \B[3]  & n172;
  assign n174 = \B[5]  & ~n93;
  assign n175 = \B[6]  & n174;
  assign n176 = ~n173 & ~n175;
  assign n177 = ~n168 & n176;
  assign n178 = ~\B[8]  & ~n177;
  assign n179 = ~\B[6]  & \B[7] ;
  assign n180 = \B[3]  & n179;
  assign n181 = \B[6]  & ~\B[7] ;
  assign n182 = ~\B[2]  & n181;
  assign n183 = ~n180 & ~n182;
  assign n184 = \B[5]  & ~n183;
  assign n185 = \B[4]  & n184;
  assign n186 = \B[4]  & \B[5] ;
  assign n187 = \B[7]  & ~n186;
  assign n188 = \B[6]  & n187;
  assign n189 = ~n185 & ~n188;
  assign n190 = ~n178 & n189;
  assign n191 = ~\B[9]  & ~n190;
  assign n192 = \B[4]  & \B[6] ;
  assign n193 = n33 & n192;
  assign n194 = ~n179 & ~n193;
  assign n195 = \B[8]  & ~n194;
  assign n196 = ~n191 & ~n195;
  assign n197 = ~\B[10]  & ~n196;
  assign n198 = \B[8]  & \B[10] ;
  assign n199 = ~\B[8]  & \B[9] ;
  assign n200 = \B[5]  & n199;
  assign n201 = ~n198 & ~n200;
  assign n202 = \B[7]  & ~n201;
  assign n203 = \B[6]  & n202;
  assign n204 = \B[5]  & \B[7] ;
  assign n205 = \B[8]  & ~n204;
  assign n206 = ~\B[10]  & ~n205;
  assign n207 = \B[9]  & ~n206;
  assign n208 = ~n203 & ~n207;
  assign \M[2]  = n197 | ~n208;
  assign n210 = \B[6]  & \B[7] ;
  assign n211 = ~\B[2]  & n210;
  assign n212 = \B[5]  & n28;
  assign n213 = n211 & n212;
  assign n214 = ~\B[5]  & n20;
  assign n215 = n103 & n214;
  assign n216 = ~n213 & ~n215;
  assign n217 = ~\B[9]  & ~n216;
  assign n218 = ~\B[10]  & n217;
  assign \M[3]  = \B[3]  | ~n218;
  assign n220 = \B[5]  & \B[6] ;
  assign n221 = \B[4]  & ~\B[7] ;
  assign n222 = n220 & n221;
  assign n223 = ~\B[5]  & ~\B[6] ;
  assign n224 = n155 & n223;
  assign n225 = ~n222 & ~n224;
  assign n226 = \B[3]  & ~n225;
  assign n227 = \B[2]  & n226;
  assign n228 = ~\B[4]  & ~n181;
  assign n229 = ~\B[7]  & ~n126;
  assign n230 = ~\B[3]  & ~n229;
  assign n231 = \B[7]  & ~n220;
  assign n232 = ~\B[6]  & ~n83;
  assign n233 = \B[5]  & n232;
  assign n234 = ~\B[9]  & ~n233;
  assign n235 = ~n231 & n234;
  assign n236 = ~n230 & n235;
  assign n237 = ~n228 & n236;
  assign n238 = ~n227 & n237;
  assign n239 = ~\B[8]  & ~n238;
  assign n240 = \B[3]  & \B[8] ;
  assign n241 = ~n65 & ~n240;
  assign n242 = \B[6]  & ~n241;
  assign n243 = \B[5]  & n242;
  assign n244 = \B[7]  & n243;
  assign n245 = ~\B[9]  & n244;
  assign n246 = \B[4]  & n245;
  assign n247 = \B[7]  & n220;
  assign n248 = \B[9]  & ~n247;
  assign n249 = ~n246 & ~n248;
  assign n250 = ~n239 & n249;
  assign \E[0]  = \B[10]  | n250;
  assign n252 = \B[6]  & \B[8] ;
  assign n253 = n204 & n252;
  assign n254 = \B[1]  & \B[3] ;
  assign n255 = \B[0]  & n254;
  assign n256 = ~\B[5]  & ~\B[7] ;
  assign n257 = ~\B[8]  & n256;
  assign n258 = n255 & n257;
  assign n259 = ~n253 & ~n258;
  assign n260 = \B[2]  & ~n259;
  assign n261 = \B[8]  & n204;
  assign n262 = \B[3]  & \B[6] ;
  assign n263 = n261 & n262;
  assign n264 = ~n260 & ~n263;
  assign n265 = \B[4]  & ~n264;
  assign n266 = n133 & n192;
  assign n267 = \B[5]  & ~n266;
  assign n268 = ~n169 & ~n267;
  assign n269 = ~\B[7]  & ~n268;
  assign n270 = ~\B[8]  & n269;
  assign n271 = ~\B[9]  & ~\B[10] ;
  assign n272 = ~n270 & n271;
  assign \E[1]  = n265 | ~n272;
  assign n274 = \B[2]  & n93;
  assign n275 = n220 & n274;
  assign n276 = ~\B[9]  & ~n275;
  assign n277 = ~\B[10]  & n276;
  assign \E[2]  = ~n53 | ~n277;
endmodule

