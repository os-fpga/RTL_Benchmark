--------------------------------------------------------------------------------
--                                                                            --
--                          V H D L    F I L E                                --
--                          COPYRIGHT (C) 2006                                --
--                                                                            --
--------------------------------------------------------------------------------
--
-- Title       : CLKGEN
-- Design      : MDCT Core
-- Author      : Michal Krepa
--
--------------------------------------------------------------------------------
--
-- File        : CLKGEN.VHD
-- Created     : Sat Mar 12 2006
--
--------------------------------------------------------------------------------
--
--  Description : Clock generator for simulation
--
--------------------------------------------------------------------------------
library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all; 

library WORK;
  use WORK.MDCT_PKG.all;
  
entity CLKGEN is
  port (   
        clk               : out STD_LOGIC
       );
end CLKGEN;

--**************************************************************************--

architecture SIM of CLKGEN is	 

  signal clk_s            : STD_LOGIC;	 

begin

  ----------------------------------------------------------------------------
  clk_gen_proc:	-- clock generator
  ----------------------------------------------------------------------------
  process
    constant PERIOD       : TIME := 1 us /(CLK_FREQ_C);
  begin
    clk_s                 <= '0';
    wait for PERIOD/2;
    clk_s                 <= '1';
    wait for PERIOD/2;
  end process;

  ----------------------------------------------------------------------------
  clk_drv:
  ----------------------------------------------------------------------------
  clk                     <= clk_s;

end SIM;
--**************************************************************************--