library ieee;
use ieee.std_logic_1164.all;

entity top is
	port( priority, req: in std_logic_vector(127 downto 0);
	grant: out std_logic_vector(127 downto 0);
	anyGrant: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838: std_logic;

begin

w0 <= priority(1) and not req(1);
w1 <= not priority(2) and not w0;
w2 <= not req(2) and not req(3);
w3 <= not w1 and w2;
w4 <= priority(3) and not req(3);
w5 <= not priority(4) and not w4;
w6 <= not priority(5) and w5;
w7 <= not w3 and w6;
w8 <= not priority(5) and req(4);
w9 <= not req(5) and not req(6);
w10 <= not w8 and w9;
w11 <= not w7 and w10;
w12 <= priority(6) and not req(6);
w13 <= not priority(7) and not w12;
w14 <= not priority(8) and w13;
w15 <= not w11 and w14;
w16 <= not priority(8) and req(7);
w17 <= not req(8) and not req(9);
w18 <= not w16 and w17;
w19 <= not w15 and w18;
w20 <= priority(9) and not req(9);
w21 <= not priority(10) and not w20;
w22 <= not priority(11) and w21;
w23 <= not w19 and w22;
w24 <= not priority(11) and req(10);
w25 <= not req(11) and not req(12);
w26 <= not w24 and w25;
w27 <= not w23 and w26;
w28 <= priority(12) and not req(12);
w29 <= not priority(13) and not w28;
w30 <= not priority(14) and w29;
w31 <= not w27 and w30;
w32 <= not priority(14) and req(13);
w33 <= not req(14) and not req(15);
w34 <= not w32 and w33;
w35 <= not w31 and w34;
w36 <= priority(15) and not req(15);
w37 <= not priority(16) and not w36;
w38 <= not priority(17) and w37;
w39 <= not w35 and w38;
w40 <= not priority(17) and req(16);
w41 <= not req(17) and not req(18);
w42 <= not w40 and w41;
w43 <= not w39 and w42;
w44 <= priority(18) and not req(18);
w45 <= not priority(19) and not w44;
w46 <= not priority(20) and w45;
w47 <= not w43 and w46;
w48 <= not priority(20) and req(19);
w49 <= not req(20) and not req(21);
w50 <= not w48 and w49;
w51 <= not w47 and w50;
w52 <= priority(21) and not req(21);
w53 <= not priority(22) and not w52;
w54 <= not priority(23) and w53;
w55 <= not w51 and w54;
w56 <= not priority(23) and req(22);
w57 <= not req(23) and not req(24);
w58 <= not w56 and w57;
w59 <= not w55 and w58;
w60 <= priority(24) and not req(24);
w61 <= not priority(25) and not w60;
w62 <= not priority(26) and w61;
w63 <= not w59 and w62;
w64 <= not priority(26) and req(25);
w65 <= not req(26) and not req(27);
w66 <= not w64 and w65;
w67 <= not w63 and w66;
w68 <= priority(27) and not req(27);
w69 <= not priority(28) and not w68;
w70 <= not priority(29) and w69;
w71 <= not w67 and w70;
w72 <= not priority(29) and req(28);
w73 <= not req(29) and not req(30);
w74 <= not w72 and w73;
w75 <= not w71 and w74;
w76 <= priority(30) and not req(30);
w77 <= not priority(31) and not w76;
w78 <= not priority(32) and w77;
w79 <= not w75 and w78;
w80 <= not priority(32) and req(31);
w81 <= not req(32) and not req(33);
w82 <= not w80 and w81;
w83 <= not w79 and w82;
w84 <= priority(33) and not req(33);
w85 <= not priority(34) and not w84;
w86 <= not priority(35) and w85;
w87 <= not w83 and w86;
w88 <= not priority(35) and req(34);
w89 <= not req(35) and not req(36);
w90 <= not w88 and w89;
w91 <= not w87 and w90;
w92 <= priority(36) and not req(36);
w93 <= not priority(37) and not w92;
w94 <= not priority(38) and w93;
w95 <= not w91 and w94;
w96 <= not priority(38) and req(37);
w97 <= not req(38) and not req(39);
w98 <= not w96 and w97;
w99 <= not w95 and w98;
w100 <= priority(39) and not req(39);
w101 <= not priority(40) and not w100;
w102 <= not priority(41) and w101;
w103 <= not w99 and w102;
w104 <= not priority(41) and req(40);
w105 <= not req(41) and not req(42);
w106 <= not w104 and w105;
w107 <= not w103 and w106;
w108 <= priority(42) and not req(42);
w109 <= not priority(43) and not w108;
w110 <= not priority(44) and w109;
w111 <= not w107 and w110;
w112 <= not priority(44) and req(43);
w113 <= not req(44) and not req(45);
w114 <= not w112 and w113;
w115 <= not w111 and w114;
w116 <= priority(45) and not req(45);
w117 <= not priority(46) and not w116;
w118 <= not priority(47) and w117;
w119 <= not w115 and w118;
w120 <= not priority(47) and req(46);
w121 <= not req(47) and not req(48);
w122 <= not w120 and w121;
w123 <= not w119 and w122;
w124 <= priority(48) and not req(48);
w125 <= not priority(49) and not w124;
w126 <= not priority(50) and w125;
w127 <= not w123 and w126;
w128 <= not priority(50) and req(49);
w129 <= not req(50) and not req(51);
w130 <= not w128 and w129;
w131 <= not w127 and w130;
w132 <= priority(51) and not req(51);
w133 <= not priority(52) and not w132;
w134 <= not priority(53) and w133;
w135 <= not w131 and w134;
w136 <= not priority(53) and req(52);
w137 <= not req(53) and not req(54);
w138 <= not w136 and w137;
w139 <= not w135 and w138;
w140 <= priority(54) and not req(54);
w141 <= not priority(55) and not w140;
w142 <= not priority(56) and w141;
w143 <= not w139 and w142;
w144 <= not priority(56) and req(55);
w145 <= not req(56) and not req(57);
w146 <= not w144 and w145;
w147 <= not w143 and w146;
w148 <= priority(57) and not req(57);
w149 <= not priority(58) and not w148;
w150 <= not priority(59) and w149;
w151 <= not w147 and w150;
w152 <= not priority(59) and req(58);
w153 <= not req(59) and not req(60);
w154 <= not w152 and w153;
w155 <= not w151 and w154;
w156 <= priority(60) and not req(60);
w157 <= not priority(61) and not w156;
w158 <= not priority(62) and w157;
w159 <= not w155 and w158;
w160 <= not priority(62) and req(61);
w161 <= not req(62) and not req(63);
w162 <= not w160 and w161;
w163 <= not w159 and w162;
w164 <= priority(63) and not req(63);
w165 <= not priority(64) and not w164;
w166 <= not priority(65) and w165;
w167 <= not w163 and w166;
w168 <= not priority(65) and req(64);
w169 <= not req(65) and not req(66);
w170 <= not w168 and w169;
w171 <= not w167 and w170;
w172 <= priority(66) and not req(66);
w173 <= not priority(67) and not w172;
w174 <= not priority(68) and w173;
w175 <= not w171 and w174;
w176 <= not priority(68) and req(67);
w177 <= not req(68) and not req(69);
w178 <= not w176 and w177;
w179 <= not w175 and w178;
w180 <= priority(69) and not req(69);
w181 <= not priority(70) and not w180;
w182 <= not priority(71) and w181;
w183 <= not w179 and w182;
w184 <= not priority(71) and req(70);
w185 <= not req(71) and not req(72);
w186 <= not w184 and w185;
w187 <= not w183 and w186;
w188 <= priority(72) and not req(72);
w189 <= not priority(73) and not w188;
w190 <= not priority(74) and w189;
w191 <= not w187 and w190;
w192 <= not priority(74) and req(73);
w193 <= not req(74) and not req(75);
w194 <= not w192 and w193;
w195 <= not w191 and w194;
w196 <= priority(75) and not req(75);
w197 <= not priority(76) and not w196;
w198 <= not priority(77) and w197;
w199 <= not w195 and w198;
w200 <= not priority(77) and req(76);
w201 <= not req(77) and not req(78);
w202 <= not w200 and w201;
w203 <= not w199 and w202;
w204 <= priority(78) and not req(78);
w205 <= not priority(79) and not w204;
w206 <= not priority(80) and w205;
w207 <= not w203 and w206;
w208 <= not priority(80) and req(79);
w209 <= not req(80) and not req(81);
w210 <= not w208 and w209;
w211 <= not w207 and w210;
w212 <= priority(81) and not req(81);
w213 <= not priority(82) and not w212;
w214 <= not priority(83) and w213;
w215 <= not w211 and w214;
w216 <= not priority(83) and req(82);
w217 <= not req(83) and not req(84);
w218 <= not w216 and w217;
w219 <= not w215 and w218;
w220 <= priority(84) and not req(84);
w221 <= not priority(85) and not w220;
w222 <= not priority(86) and w221;
w223 <= not w219 and w222;
w224 <= not priority(86) and req(85);
w225 <= not req(86) and not req(87);
w226 <= not w224 and w225;
w227 <= not w223 and w226;
w228 <= priority(87) and not req(87);
w229 <= not priority(88) and not w228;
w230 <= not priority(89) and w229;
w231 <= not w227 and w230;
w232 <= not priority(89) and req(88);
w233 <= not req(89) and not req(90);
w234 <= not w232 and w233;
w235 <= not w231 and w234;
w236 <= priority(90) and not req(90);
w237 <= not priority(91) and not w236;
w238 <= not priority(92) and w237;
w239 <= not w235 and w238;
w240 <= not priority(92) and req(91);
w241 <= not req(92) and not req(93);
w242 <= not w240 and w241;
w243 <= not w239 and w242;
w244 <= priority(93) and not req(93);
w245 <= not priority(94) and not w244;
w246 <= not priority(95) and w245;
w247 <= not w243 and w246;
w248 <= not priority(95) and req(94);
w249 <= not req(95) and not req(96);
w250 <= not w248 and w249;
w251 <= not w247 and w250;
w252 <= priority(96) and not req(96);
w253 <= not priority(97) and not w252;
w254 <= not priority(98) and w253;
w255 <= not w251 and w254;
w256 <= not priority(98) and req(97);
w257 <= not req(98) and not req(99);
w258 <= not w256 and w257;
w259 <= not w255 and w258;
w260 <= priority(99) and not req(99);
w261 <= not priority(100) and not w260;
w262 <= not priority(101) and w261;
w263 <= not w259 and w262;
w264 <= not priority(101) and req(100);
w265 <= not req(101) and not req(102);
w266 <= not w264 and w265;
w267 <= not w263 and w266;
w268 <= priority(102) and not req(102);
w269 <= not priority(103) and not w268;
w270 <= not priority(104) and w269;
w271 <= not w267 and w270;
w272 <= not priority(104) and req(103);
w273 <= not req(104) and not req(105);
w274 <= not w272 and w273;
w275 <= not w271 and w274;
w276 <= priority(105) and not req(105);
w277 <= not priority(106) and not w276;
w278 <= not priority(107) and w277;
w279 <= not w275 and w278;
w280 <= not priority(107) and req(106);
w281 <= not req(107) and not req(108);
w282 <= not w280 and w281;
w283 <= not w279 and w282;
w284 <= priority(108) and not req(108);
w285 <= not priority(109) and not w284;
w286 <= not priority(110) and w285;
w287 <= not w283 and w286;
w288 <= not priority(110) and req(109);
w289 <= not req(110) and not req(111);
w290 <= not w288 and w289;
w291 <= not w287 and w290;
w292 <= priority(111) and not req(111);
w293 <= not priority(112) and not w292;
w294 <= not priority(113) and w293;
w295 <= not w291 and w294;
w296 <= not priority(113) and req(112);
w297 <= not req(113) and not req(114);
w298 <= not w296 and w297;
w299 <= not w295 and w298;
w300 <= priority(114) and not req(114);
w301 <= not priority(115) and not w300;
w302 <= not priority(116) and w301;
w303 <= not w299 and w302;
w304 <= not priority(116) and req(115);
w305 <= not req(116) and not req(117);
w306 <= not w304 and w305;
w307 <= not w303 and w306;
w308 <= priority(117) and not req(117);
w309 <= not priority(118) and not w308;
w310 <= not priority(119) and w309;
w311 <= not w307 and w310;
w312 <= not priority(119) and req(118);
w313 <= not req(119) and not req(120);
w314 <= not w312 and w313;
w315 <= not w311 and w314;
w316 <= priority(120) and not req(120);
w317 <= not priority(121) and not w316;
w318 <= not priority(122) and w317;
w319 <= not w315 and w318;
w320 <= not priority(122) and req(121);
w321 <= not req(122) and not req(123);
w322 <= not w320 and w321;
w323 <= not w319 and w322;
w324 <= priority(123) and not req(123);
w325 <= not priority(124) and not w324;
w326 <= not priority(125) and w325;
w327 <= not w323 and w326;
w328 <= not priority(125) and req(124);
w329 <= not req(125) and not req(126);
w330 <= not w328 and w329;
w331 <= not w327 and w330;
w332 <= priority(126) and not req(126);
w333 <= not priority(127) and not w332;
w334 <= not priority(0) and w333;
w335 <= not w331 and w334;
w336 <= not priority(0) and req(127);
w337 <= req(0) and not w336;
w338 <= not w335 and w337;
w339 <= priority(2) and not req(2);
w340 <= not priority(3) and not w339;
w341 <= not req(3) and not req(4);
w342 <= not w340 and w341;
w343 <= priority(4) and not req(4);
w344 <= not priority(5) and not w343;
w345 <= not priority(6) and w344;
w346 <= not w342 and w345;
w347 <= not priority(6) and req(5);
w348 <= not req(6) and not req(7);
w349 <= not w347 and w348;
w350 <= not w346 and w349;
w351 <= priority(7) and not req(7);
w352 <= not priority(8) and not w351;
w353 <= not priority(9) and w352;
w354 <= not w350 and w353;
w355 <= not priority(9) and req(8);
w356 <= not req(9) and not req(10);
w357 <= not w355 and w356;
w358 <= not w354 and w357;
w359 <= priority(10) and not req(10);
w360 <= not priority(11) and not w359;
w361 <= not priority(12) and w360;
w362 <= not w358 and w361;
w363 <= not priority(12) and req(11);
w364 <= not req(12) and not req(13);
w365 <= not w363 and w364;
w366 <= not w362 and w365;
w367 <= priority(13) and not req(13);
w368 <= not priority(14) and not w367;
w369 <= not priority(15) and w368;
w370 <= not w366 and w369;
w371 <= not priority(15) and req(14);
w372 <= not req(15) and not req(16);
w373 <= not w371 and w372;
w374 <= not w370 and w373;
w375 <= priority(16) and not req(16);
w376 <= not priority(17) and not w375;
w377 <= not priority(18) and w376;
w378 <= not w374 and w377;
w379 <= not priority(18) and req(17);
w380 <= not req(18) and not req(19);
w381 <= not w379 and w380;
w382 <= not w378 and w381;
w383 <= priority(19) and not req(19);
w384 <= not priority(20) and not w383;
w385 <= not priority(21) and w384;
w386 <= not w382 and w385;
w387 <= not priority(21) and req(20);
w388 <= not req(21) and not req(22);
w389 <= not w387 and w388;
w390 <= not w386 and w389;
w391 <= priority(22) and not req(22);
w392 <= not priority(23) and not w391;
w393 <= not priority(24) and w392;
w394 <= not w390 and w393;
w395 <= not priority(24) and req(23);
w396 <= not req(24) and not req(25);
w397 <= not w395 and w396;
w398 <= not w394 and w397;
w399 <= priority(25) and not req(25);
w400 <= not priority(26) and not w399;
w401 <= not priority(27) and w400;
w402 <= not w398 and w401;
w403 <= not priority(27) and req(26);
w404 <= not req(27) and not req(28);
w405 <= not w403 and w404;
w406 <= not w402 and w405;
w407 <= priority(28) and not req(28);
w408 <= not priority(29) and not w407;
w409 <= not priority(30) and w408;
w410 <= not w406 and w409;
w411 <= not priority(30) and req(29);
w412 <= not req(30) and not req(31);
w413 <= not w411 and w412;
w414 <= not w410 and w413;
w415 <= priority(31) and not req(31);
w416 <= not priority(32) and not w415;
w417 <= not priority(33) and w416;
w418 <= not w414 and w417;
w419 <= not priority(33) and req(32);
w420 <= not req(33) and not req(34);
w421 <= not w419 and w420;
w422 <= not w418 and w421;
w423 <= priority(34) and not req(34);
w424 <= not priority(35) and not w423;
w425 <= not priority(36) and w424;
w426 <= not w422 and w425;
w427 <= not priority(36) and req(35);
w428 <= not req(36) and not req(37);
w429 <= not w427 and w428;
w430 <= not w426 and w429;
w431 <= priority(37) and not req(37);
w432 <= not priority(38) and not w431;
w433 <= not priority(39) and w432;
w434 <= not w430 and w433;
w435 <= not priority(39) and req(38);
w436 <= not req(39) and not req(40);
w437 <= not w435 and w436;
w438 <= not w434 and w437;
w439 <= priority(40) and not req(40);
w440 <= not priority(41) and not w439;
w441 <= not priority(42) and w440;
w442 <= not w438 and w441;
w443 <= not priority(42) and req(41);
w444 <= not req(42) and not req(43);
w445 <= not w443 and w444;
w446 <= not w442 and w445;
w447 <= priority(43) and not req(43);
w448 <= not priority(44) and not w447;
w449 <= not priority(45) and w448;
w450 <= not w446 and w449;
w451 <= not priority(45) and req(44);
w452 <= not req(45) and not req(46);
w453 <= not w451 and w452;
w454 <= not w450 and w453;
w455 <= priority(46) and not req(46);
w456 <= not priority(47) and not w455;
w457 <= not priority(48) and w456;
w458 <= not w454 and w457;
w459 <= not priority(48) and req(47);
w460 <= not req(48) and not req(49);
w461 <= not w459 and w460;
w462 <= not w458 and w461;
w463 <= priority(49) and not req(49);
w464 <= not priority(50) and not w463;
w465 <= not priority(51) and w464;
w466 <= not w462 and w465;
w467 <= not priority(51) and req(50);
w468 <= not req(51) and not req(52);
w469 <= not w467 and w468;
w470 <= not w466 and w469;
w471 <= priority(52) and not req(52);
w472 <= not priority(53) and not w471;
w473 <= not priority(54) and w472;
w474 <= not w470 and w473;
w475 <= not priority(54) and req(53);
w476 <= not req(54) and not req(55);
w477 <= not w475 and w476;
w478 <= not w474 and w477;
w479 <= priority(55) and not req(55);
w480 <= not priority(56) and not w479;
w481 <= not priority(57) and w480;
w482 <= not w478 and w481;
w483 <= not priority(57) and req(56);
w484 <= not req(57) and not req(58);
w485 <= not w483 and w484;
w486 <= not w482 and w485;
w487 <= priority(58) and not req(58);
w488 <= not priority(59) and not w487;
w489 <= not priority(60) and w488;
w490 <= not w486 and w489;
w491 <= not priority(60) and req(59);
w492 <= not req(60) and not req(61);
w493 <= not w491 and w492;
w494 <= not w490 and w493;
w495 <= priority(61) and not req(61);
w496 <= not priority(62) and not w495;
w497 <= not priority(63) and w496;
w498 <= not w494 and w497;
w499 <= not priority(63) and req(62);
w500 <= not req(63) and not req(64);
w501 <= not w499 and w500;
w502 <= not w498 and w501;
w503 <= priority(64) and not req(64);
w504 <= not priority(65) and not w503;
w505 <= not priority(66) and w504;
w506 <= not w502 and w505;
w507 <= not priority(66) and req(65);
w508 <= not req(66) and not req(67);
w509 <= not w507 and w508;
w510 <= not w506 and w509;
w511 <= priority(67) and not req(67);
w512 <= not priority(68) and not w511;
w513 <= not priority(69) and w512;
w514 <= not w510 and w513;
w515 <= not priority(69) and req(68);
w516 <= not req(69) and not req(70);
w517 <= not w515 and w516;
w518 <= not w514 and w517;
w519 <= priority(70) and not req(70);
w520 <= not priority(71) and not w519;
w521 <= not priority(72) and w520;
w522 <= not w518 and w521;
w523 <= not priority(72) and req(71);
w524 <= not req(72) and not req(73);
w525 <= not w523 and w524;
w526 <= not w522 and w525;
w527 <= priority(73) and not req(73);
w528 <= not priority(74) and not w527;
w529 <= not priority(75) and w528;
w530 <= not w526 and w529;
w531 <= not priority(75) and req(74);
w532 <= not req(75) and not req(76);
w533 <= not w531 and w532;
w534 <= not w530 and w533;
w535 <= priority(76) and not req(76);
w536 <= not priority(77) and not w535;
w537 <= not priority(78) and w536;
w538 <= not w534 and w537;
w539 <= not priority(78) and req(77);
w540 <= not req(78) and not req(79);
w541 <= not w539 and w540;
w542 <= not w538 and w541;
w543 <= priority(79) and not req(79);
w544 <= not priority(80) and not w543;
w545 <= not priority(81) and w544;
w546 <= not w542 and w545;
w547 <= not priority(81) and req(80);
w548 <= not req(81) and not req(82);
w549 <= not w547 and w548;
w550 <= not w546 and w549;
w551 <= priority(82) and not req(82);
w552 <= not priority(83) and not w551;
w553 <= not priority(84) and w552;
w554 <= not w550 and w553;
w555 <= not priority(84) and req(83);
w556 <= not req(84) and not req(85);
w557 <= not w555 and w556;
w558 <= not w554 and w557;
w559 <= priority(85) and not req(85);
w560 <= not priority(86) and not w559;
w561 <= not priority(87) and w560;
w562 <= not w558 and w561;
w563 <= not priority(87) and req(86);
w564 <= not req(87) and not req(88);
w565 <= not w563 and w564;
w566 <= not w562 and w565;
w567 <= priority(88) and not req(88);
w568 <= not priority(89) and not w567;
w569 <= not priority(90) and w568;
w570 <= not w566 and w569;
w571 <= not priority(90) and req(89);
w572 <= not req(90) and not req(91);
w573 <= not w571 and w572;
w574 <= not w570 and w573;
w575 <= priority(91) and not req(91);
w576 <= not priority(92) and not w575;
w577 <= not priority(93) and w576;
w578 <= not w574 and w577;
w579 <= not priority(93) and req(92);
w580 <= not req(93) and not req(94);
w581 <= not w579 and w580;
w582 <= not w578 and w581;
w583 <= priority(94) and not req(94);
w584 <= not priority(95) and not w583;
w585 <= not priority(96) and w584;
w586 <= not w582 and w585;
w587 <= not priority(96) and req(95);
w588 <= not req(96) and not req(97);
w589 <= not w587 and w588;
w590 <= not w586 and w589;
w591 <= priority(97) and not req(97);
w592 <= not priority(98) and not w591;
w593 <= not priority(99) and w592;
w594 <= not w590 and w593;
w595 <= not priority(99) and req(98);
w596 <= not req(99) and not req(100);
w597 <= not w595 and w596;
w598 <= not w594 and w597;
w599 <= priority(100) and not req(100);
w600 <= not priority(101) and not w599;
w601 <= not priority(102) and w600;
w602 <= not w598 and w601;
w603 <= not priority(102) and req(101);
w604 <= not req(102) and not req(103);
w605 <= not w603 and w604;
w606 <= not w602 and w605;
w607 <= priority(103) and not req(103);
w608 <= not priority(104) and not w607;
w609 <= not priority(105) and w608;
w610 <= not w606 and w609;
w611 <= not priority(105) and req(104);
w612 <= not req(105) and not req(106);
w613 <= not w611 and w612;
w614 <= not w610 and w613;
w615 <= priority(106) and not req(106);
w616 <= not priority(107) and not w615;
w617 <= not priority(108) and w616;
w618 <= not w614 and w617;
w619 <= not priority(108) and req(107);
w620 <= not req(108) and not req(109);
w621 <= not w619 and w620;
w622 <= not w618 and w621;
w623 <= priority(109) and not req(109);
w624 <= not priority(110) and not w623;
w625 <= not priority(111) and w624;
w626 <= not w622 and w625;
w627 <= not priority(111) and req(110);
w628 <= not req(111) and not req(112);
w629 <= not w627 and w628;
w630 <= not w626 and w629;
w631 <= priority(112) and not req(112);
w632 <= not priority(113) and not w631;
w633 <= not priority(114) and w632;
w634 <= not w630 and w633;
w635 <= not priority(114) and req(113);
w636 <= not req(114) and not req(115);
w637 <= not w635 and w636;
w638 <= not w634 and w637;
w639 <= priority(115) and not req(115);
w640 <= not priority(116) and not w639;
w641 <= not priority(117) and w640;
w642 <= not w638 and w641;
w643 <= not priority(117) and req(116);
w644 <= not req(117) and not req(118);
w645 <= not w643 and w644;
w646 <= not w642 and w645;
w647 <= priority(118) and not req(118);
w648 <= not priority(119) and not w647;
w649 <= not priority(120) and w648;
w650 <= not w646 and w649;
w651 <= not priority(120) and req(119);
w652 <= not req(120) and not req(121);
w653 <= not w651 and w652;
w654 <= not w650 and w653;
w655 <= priority(121) and not req(121);
w656 <= not priority(122) and not w655;
w657 <= not priority(123) and w656;
w658 <= not w654 and w657;
w659 <= not priority(123) and req(122);
w660 <= not req(123) and not req(124);
w661 <= not w659 and w660;
w662 <= not w658 and w661;
w663 <= priority(124) and not req(124);
w664 <= not priority(125) and not w663;
w665 <= not priority(126) and w664;
w666 <= not w662 and w665;
w667 <= not priority(126) and req(125);
w668 <= not req(126) and not req(127);
w669 <= not w667 and w668;
w670 <= not w666 and w669;
w671 <= priority(127) and not req(127);
w672 <= not priority(0) and not w671;
w673 <= not priority(1) and w672;
w674 <= not w670 and w673;
w675 <= not priority(1) and req(0);
w676 <= req(1) and not w675;
w677 <= not w674 and w676;
w678 <= not req(4) and not req(5);
w679 <= not w5 and w678;
w680 <= priority(5) and not req(5);
w681 <= not priority(6) and not w680;
w682 <= not priority(7) and w681;
w683 <= not w679 and w682;
w684 <= not priority(7) and req(6);
w685 <= not req(7) and not req(8);
w686 <= not w684 and w685;
w687 <= not w683 and w686;
w688 <= priority(8) and not req(8);
w689 <= not priority(9) and not w688;
w690 <= not priority(10) and w689;
w691 <= not w687 and w690;
w692 <= not priority(10) and req(9);
w693 <= not req(10) and not req(11);
w694 <= not w692 and w693;
w695 <= not w691 and w694;
w696 <= priority(11) and not req(11);
w697 <= not priority(12) and not w696;
w698 <= not priority(13) and w697;
w699 <= not w695 and w698;
w700 <= not priority(13) and req(12);
w701 <= not req(13) and not req(14);
w702 <= not w700 and w701;
w703 <= not w699 and w702;
w704 <= priority(14) and not req(14);
w705 <= not priority(15) and not w704;
w706 <= not priority(16) and w705;
w707 <= not w703 and w706;
w708 <= not priority(16) and req(15);
w709 <= not req(16) and not req(17);
w710 <= not w708 and w709;
w711 <= not w707 and w710;
w712 <= priority(17) and not req(17);
w713 <= not priority(18) and not w712;
w714 <= not priority(19) and w713;
w715 <= not w711 and w714;
w716 <= not priority(19) and req(18);
w717 <= not req(19) and not req(20);
w718 <= not w716 and w717;
w719 <= not w715 and w718;
w720 <= priority(20) and not req(20);
w721 <= not priority(21) and not w720;
w722 <= not priority(22) and w721;
w723 <= not w719 and w722;
w724 <= not priority(22) and req(21);
w725 <= not req(22) and not req(23);
w726 <= not w724 and w725;
w727 <= not w723 and w726;
w728 <= priority(23) and not req(23);
w729 <= not priority(24) and not w728;
w730 <= not priority(25) and w729;
w731 <= not w727 and w730;
w732 <= not priority(25) and req(24);
w733 <= not req(25) and not req(26);
w734 <= not w732 and w733;
w735 <= not w731 and w734;
w736 <= priority(26) and not req(26);
w737 <= not priority(27) and not w736;
w738 <= not priority(28) and w737;
w739 <= not w735 and w738;
w740 <= not priority(28) and req(27);
w741 <= not req(28) and not req(29);
w742 <= not w740 and w741;
w743 <= not w739 and w742;
w744 <= priority(29) and not req(29);
w745 <= not priority(30) and not w744;
w746 <= not priority(31) and w745;
w747 <= not w743 and w746;
w748 <= not priority(31) and req(30);
w749 <= not req(31) and not req(32);
w750 <= not w748 and w749;
w751 <= not w747 and w750;
w752 <= priority(32) and not req(32);
w753 <= not priority(33) and not w752;
w754 <= not priority(34) and w753;
w755 <= not w751 and w754;
w756 <= not priority(34) and req(33);
w757 <= not req(34) and not req(35);
w758 <= not w756 and w757;
w759 <= not w755 and w758;
w760 <= priority(35) and not req(35);
w761 <= not priority(36) and not w760;
w762 <= not priority(37) and w761;
w763 <= not w759 and w762;
w764 <= not priority(37) and req(36);
w765 <= not req(37) and not req(38);
w766 <= not w764 and w765;
w767 <= not w763 and w766;
w768 <= priority(38) and not req(38);
w769 <= not priority(39) and not w768;
w770 <= not priority(40) and w769;
w771 <= not w767 and w770;
w772 <= not priority(40) and req(39);
w773 <= not req(40) and not req(41);
w774 <= not w772 and w773;
w775 <= not w771 and w774;
w776 <= priority(41) and not req(41);
w777 <= not priority(42) and not w776;
w778 <= not priority(43) and w777;
w779 <= not w775 and w778;
w780 <= not priority(43) and req(42);
w781 <= not req(43) and not req(44);
w782 <= not w780 and w781;
w783 <= not w779 and w782;
w784 <= priority(44) and not req(44);
w785 <= not priority(45) and not w784;
w786 <= not priority(46) and w785;
w787 <= not w783 and w786;
w788 <= not priority(46) and req(45);
w789 <= not req(46) and not req(47);
w790 <= not w788 and w789;
w791 <= not w787 and w790;
w792 <= priority(47) and not req(47);
w793 <= not priority(48) and not w792;
w794 <= not priority(49) and w793;
w795 <= not w791 and w794;
w796 <= not priority(49) and req(48);
w797 <= not req(49) and not req(50);
w798 <= not w796 and w797;
w799 <= not w795 and w798;
w800 <= priority(50) and not req(50);
w801 <= not priority(51) and not w800;
w802 <= not priority(52) and w801;
w803 <= not w799 and w802;
w804 <= not priority(52) and req(51);
w805 <= not req(52) and not req(53);
w806 <= not w804 and w805;
w807 <= not w803 and w806;
w808 <= priority(53) and not req(53);
w809 <= not priority(54) and not w808;
w810 <= not priority(55) and w809;
w811 <= not w807 and w810;
w812 <= not priority(55) and req(54);
w813 <= not req(55) and not req(56);
w814 <= not w812 and w813;
w815 <= not w811 and w814;
w816 <= priority(56) and not req(56);
w817 <= not priority(57) and not w816;
w818 <= not priority(58) and w817;
w819 <= not w815 and w818;
w820 <= not priority(58) and req(57);
w821 <= not req(58) and not req(59);
w822 <= not w820 and w821;
w823 <= not w819 and w822;
w824 <= priority(59) and not req(59);
w825 <= not priority(60) and not w824;
w826 <= not priority(61) and w825;
w827 <= not w823 and w826;
w828 <= not priority(61) and req(60);
w829 <= not req(61) and not req(62);
w830 <= not w828 and w829;
w831 <= not w827 and w830;
w832 <= priority(62) and not req(62);
w833 <= not priority(63) and not w832;
w834 <= not priority(64) and w833;
w835 <= not w831 and w834;
w836 <= not priority(64) and req(63);
w837 <= not req(64) and not req(65);
w838 <= not w836 and w837;
w839 <= not w835 and w838;
w840 <= priority(65) and not req(65);
w841 <= not priority(66) and not w840;
w842 <= not priority(67) and w841;
w843 <= not w839 and w842;
w844 <= not priority(67) and req(66);
w845 <= not req(67) and not req(68);
w846 <= not w844 and w845;
w847 <= not w843 and w846;
w848 <= priority(68) and not req(68);
w849 <= not priority(69) and not w848;
w850 <= not priority(70) and w849;
w851 <= not w847 and w850;
w852 <= not priority(70) and req(69);
w853 <= not req(70) and not req(71);
w854 <= not w852 and w853;
w855 <= not w851 and w854;
w856 <= priority(71) and not req(71);
w857 <= not priority(72) and not w856;
w858 <= not priority(73) and w857;
w859 <= not w855 and w858;
w860 <= not priority(73) and req(72);
w861 <= not req(73) and not req(74);
w862 <= not w860 and w861;
w863 <= not w859 and w862;
w864 <= priority(74) and not req(74);
w865 <= not priority(75) and not w864;
w866 <= not priority(76) and w865;
w867 <= not w863 and w866;
w868 <= not priority(76) and req(75);
w869 <= not req(76) and not req(77);
w870 <= not w868 and w869;
w871 <= not w867 and w870;
w872 <= priority(77) and not req(77);
w873 <= not priority(78) and not w872;
w874 <= not priority(79) and w873;
w875 <= not w871 and w874;
w876 <= not priority(79) and req(78);
w877 <= not req(79) and not req(80);
w878 <= not w876 and w877;
w879 <= not w875 and w878;
w880 <= priority(80) and not req(80);
w881 <= not priority(81) and not w880;
w882 <= not priority(82) and w881;
w883 <= not w879 and w882;
w884 <= not priority(82) and req(81);
w885 <= not req(82) and not req(83);
w886 <= not w884 and w885;
w887 <= not w883 and w886;
w888 <= priority(83) and not req(83);
w889 <= not priority(84) and not w888;
w890 <= not priority(85) and w889;
w891 <= not w887 and w890;
w892 <= not priority(85) and req(84);
w893 <= not req(85) and not req(86);
w894 <= not w892 and w893;
w895 <= not w891 and w894;
w896 <= priority(86) and not req(86);
w897 <= not priority(87) and not w896;
w898 <= not priority(88) and w897;
w899 <= not w895 and w898;
w900 <= not priority(88) and req(87);
w901 <= not req(88) and not req(89);
w902 <= not w900 and w901;
w903 <= not w899 and w902;
w904 <= priority(89) and not req(89);
w905 <= not priority(90) and not w904;
w906 <= not priority(91) and w905;
w907 <= not w903 and w906;
w908 <= not priority(91) and req(90);
w909 <= not req(91) and not req(92);
w910 <= not w908 and w909;
w911 <= not w907 and w910;
w912 <= priority(92) and not req(92);
w913 <= not priority(93) and not w912;
w914 <= not priority(94) and w913;
w915 <= not w911 and w914;
w916 <= not priority(94) and req(93);
w917 <= not req(94) and not req(95);
w918 <= not w916 and w917;
w919 <= not w915 and w918;
w920 <= priority(95) and not req(95);
w921 <= not priority(96) and not w920;
w922 <= not priority(97) and w921;
w923 <= not w919 and w922;
w924 <= not priority(97) and req(96);
w925 <= not req(97) and not req(98);
w926 <= not w924 and w925;
w927 <= not w923 and w926;
w928 <= priority(98) and not req(98);
w929 <= not priority(99) and not w928;
w930 <= not priority(100) and w929;
w931 <= not w927 and w930;
w932 <= not priority(100) and req(99);
w933 <= not req(100) and not req(101);
w934 <= not w932 and w933;
w935 <= not w931 and w934;
w936 <= priority(101) and not req(101);
w937 <= not priority(102) and not w936;
w938 <= not priority(103) and w937;
w939 <= not w935 and w938;
w940 <= not priority(103) and req(102);
w941 <= not req(103) and not req(104);
w942 <= not w940 and w941;
w943 <= not w939 and w942;
w944 <= priority(104) and not req(104);
w945 <= not priority(105) and not w944;
w946 <= not priority(106) and w945;
w947 <= not w943 and w946;
w948 <= not priority(106) and req(105);
w949 <= not req(106) and not req(107);
w950 <= not w948 and w949;
w951 <= not w947 and w950;
w952 <= priority(107) and not req(107);
w953 <= not priority(108) and not w952;
w954 <= not priority(109) and w953;
w955 <= not w951 and w954;
w956 <= not priority(109) and req(108);
w957 <= not req(109) and not req(110);
w958 <= not w956 and w957;
w959 <= not w955 and w958;
w960 <= priority(110) and not req(110);
w961 <= not priority(111) and not w960;
w962 <= not priority(112) and w961;
w963 <= not w959 and w962;
w964 <= not priority(112) and req(111);
w965 <= not req(112) and not req(113);
w966 <= not w964 and w965;
w967 <= not w963 and w966;
w968 <= priority(113) and not req(113);
w969 <= not priority(114) and not w968;
w970 <= not priority(115) and w969;
w971 <= not w967 and w970;
w972 <= not priority(115) and req(114);
w973 <= not req(115) and not req(116);
w974 <= not w972 and w973;
w975 <= not w971 and w974;
w976 <= priority(116) and not req(116);
w977 <= not priority(117) and not w976;
w978 <= not priority(118) and w977;
w979 <= not w975 and w978;
w980 <= not priority(118) and req(117);
w981 <= not req(118) and not req(119);
w982 <= not w980 and w981;
w983 <= not w979 and w982;
w984 <= priority(119) and not req(119);
w985 <= not priority(120) and not w984;
w986 <= not priority(121) and w985;
w987 <= not w983 and w986;
w988 <= not priority(121) and req(120);
w989 <= not req(121) and not req(122);
w990 <= not w988 and w989;
w991 <= not w987 and w990;
w992 <= priority(122) and not req(122);
w993 <= not priority(123) and not w992;
w994 <= not priority(124) and w993;
w995 <= not w991 and w994;
w996 <= not priority(124) and req(123);
w997 <= not req(124) and not req(125);
w998 <= not w996 and w997;
w999 <= not w995 and w998;
w1000 <= priority(125) and not req(125);
w1001 <= not priority(126) and not w1000;
w1002 <= not priority(127) and w1001;
w1003 <= not w999 and w1002;
w1004 <= not priority(127) and req(126);
w1005 <= not req(0) and not req(127);
w1006 <= not w1004 and w1005;
w1007 <= not w1003 and w1006;
w1008 <= priority(0) and not req(0);
w1009 <= not priority(1) and not w1008;
w1010 <= not priority(2) and w1009;
w1011 <= not w1007 and w1010;
w1012 <= not priority(2) and req(1);
w1013 <= req(2) and not w1012;
w1014 <= not w1011 and w1013;
w1015 <= w9 and not w344;
w1016 <= w14 and not w1015;
w1017 <= w18 and not w1016;
w1018 <= w22 and not w1017;
w1019 <= w26 and not w1018;
w1020 <= w30 and not w1019;
w1021 <= w34 and not w1020;
w1022 <= w38 and not w1021;
w1023 <= w42 and not w1022;
w1024 <= w46 and not w1023;
w1025 <= w50 and not w1024;
w1026 <= w54 and not w1025;
w1027 <= w58 and not w1026;
w1028 <= w62 and not w1027;
w1029 <= w66 and not w1028;
w1030 <= w70 and not w1029;
w1031 <= w74 and not w1030;
w1032 <= w78 and not w1031;
w1033 <= w82 and not w1032;
w1034 <= w86 and not w1033;
w1035 <= w90 and not w1034;
w1036 <= w94 and not w1035;
w1037 <= w98 and not w1036;
w1038 <= w102 and not w1037;
w1039 <= w106 and not w1038;
w1040 <= w110 and not w1039;
w1041 <= w114 and not w1040;
w1042 <= w118 and not w1041;
w1043 <= w122 and not w1042;
w1044 <= w126 and not w1043;
w1045 <= w130 and not w1044;
w1046 <= w134 and not w1045;
w1047 <= w138 and not w1046;
w1048 <= w142 and not w1047;
w1049 <= w146 and not w1048;
w1050 <= w150 and not w1049;
w1051 <= w154 and not w1050;
w1052 <= w158 and not w1051;
w1053 <= w162 and not w1052;
w1054 <= w166 and not w1053;
w1055 <= w170 and not w1054;
w1056 <= w174 and not w1055;
w1057 <= w178 and not w1056;
w1058 <= w182 and not w1057;
w1059 <= w186 and not w1058;
w1060 <= w190 and not w1059;
w1061 <= w194 and not w1060;
w1062 <= w198 and not w1061;
w1063 <= w202 and not w1062;
w1064 <= w206 and not w1063;
w1065 <= w210 and not w1064;
w1066 <= w214 and not w1065;
w1067 <= w218 and not w1066;
w1068 <= w222 and not w1067;
w1069 <= w226 and not w1068;
w1070 <= w230 and not w1069;
w1071 <= w234 and not w1070;
w1072 <= w238 and not w1071;
w1073 <= w242 and not w1072;
w1074 <= w246 and not w1073;
w1075 <= w250 and not w1074;
w1076 <= w254 and not w1075;
w1077 <= w258 and not w1076;
w1078 <= w262 and not w1077;
w1079 <= w266 and not w1078;
w1080 <= w270 and not w1079;
w1081 <= w274 and not w1080;
w1082 <= w278 and not w1081;
w1083 <= w282 and not w1082;
w1084 <= w286 and not w1083;
w1085 <= w290 and not w1084;
w1086 <= w294 and not w1085;
w1087 <= w298 and not w1086;
w1088 <= w302 and not w1087;
w1089 <= w306 and not w1088;
w1090 <= w310 and not w1089;
w1091 <= w314 and not w1090;
w1092 <= w318 and not w1091;
w1093 <= w322 and not w1092;
w1094 <= w326 and not w1093;
w1095 <= w330 and not w1094;
w1096 <= w334 and not w1095;
w1097 <= not req(0) and not req(1);
w1098 <= not w336 and w1097;
w1099 <= not w1096 and w1098;
w1100 <= not priority(3) and w1;
w1101 <= not w1099 and w1100;
w1102 <= not priority(3) and req(2);
w1103 <= req(3) and not w1102;
w1104 <= not w1101 and w1103;
w1105 <= w348 and not w681;
w1106 <= w353 and not w1105;
w1107 <= w357 and not w1106;
w1108 <= w361 and not w1107;
w1109 <= w365 and not w1108;
w1110 <= w369 and not w1109;
w1111 <= w373 and not w1110;
w1112 <= w377 and not w1111;
w1113 <= w381 and not w1112;
w1114 <= w385 and not w1113;
w1115 <= w389 and not w1114;
w1116 <= w393 and not w1115;
w1117 <= w397 and not w1116;
w1118 <= w401 and not w1117;
w1119 <= w405 and not w1118;
w1120 <= w409 and not w1119;
w1121 <= w413 and not w1120;
w1122 <= w417 and not w1121;
w1123 <= w421 and not w1122;
w1124 <= w425 and not w1123;
w1125 <= w429 and not w1124;
w1126 <= w433 and not w1125;
w1127 <= w437 and not w1126;
w1128 <= w441 and not w1127;
w1129 <= w445 and not w1128;
w1130 <= w449 and not w1129;
w1131 <= w453 and not w1130;
w1132 <= w457 and not w1131;
w1133 <= w461 and not w1132;
w1134 <= w465 and not w1133;
w1135 <= w469 and not w1134;
w1136 <= w473 and not w1135;
w1137 <= w477 and not w1136;
w1138 <= w481 and not w1137;
w1139 <= w485 and not w1138;
w1140 <= w489 and not w1139;
w1141 <= w493 and not w1140;
w1142 <= w497 and not w1141;
w1143 <= w501 and not w1142;
w1144 <= w505 and not w1143;
w1145 <= w509 and not w1144;
w1146 <= w513 and not w1145;
w1147 <= w517 and not w1146;
w1148 <= w521 and not w1147;
w1149 <= w525 and not w1148;
w1150 <= w529 and not w1149;
w1151 <= w533 and not w1150;
w1152 <= w537 and not w1151;
w1153 <= w541 and not w1152;
w1154 <= w545 and not w1153;
w1155 <= w549 and not w1154;
w1156 <= w553 and not w1155;
w1157 <= w557 and not w1156;
w1158 <= w561 and not w1157;
w1159 <= w565 and not w1158;
w1160 <= w569 and not w1159;
w1161 <= w573 and not w1160;
w1162 <= w577 and not w1161;
w1163 <= w581 and not w1162;
w1164 <= w585 and not w1163;
w1165 <= w589 and not w1164;
w1166 <= w593 and not w1165;
w1167 <= w597 and not w1166;
w1168 <= w601 and not w1167;
w1169 <= w605 and not w1168;
w1170 <= w609 and not w1169;
w1171 <= w613 and not w1170;
w1172 <= w617 and not w1171;
w1173 <= w621 and not w1172;
w1174 <= w625 and not w1173;
w1175 <= w629 and not w1174;
w1176 <= w633 and not w1175;
w1177 <= w637 and not w1176;
w1178 <= w641 and not w1177;
w1179 <= w645 and not w1178;
w1180 <= w649 and not w1179;
w1181 <= w653 and not w1180;
w1182 <= w657 and not w1181;
w1183 <= w661 and not w1182;
w1184 <= w665 and not w1183;
w1185 <= w669 and not w1184;
w1186 <= w673 and not w1185;
w1187 <= not req(1) and not req(2);
w1188 <= not w675 and w1187;
w1189 <= not w1186 and w1188;
w1190 <= not priority(4) and w340;
w1191 <= not w1189 and w1190;
w1192 <= not priority(4) and req(3);
w1193 <= req(4) and not w1192;
w1194 <= not w1191 and w1193;
w1195 <= not w13 and w685;
w1196 <= w690 and not w1195;
w1197 <= w694 and not w1196;
w1198 <= w698 and not w1197;
w1199 <= w702 and not w1198;
w1200 <= w706 and not w1199;
w1201 <= w710 and not w1200;
w1202 <= w714 and not w1201;
w1203 <= w718 and not w1202;
w1204 <= w722 and not w1203;
w1205 <= w726 and not w1204;
w1206 <= w730 and not w1205;
w1207 <= w734 and not w1206;
w1208 <= w738 and not w1207;
w1209 <= w742 and not w1208;
w1210 <= w746 and not w1209;
w1211 <= w750 and not w1210;
w1212 <= w754 and not w1211;
w1213 <= w758 and not w1212;
w1214 <= w762 and not w1213;
w1215 <= w766 and not w1214;
w1216 <= w770 and not w1215;
w1217 <= w774 and not w1216;
w1218 <= w778 and not w1217;
w1219 <= w782 and not w1218;
w1220 <= w786 and not w1219;
w1221 <= w790 and not w1220;
w1222 <= w794 and not w1221;
w1223 <= w798 and not w1222;
w1224 <= w802 and not w1223;
w1225 <= w806 and not w1224;
w1226 <= w810 and not w1225;
w1227 <= w814 and not w1226;
w1228 <= w818 and not w1227;
w1229 <= w822 and not w1228;
w1230 <= w826 and not w1229;
w1231 <= w830 and not w1230;
w1232 <= w834 and not w1231;
w1233 <= w838 and not w1232;
w1234 <= w842 and not w1233;
w1235 <= w846 and not w1234;
w1236 <= w850 and not w1235;
w1237 <= w854 and not w1236;
w1238 <= w858 and not w1237;
w1239 <= w862 and not w1238;
w1240 <= w866 and not w1239;
w1241 <= w870 and not w1240;
w1242 <= w874 and not w1241;
w1243 <= w878 and not w1242;
w1244 <= w882 and not w1243;
w1245 <= w886 and not w1244;
w1246 <= w890 and not w1245;
w1247 <= w894 and not w1246;
w1248 <= w898 and not w1247;
w1249 <= w902 and not w1248;
w1250 <= w906 and not w1249;
w1251 <= w910 and not w1250;
w1252 <= w914 and not w1251;
w1253 <= w918 and not w1252;
w1254 <= w922 and not w1253;
w1255 <= w926 and not w1254;
w1256 <= w930 and not w1255;
w1257 <= w934 and not w1256;
w1258 <= w938 and not w1257;
w1259 <= w942 and not w1258;
w1260 <= w946 and not w1259;
w1261 <= w950 and not w1260;
w1262 <= w954 and not w1261;
w1263 <= w958 and not w1262;
w1264 <= w962 and not w1263;
w1265 <= w966 and not w1264;
w1266 <= w970 and not w1265;
w1267 <= w974 and not w1266;
w1268 <= w978 and not w1267;
w1269 <= w982 and not w1268;
w1270 <= w986 and not w1269;
w1271 <= w990 and not w1270;
w1272 <= w994 and not w1271;
w1273 <= w998 and not w1272;
w1274 <= w1002 and not w1273;
w1275 <= w1006 and not w1274;
w1276 <= w1010 and not w1275;
w1277 <= w2 and not w1012;
w1278 <= not w1276 and w1277;
w1279 <= w6 and not w1278;
w1280 <= req(5) and not w8;
w1281 <= not w1279 and w1280;
w1282 <= w17 and not w352;
w1283 <= w22 and not w1282;
w1284 <= w26 and not w1283;
w1285 <= w30 and not w1284;
w1286 <= w34 and not w1285;
w1287 <= w38 and not w1286;
w1288 <= w42 and not w1287;
w1289 <= w46 and not w1288;
w1290 <= w50 and not w1289;
w1291 <= w54 and not w1290;
w1292 <= w58 and not w1291;
w1293 <= w62 and not w1292;
w1294 <= w66 and not w1293;
w1295 <= w70 and not w1294;
w1296 <= w74 and not w1295;
w1297 <= w78 and not w1296;
w1298 <= w82 and not w1297;
w1299 <= w86 and not w1298;
w1300 <= w90 and not w1299;
w1301 <= w94 and not w1300;
w1302 <= w98 and not w1301;
w1303 <= w102 and not w1302;
w1304 <= w106 and not w1303;
w1305 <= w110 and not w1304;
w1306 <= w114 and not w1305;
w1307 <= w118 and not w1306;
w1308 <= w122 and not w1307;
w1309 <= w126 and not w1308;
w1310 <= w130 and not w1309;
w1311 <= w134 and not w1310;
w1312 <= w138 and not w1311;
w1313 <= w142 and not w1312;
w1314 <= w146 and not w1313;
w1315 <= w150 and not w1314;
w1316 <= w154 and not w1315;
w1317 <= w158 and not w1316;
w1318 <= w162 and not w1317;
w1319 <= w166 and not w1318;
w1320 <= w170 and not w1319;
w1321 <= w174 and not w1320;
w1322 <= w178 and not w1321;
w1323 <= w182 and not w1322;
w1324 <= w186 and not w1323;
w1325 <= w190 and not w1324;
w1326 <= w194 and not w1325;
w1327 <= w198 and not w1326;
w1328 <= w202 and not w1327;
w1329 <= w206 and not w1328;
w1330 <= w210 and not w1329;
w1331 <= w214 and not w1330;
w1332 <= w218 and not w1331;
w1333 <= w222 and not w1332;
w1334 <= w226 and not w1333;
w1335 <= w230 and not w1334;
w1336 <= w234 and not w1335;
w1337 <= w238 and not w1336;
w1338 <= w242 and not w1337;
w1339 <= w246 and not w1338;
w1340 <= w250 and not w1339;
w1341 <= w254 and not w1340;
w1342 <= w258 and not w1341;
w1343 <= w262 and not w1342;
w1344 <= w266 and not w1343;
w1345 <= w270 and not w1344;
w1346 <= w274 and not w1345;
w1347 <= w278 and not w1346;
w1348 <= w282 and not w1347;
w1349 <= w286 and not w1348;
w1350 <= w290 and not w1349;
w1351 <= w294 and not w1350;
w1352 <= w298 and not w1351;
w1353 <= w302 and not w1352;
w1354 <= w306 and not w1353;
w1355 <= w310 and not w1354;
w1356 <= w314 and not w1355;
w1357 <= w318 and not w1356;
w1358 <= w322 and not w1357;
w1359 <= w326 and not w1358;
w1360 <= w330 and not w1359;
w1361 <= w334 and not w1360;
w1362 <= w1098 and not w1361;
w1363 <= w1100 and not w1362;
w1364 <= w341 and not w1102;
w1365 <= not w1363 and w1364;
w1366 <= w345 and not w1365;
w1367 <= req(6) and not w347;
w1368 <= not w1366 and w1367;
w1369 <= w356 and not w689;
w1370 <= w361 and not w1369;
w1371 <= w365 and not w1370;
w1372 <= w369 and not w1371;
w1373 <= w373 and not w1372;
w1374 <= w377 and not w1373;
w1375 <= w381 and not w1374;
w1376 <= w385 and not w1375;
w1377 <= w389 and not w1376;
w1378 <= w393 and not w1377;
w1379 <= w397 and not w1378;
w1380 <= w401 and not w1379;
w1381 <= w405 and not w1380;
w1382 <= w409 and not w1381;
w1383 <= w413 and not w1382;
w1384 <= w417 and not w1383;
w1385 <= w421 and not w1384;
w1386 <= w425 and not w1385;
w1387 <= w429 and not w1386;
w1388 <= w433 and not w1387;
w1389 <= w437 and not w1388;
w1390 <= w441 and not w1389;
w1391 <= w445 and not w1390;
w1392 <= w449 and not w1391;
w1393 <= w453 and not w1392;
w1394 <= w457 and not w1393;
w1395 <= w461 and not w1394;
w1396 <= w465 and not w1395;
w1397 <= w469 and not w1396;
w1398 <= w473 and not w1397;
w1399 <= w477 and not w1398;
w1400 <= w481 and not w1399;
w1401 <= w485 and not w1400;
w1402 <= w489 and not w1401;
w1403 <= w493 and not w1402;
w1404 <= w497 and not w1403;
w1405 <= w501 and not w1404;
w1406 <= w505 and not w1405;
w1407 <= w509 and not w1406;
w1408 <= w513 and not w1407;
w1409 <= w517 and not w1408;
w1410 <= w521 and not w1409;
w1411 <= w525 and not w1410;
w1412 <= w529 and not w1411;
w1413 <= w533 and not w1412;
w1414 <= w537 and not w1413;
w1415 <= w541 and not w1414;
w1416 <= w545 and not w1415;
w1417 <= w549 and not w1416;
w1418 <= w553 and not w1417;
w1419 <= w557 and not w1418;
w1420 <= w561 and not w1419;
w1421 <= w565 and not w1420;
w1422 <= w569 and not w1421;
w1423 <= w573 and not w1422;
w1424 <= w577 and not w1423;
w1425 <= w581 and not w1424;
w1426 <= w585 and not w1425;
w1427 <= w589 and not w1426;
w1428 <= w593 and not w1427;
w1429 <= w597 and not w1428;
w1430 <= w601 and not w1429;
w1431 <= w605 and not w1430;
w1432 <= w609 and not w1431;
w1433 <= w613 and not w1432;
w1434 <= w617 and not w1433;
w1435 <= w621 and not w1434;
w1436 <= w625 and not w1435;
w1437 <= w629 and not w1436;
w1438 <= w633 and not w1437;
w1439 <= w637 and not w1438;
w1440 <= w641 and not w1439;
w1441 <= w645 and not w1440;
w1442 <= w649 and not w1441;
w1443 <= w653 and not w1442;
w1444 <= w657 and not w1443;
w1445 <= w661 and not w1444;
w1446 <= w665 and not w1445;
w1447 <= w669 and not w1446;
w1448 <= w673 and not w1447;
w1449 <= w1188 and not w1448;
w1450 <= w1190 and not w1449;
w1451 <= w678 and not w1192;
w1452 <= not w1450 and w1451;
w1453 <= w682 and not w1452;
w1454 <= req(7) and not w684;
w1455 <= not w1453 and w1454;
w1456 <= not w21 and w693;
w1457 <= w698 and not w1456;
w1458 <= w702 and not w1457;
w1459 <= w706 and not w1458;
w1460 <= w710 and not w1459;
w1461 <= w714 and not w1460;
w1462 <= w718 and not w1461;
w1463 <= w722 and not w1462;
w1464 <= w726 and not w1463;
w1465 <= w730 and not w1464;
w1466 <= w734 and not w1465;
w1467 <= w738 and not w1466;
w1468 <= w742 and not w1467;
w1469 <= w746 and not w1468;
w1470 <= w750 and not w1469;
w1471 <= w754 and not w1470;
w1472 <= w758 and not w1471;
w1473 <= w762 and not w1472;
w1474 <= w766 and not w1473;
w1475 <= w770 and not w1474;
w1476 <= w774 and not w1475;
w1477 <= w778 and not w1476;
w1478 <= w782 and not w1477;
w1479 <= w786 and not w1478;
w1480 <= w790 and not w1479;
w1481 <= w794 and not w1480;
w1482 <= w798 and not w1481;
w1483 <= w802 and not w1482;
w1484 <= w806 and not w1483;
w1485 <= w810 and not w1484;
w1486 <= w814 and not w1485;
w1487 <= w818 and not w1486;
w1488 <= w822 and not w1487;
w1489 <= w826 and not w1488;
w1490 <= w830 and not w1489;
w1491 <= w834 and not w1490;
w1492 <= w838 and not w1491;
w1493 <= w842 and not w1492;
w1494 <= w846 and not w1493;
w1495 <= w850 and not w1494;
w1496 <= w854 and not w1495;
w1497 <= w858 and not w1496;
w1498 <= w862 and not w1497;
w1499 <= w866 and not w1498;
w1500 <= w870 and not w1499;
w1501 <= w874 and not w1500;
w1502 <= w878 and not w1501;
w1503 <= w882 and not w1502;
w1504 <= w886 and not w1503;
w1505 <= w890 and not w1504;
w1506 <= w894 and not w1505;
w1507 <= w898 and not w1506;
w1508 <= w902 and not w1507;
w1509 <= w906 and not w1508;
w1510 <= w910 and not w1509;
w1511 <= w914 and not w1510;
w1512 <= w918 and not w1511;
w1513 <= w922 and not w1512;
w1514 <= w926 and not w1513;
w1515 <= w930 and not w1514;
w1516 <= w934 and not w1515;
w1517 <= w938 and not w1516;
w1518 <= w942 and not w1517;
w1519 <= w946 and not w1518;
w1520 <= w950 and not w1519;
w1521 <= w954 and not w1520;
w1522 <= w958 and not w1521;
w1523 <= w962 and not w1522;
w1524 <= w966 and not w1523;
w1525 <= w970 and not w1524;
w1526 <= w974 and not w1525;
w1527 <= w978 and not w1526;
w1528 <= w982 and not w1527;
w1529 <= w986 and not w1528;
w1530 <= w990 and not w1529;
w1531 <= w994 and not w1530;
w1532 <= w998 and not w1531;
w1533 <= w1002 and not w1532;
w1534 <= w1006 and not w1533;
w1535 <= w1010 and not w1534;
w1536 <= w1277 and not w1535;
w1537 <= w6 and not w1536;
w1538 <= w10 and not w1537;
w1539 <= w14 and not w1538;
w1540 <= req(8) and not w16;
w1541 <= not w1539 and w1540;
w1542 <= w25 and not w360;
w1543 <= w30 and not w1542;
w1544 <= w34 and not w1543;
w1545 <= w38 and not w1544;
w1546 <= w42 and not w1545;
w1547 <= w46 and not w1546;
w1548 <= w50 and not w1547;
w1549 <= w54 and not w1548;
w1550 <= w58 and not w1549;
w1551 <= w62 and not w1550;
w1552 <= w66 and not w1551;
w1553 <= w70 and not w1552;
w1554 <= w74 and not w1553;
w1555 <= w78 and not w1554;
w1556 <= w82 and not w1555;
w1557 <= w86 and not w1556;
w1558 <= w90 and not w1557;
w1559 <= w94 and not w1558;
w1560 <= w98 and not w1559;
w1561 <= w102 and not w1560;
w1562 <= w106 and not w1561;
w1563 <= w110 and not w1562;
w1564 <= w114 and not w1563;
w1565 <= w118 and not w1564;
w1566 <= w122 and not w1565;
w1567 <= w126 and not w1566;
w1568 <= w130 and not w1567;
w1569 <= w134 and not w1568;
w1570 <= w138 and not w1569;
w1571 <= w142 and not w1570;
w1572 <= w146 and not w1571;
w1573 <= w150 and not w1572;
w1574 <= w154 and not w1573;
w1575 <= w158 and not w1574;
w1576 <= w162 and not w1575;
w1577 <= w166 and not w1576;
w1578 <= w170 and not w1577;
w1579 <= w174 and not w1578;
w1580 <= w178 and not w1579;
w1581 <= w182 and not w1580;
w1582 <= w186 and not w1581;
w1583 <= w190 and not w1582;
w1584 <= w194 and not w1583;
w1585 <= w198 and not w1584;
w1586 <= w202 and not w1585;
w1587 <= w206 and not w1586;
w1588 <= w210 and not w1587;
w1589 <= w214 and not w1588;
w1590 <= w218 and not w1589;
w1591 <= w222 and not w1590;
w1592 <= w226 and not w1591;
w1593 <= w230 and not w1592;
w1594 <= w234 and not w1593;
w1595 <= w238 and not w1594;
w1596 <= w242 and not w1595;
w1597 <= w246 and not w1596;
w1598 <= w250 and not w1597;
w1599 <= w254 and not w1598;
w1600 <= w258 and not w1599;
w1601 <= w262 and not w1600;
w1602 <= w266 and not w1601;
w1603 <= w270 and not w1602;
w1604 <= w274 and not w1603;
w1605 <= w278 and not w1604;
w1606 <= w282 and not w1605;
w1607 <= w286 and not w1606;
w1608 <= w290 and not w1607;
w1609 <= w294 and not w1608;
w1610 <= w298 and not w1609;
w1611 <= w302 and not w1610;
w1612 <= w306 and not w1611;
w1613 <= w310 and not w1612;
w1614 <= w314 and not w1613;
w1615 <= w318 and not w1614;
w1616 <= w322 and not w1615;
w1617 <= w326 and not w1616;
w1618 <= w330 and not w1617;
w1619 <= w334 and not w1618;
w1620 <= w1098 and not w1619;
w1621 <= w1100 and not w1620;
w1622 <= w1364 and not w1621;
w1623 <= w345 and not w1622;
w1624 <= w349 and not w1623;
w1625 <= w353 and not w1624;
w1626 <= req(9) and not w355;
w1627 <= not w1625 and w1626;
w1628 <= w364 and not w697;
w1629 <= w369 and not w1628;
w1630 <= w373 and not w1629;
w1631 <= w377 and not w1630;
w1632 <= w381 and not w1631;
w1633 <= w385 and not w1632;
w1634 <= w389 and not w1633;
w1635 <= w393 and not w1634;
w1636 <= w397 and not w1635;
w1637 <= w401 and not w1636;
w1638 <= w405 and not w1637;
w1639 <= w409 and not w1638;
w1640 <= w413 and not w1639;
w1641 <= w417 and not w1640;
w1642 <= w421 and not w1641;
w1643 <= w425 and not w1642;
w1644 <= w429 and not w1643;
w1645 <= w433 and not w1644;
w1646 <= w437 and not w1645;
w1647 <= w441 and not w1646;
w1648 <= w445 and not w1647;
w1649 <= w449 and not w1648;
w1650 <= w453 and not w1649;
w1651 <= w457 and not w1650;
w1652 <= w461 and not w1651;
w1653 <= w465 and not w1652;
w1654 <= w469 and not w1653;
w1655 <= w473 and not w1654;
w1656 <= w477 and not w1655;
w1657 <= w481 and not w1656;
w1658 <= w485 and not w1657;
w1659 <= w489 and not w1658;
w1660 <= w493 and not w1659;
w1661 <= w497 and not w1660;
w1662 <= w501 and not w1661;
w1663 <= w505 and not w1662;
w1664 <= w509 and not w1663;
w1665 <= w513 and not w1664;
w1666 <= w517 and not w1665;
w1667 <= w521 and not w1666;
w1668 <= w525 and not w1667;
w1669 <= w529 and not w1668;
w1670 <= w533 and not w1669;
w1671 <= w537 and not w1670;
w1672 <= w541 and not w1671;
w1673 <= w545 and not w1672;
w1674 <= w549 and not w1673;
w1675 <= w553 and not w1674;
w1676 <= w557 and not w1675;
w1677 <= w561 and not w1676;
w1678 <= w565 and not w1677;
w1679 <= w569 and not w1678;
w1680 <= w573 and not w1679;
w1681 <= w577 and not w1680;
w1682 <= w581 and not w1681;
w1683 <= w585 and not w1682;
w1684 <= w589 and not w1683;
w1685 <= w593 and not w1684;
w1686 <= w597 and not w1685;
w1687 <= w601 and not w1686;
w1688 <= w605 and not w1687;
w1689 <= w609 and not w1688;
w1690 <= w613 and not w1689;
w1691 <= w617 and not w1690;
w1692 <= w621 and not w1691;
w1693 <= w625 and not w1692;
w1694 <= w629 and not w1693;
w1695 <= w633 and not w1694;
w1696 <= w637 and not w1695;
w1697 <= w641 and not w1696;
w1698 <= w645 and not w1697;
w1699 <= w649 and not w1698;
w1700 <= w653 and not w1699;
w1701 <= w657 and not w1700;
w1702 <= w661 and not w1701;
w1703 <= w665 and not w1702;
w1704 <= w669 and not w1703;
w1705 <= w673 and not w1704;
w1706 <= w1188 and not w1705;
w1707 <= w1190 and not w1706;
w1708 <= w1451 and not w1707;
w1709 <= w682 and not w1708;
w1710 <= w686 and not w1709;
w1711 <= w690 and not w1710;
w1712 <= req(10) and not w692;
w1713 <= not w1711 and w1712;
w1714 <= not w29 and w701;
w1715 <= w706 and not w1714;
w1716 <= w710 and not w1715;
w1717 <= w714 and not w1716;
w1718 <= w718 and not w1717;
w1719 <= w722 and not w1718;
w1720 <= w726 and not w1719;
w1721 <= w730 and not w1720;
w1722 <= w734 and not w1721;
w1723 <= w738 and not w1722;
w1724 <= w742 and not w1723;
w1725 <= w746 and not w1724;
w1726 <= w750 and not w1725;
w1727 <= w754 and not w1726;
w1728 <= w758 and not w1727;
w1729 <= w762 and not w1728;
w1730 <= w766 and not w1729;
w1731 <= w770 and not w1730;
w1732 <= w774 and not w1731;
w1733 <= w778 and not w1732;
w1734 <= w782 and not w1733;
w1735 <= w786 and not w1734;
w1736 <= w790 and not w1735;
w1737 <= w794 and not w1736;
w1738 <= w798 and not w1737;
w1739 <= w802 and not w1738;
w1740 <= w806 and not w1739;
w1741 <= w810 and not w1740;
w1742 <= w814 and not w1741;
w1743 <= w818 and not w1742;
w1744 <= w822 and not w1743;
w1745 <= w826 and not w1744;
w1746 <= w830 and not w1745;
w1747 <= w834 and not w1746;
w1748 <= w838 and not w1747;
w1749 <= w842 and not w1748;
w1750 <= w846 and not w1749;
w1751 <= w850 and not w1750;
w1752 <= w854 and not w1751;
w1753 <= w858 and not w1752;
w1754 <= w862 and not w1753;
w1755 <= w866 and not w1754;
w1756 <= w870 and not w1755;
w1757 <= w874 and not w1756;
w1758 <= w878 and not w1757;
w1759 <= w882 and not w1758;
w1760 <= w886 and not w1759;
w1761 <= w890 and not w1760;
w1762 <= w894 and not w1761;
w1763 <= w898 and not w1762;
w1764 <= w902 and not w1763;
w1765 <= w906 and not w1764;
w1766 <= w910 and not w1765;
w1767 <= w914 and not w1766;
w1768 <= w918 and not w1767;
w1769 <= w922 and not w1768;
w1770 <= w926 and not w1769;
w1771 <= w930 and not w1770;
w1772 <= w934 and not w1771;
w1773 <= w938 and not w1772;
w1774 <= w942 and not w1773;
w1775 <= w946 and not w1774;
w1776 <= w950 and not w1775;
w1777 <= w954 and not w1776;
w1778 <= w958 and not w1777;
w1779 <= w962 and not w1778;
w1780 <= w966 and not w1779;
w1781 <= w970 and not w1780;
w1782 <= w974 and not w1781;
w1783 <= w978 and not w1782;
w1784 <= w982 and not w1783;
w1785 <= w986 and not w1784;
w1786 <= w990 and not w1785;
w1787 <= w994 and not w1786;
w1788 <= w998 and not w1787;
w1789 <= w1002 and not w1788;
w1790 <= w1006 and not w1789;
w1791 <= w1010 and not w1790;
w1792 <= w1277 and not w1791;
w1793 <= w6 and not w1792;
w1794 <= w10 and not w1793;
w1795 <= w14 and not w1794;
w1796 <= w18 and not w1795;
w1797 <= w22 and not w1796;
w1798 <= req(11) and not w24;
w1799 <= not w1797 and w1798;
w1800 <= w33 and not w368;
w1801 <= w38 and not w1800;
w1802 <= w42 and not w1801;
w1803 <= w46 and not w1802;
w1804 <= w50 and not w1803;
w1805 <= w54 and not w1804;
w1806 <= w58 and not w1805;
w1807 <= w62 and not w1806;
w1808 <= w66 and not w1807;
w1809 <= w70 and not w1808;
w1810 <= w74 and not w1809;
w1811 <= w78 and not w1810;
w1812 <= w82 and not w1811;
w1813 <= w86 and not w1812;
w1814 <= w90 and not w1813;
w1815 <= w94 and not w1814;
w1816 <= w98 and not w1815;
w1817 <= w102 and not w1816;
w1818 <= w106 and not w1817;
w1819 <= w110 and not w1818;
w1820 <= w114 and not w1819;
w1821 <= w118 and not w1820;
w1822 <= w122 and not w1821;
w1823 <= w126 and not w1822;
w1824 <= w130 and not w1823;
w1825 <= w134 and not w1824;
w1826 <= w138 and not w1825;
w1827 <= w142 and not w1826;
w1828 <= w146 and not w1827;
w1829 <= w150 and not w1828;
w1830 <= w154 and not w1829;
w1831 <= w158 and not w1830;
w1832 <= w162 and not w1831;
w1833 <= w166 and not w1832;
w1834 <= w170 and not w1833;
w1835 <= w174 and not w1834;
w1836 <= w178 and not w1835;
w1837 <= w182 and not w1836;
w1838 <= w186 and not w1837;
w1839 <= w190 and not w1838;
w1840 <= w194 and not w1839;
w1841 <= w198 and not w1840;
w1842 <= w202 and not w1841;
w1843 <= w206 and not w1842;
w1844 <= w210 and not w1843;
w1845 <= w214 and not w1844;
w1846 <= w218 and not w1845;
w1847 <= w222 and not w1846;
w1848 <= w226 and not w1847;
w1849 <= w230 and not w1848;
w1850 <= w234 and not w1849;
w1851 <= w238 and not w1850;
w1852 <= w242 and not w1851;
w1853 <= w246 and not w1852;
w1854 <= w250 and not w1853;
w1855 <= w254 and not w1854;
w1856 <= w258 and not w1855;
w1857 <= w262 and not w1856;
w1858 <= w266 and not w1857;
w1859 <= w270 and not w1858;
w1860 <= w274 and not w1859;
w1861 <= w278 and not w1860;
w1862 <= w282 and not w1861;
w1863 <= w286 and not w1862;
w1864 <= w290 and not w1863;
w1865 <= w294 and not w1864;
w1866 <= w298 and not w1865;
w1867 <= w302 and not w1866;
w1868 <= w306 and not w1867;
w1869 <= w310 and not w1868;
w1870 <= w314 and not w1869;
w1871 <= w318 and not w1870;
w1872 <= w322 and not w1871;
w1873 <= w326 and not w1872;
w1874 <= w330 and not w1873;
w1875 <= w334 and not w1874;
w1876 <= w1098 and not w1875;
w1877 <= w1100 and not w1876;
w1878 <= w1364 and not w1877;
w1879 <= w345 and not w1878;
w1880 <= w349 and not w1879;
w1881 <= w353 and not w1880;
w1882 <= w357 and not w1881;
w1883 <= w361 and not w1882;
w1884 <= req(12) and not w363;
w1885 <= not w1883 and w1884;
w1886 <= w372 and not w705;
w1887 <= w377 and not w1886;
w1888 <= w381 and not w1887;
w1889 <= w385 and not w1888;
w1890 <= w389 and not w1889;
w1891 <= w393 and not w1890;
w1892 <= w397 and not w1891;
w1893 <= w401 and not w1892;
w1894 <= w405 and not w1893;
w1895 <= w409 and not w1894;
w1896 <= w413 and not w1895;
w1897 <= w417 and not w1896;
w1898 <= w421 and not w1897;
w1899 <= w425 and not w1898;
w1900 <= w429 and not w1899;
w1901 <= w433 and not w1900;
w1902 <= w437 and not w1901;
w1903 <= w441 and not w1902;
w1904 <= w445 and not w1903;
w1905 <= w449 and not w1904;
w1906 <= w453 and not w1905;
w1907 <= w457 and not w1906;
w1908 <= w461 and not w1907;
w1909 <= w465 and not w1908;
w1910 <= w469 and not w1909;
w1911 <= w473 and not w1910;
w1912 <= w477 and not w1911;
w1913 <= w481 and not w1912;
w1914 <= w485 and not w1913;
w1915 <= w489 and not w1914;
w1916 <= w493 and not w1915;
w1917 <= w497 and not w1916;
w1918 <= w501 and not w1917;
w1919 <= w505 and not w1918;
w1920 <= w509 and not w1919;
w1921 <= w513 and not w1920;
w1922 <= w517 and not w1921;
w1923 <= w521 and not w1922;
w1924 <= w525 and not w1923;
w1925 <= w529 and not w1924;
w1926 <= w533 and not w1925;
w1927 <= w537 and not w1926;
w1928 <= w541 and not w1927;
w1929 <= w545 and not w1928;
w1930 <= w549 and not w1929;
w1931 <= w553 and not w1930;
w1932 <= w557 and not w1931;
w1933 <= w561 and not w1932;
w1934 <= w565 and not w1933;
w1935 <= w569 and not w1934;
w1936 <= w573 and not w1935;
w1937 <= w577 and not w1936;
w1938 <= w581 and not w1937;
w1939 <= w585 and not w1938;
w1940 <= w589 and not w1939;
w1941 <= w593 and not w1940;
w1942 <= w597 and not w1941;
w1943 <= w601 and not w1942;
w1944 <= w605 and not w1943;
w1945 <= w609 and not w1944;
w1946 <= w613 and not w1945;
w1947 <= w617 and not w1946;
w1948 <= w621 and not w1947;
w1949 <= w625 and not w1948;
w1950 <= w629 and not w1949;
w1951 <= w633 and not w1950;
w1952 <= w637 and not w1951;
w1953 <= w641 and not w1952;
w1954 <= w645 and not w1953;
w1955 <= w649 and not w1954;
w1956 <= w653 and not w1955;
w1957 <= w657 and not w1956;
w1958 <= w661 and not w1957;
w1959 <= w665 and not w1958;
w1960 <= w669 and not w1959;
w1961 <= w673 and not w1960;
w1962 <= w1188 and not w1961;
w1963 <= w1190 and not w1962;
w1964 <= w1451 and not w1963;
w1965 <= w682 and not w1964;
w1966 <= w686 and not w1965;
w1967 <= w690 and not w1966;
w1968 <= w694 and not w1967;
w1969 <= w698 and not w1968;
w1970 <= req(13) and not w700;
w1971 <= not w1969 and w1970;
w1972 <= not w37 and w709;
w1973 <= w714 and not w1972;
w1974 <= w718 and not w1973;
w1975 <= w722 and not w1974;
w1976 <= w726 and not w1975;
w1977 <= w730 and not w1976;
w1978 <= w734 and not w1977;
w1979 <= w738 and not w1978;
w1980 <= w742 and not w1979;
w1981 <= w746 and not w1980;
w1982 <= w750 and not w1981;
w1983 <= w754 and not w1982;
w1984 <= w758 and not w1983;
w1985 <= w762 and not w1984;
w1986 <= w766 and not w1985;
w1987 <= w770 and not w1986;
w1988 <= w774 and not w1987;
w1989 <= w778 and not w1988;
w1990 <= w782 and not w1989;
w1991 <= w786 and not w1990;
w1992 <= w790 and not w1991;
w1993 <= w794 and not w1992;
w1994 <= w798 and not w1993;
w1995 <= w802 and not w1994;
w1996 <= w806 and not w1995;
w1997 <= w810 and not w1996;
w1998 <= w814 and not w1997;
w1999 <= w818 and not w1998;
w2000 <= w822 and not w1999;
w2001 <= w826 and not w2000;
w2002 <= w830 and not w2001;
w2003 <= w834 and not w2002;
w2004 <= w838 and not w2003;
w2005 <= w842 and not w2004;
w2006 <= w846 and not w2005;
w2007 <= w850 and not w2006;
w2008 <= w854 and not w2007;
w2009 <= w858 and not w2008;
w2010 <= w862 and not w2009;
w2011 <= w866 and not w2010;
w2012 <= w870 and not w2011;
w2013 <= w874 and not w2012;
w2014 <= w878 and not w2013;
w2015 <= w882 and not w2014;
w2016 <= w886 and not w2015;
w2017 <= w890 and not w2016;
w2018 <= w894 and not w2017;
w2019 <= w898 and not w2018;
w2020 <= w902 and not w2019;
w2021 <= w906 and not w2020;
w2022 <= w910 and not w2021;
w2023 <= w914 and not w2022;
w2024 <= w918 and not w2023;
w2025 <= w922 and not w2024;
w2026 <= w926 and not w2025;
w2027 <= w930 and not w2026;
w2028 <= w934 and not w2027;
w2029 <= w938 and not w2028;
w2030 <= w942 and not w2029;
w2031 <= w946 and not w2030;
w2032 <= w950 and not w2031;
w2033 <= w954 and not w2032;
w2034 <= w958 and not w2033;
w2035 <= w962 and not w2034;
w2036 <= w966 and not w2035;
w2037 <= w970 and not w2036;
w2038 <= w974 and not w2037;
w2039 <= w978 and not w2038;
w2040 <= w982 and not w2039;
w2041 <= w986 and not w2040;
w2042 <= w990 and not w2041;
w2043 <= w994 and not w2042;
w2044 <= w998 and not w2043;
w2045 <= w1002 and not w2044;
w2046 <= w1006 and not w2045;
w2047 <= w1010 and not w2046;
w2048 <= w1277 and not w2047;
w2049 <= w6 and not w2048;
w2050 <= w10 and not w2049;
w2051 <= w14 and not w2050;
w2052 <= w18 and not w2051;
w2053 <= w22 and not w2052;
w2054 <= w26 and not w2053;
w2055 <= w30 and not w2054;
w2056 <= req(14) and not w32;
w2057 <= not w2055 and w2056;
w2058 <= w41 and not w376;
w2059 <= w46 and not w2058;
w2060 <= w50 and not w2059;
w2061 <= w54 and not w2060;
w2062 <= w58 and not w2061;
w2063 <= w62 and not w2062;
w2064 <= w66 and not w2063;
w2065 <= w70 and not w2064;
w2066 <= w74 and not w2065;
w2067 <= w78 and not w2066;
w2068 <= w82 and not w2067;
w2069 <= w86 and not w2068;
w2070 <= w90 and not w2069;
w2071 <= w94 and not w2070;
w2072 <= w98 and not w2071;
w2073 <= w102 and not w2072;
w2074 <= w106 and not w2073;
w2075 <= w110 and not w2074;
w2076 <= w114 and not w2075;
w2077 <= w118 and not w2076;
w2078 <= w122 and not w2077;
w2079 <= w126 and not w2078;
w2080 <= w130 and not w2079;
w2081 <= w134 and not w2080;
w2082 <= w138 and not w2081;
w2083 <= w142 and not w2082;
w2084 <= w146 and not w2083;
w2085 <= w150 and not w2084;
w2086 <= w154 and not w2085;
w2087 <= w158 and not w2086;
w2088 <= w162 and not w2087;
w2089 <= w166 and not w2088;
w2090 <= w170 and not w2089;
w2091 <= w174 and not w2090;
w2092 <= w178 and not w2091;
w2093 <= w182 and not w2092;
w2094 <= w186 and not w2093;
w2095 <= w190 and not w2094;
w2096 <= w194 and not w2095;
w2097 <= w198 and not w2096;
w2098 <= w202 and not w2097;
w2099 <= w206 and not w2098;
w2100 <= w210 and not w2099;
w2101 <= w214 and not w2100;
w2102 <= w218 and not w2101;
w2103 <= w222 and not w2102;
w2104 <= w226 and not w2103;
w2105 <= w230 and not w2104;
w2106 <= w234 and not w2105;
w2107 <= w238 and not w2106;
w2108 <= w242 and not w2107;
w2109 <= w246 and not w2108;
w2110 <= w250 and not w2109;
w2111 <= w254 and not w2110;
w2112 <= w258 and not w2111;
w2113 <= w262 and not w2112;
w2114 <= w266 and not w2113;
w2115 <= w270 and not w2114;
w2116 <= w274 and not w2115;
w2117 <= w278 and not w2116;
w2118 <= w282 and not w2117;
w2119 <= w286 and not w2118;
w2120 <= w290 and not w2119;
w2121 <= w294 and not w2120;
w2122 <= w298 and not w2121;
w2123 <= w302 and not w2122;
w2124 <= w306 and not w2123;
w2125 <= w310 and not w2124;
w2126 <= w314 and not w2125;
w2127 <= w318 and not w2126;
w2128 <= w322 and not w2127;
w2129 <= w326 and not w2128;
w2130 <= w330 and not w2129;
w2131 <= w334 and not w2130;
w2132 <= w1098 and not w2131;
w2133 <= w1100 and not w2132;
w2134 <= w1364 and not w2133;
w2135 <= w345 and not w2134;
w2136 <= w349 and not w2135;
w2137 <= w353 and not w2136;
w2138 <= w357 and not w2137;
w2139 <= w361 and not w2138;
w2140 <= w365 and not w2139;
w2141 <= w369 and not w2140;
w2142 <= req(15) and not w371;
w2143 <= not w2141 and w2142;
w2144 <= w380 and not w713;
w2145 <= w385 and not w2144;
w2146 <= w389 and not w2145;
w2147 <= w393 and not w2146;
w2148 <= w397 and not w2147;
w2149 <= w401 and not w2148;
w2150 <= w405 and not w2149;
w2151 <= w409 and not w2150;
w2152 <= w413 and not w2151;
w2153 <= w417 and not w2152;
w2154 <= w421 and not w2153;
w2155 <= w425 and not w2154;
w2156 <= w429 and not w2155;
w2157 <= w433 and not w2156;
w2158 <= w437 and not w2157;
w2159 <= w441 and not w2158;
w2160 <= w445 and not w2159;
w2161 <= w449 and not w2160;
w2162 <= w453 and not w2161;
w2163 <= w457 and not w2162;
w2164 <= w461 and not w2163;
w2165 <= w465 and not w2164;
w2166 <= w469 and not w2165;
w2167 <= w473 and not w2166;
w2168 <= w477 and not w2167;
w2169 <= w481 and not w2168;
w2170 <= w485 and not w2169;
w2171 <= w489 and not w2170;
w2172 <= w493 and not w2171;
w2173 <= w497 and not w2172;
w2174 <= w501 and not w2173;
w2175 <= w505 and not w2174;
w2176 <= w509 and not w2175;
w2177 <= w513 and not w2176;
w2178 <= w517 and not w2177;
w2179 <= w521 and not w2178;
w2180 <= w525 and not w2179;
w2181 <= w529 and not w2180;
w2182 <= w533 and not w2181;
w2183 <= w537 and not w2182;
w2184 <= w541 and not w2183;
w2185 <= w545 and not w2184;
w2186 <= w549 and not w2185;
w2187 <= w553 and not w2186;
w2188 <= w557 and not w2187;
w2189 <= w561 and not w2188;
w2190 <= w565 and not w2189;
w2191 <= w569 and not w2190;
w2192 <= w573 and not w2191;
w2193 <= w577 and not w2192;
w2194 <= w581 and not w2193;
w2195 <= w585 and not w2194;
w2196 <= w589 and not w2195;
w2197 <= w593 and not w2196;
w2198 <= w597 and not w2197;
w2199 <= w601 and not w2198;
w2200 <= w605 and not w2199;
w2201 <= w609 and not w2200;
w2202 <= w613 and not w2201;
w2203 <= w617 and not w2202;
w2204 <= w621 and not w2203;
w2205 <= w625 and not w2204;
w2206 <= w629 and not w2205;
w2207 <= w633 and not w2206;
w2208 <= w637 and not w2207;
w2209 <= w641 and not w2208;
w2210 <= w645 and not w2209;
w2211 <= w649 and not w2210;
w2212 <= w653 and not w2211;
w2213 <= w657 and not w2212;
w2214 <= w661 and not w2213;
w2215 <= w665 and not w2214;
w2216 <= w669 and not w2215;
w2217 <= w673 and not w2216;
w2218 <= w1188 and not w2217;
w2219 <= w1190 and not w2218;
w2220 <= w1451 and not w2219;
w2221 <= w682 and not w2220;
w2222 <= w686 and not w2221;
w2223 <= w690 and not w2222;
w2224 <= w694 and not w2223;
w2225 <= w698 and not w2224;
w2226 <= w702 and not w2225;
w2227 <= w706 and not w2226;
w2228 <= req(16) and not w708;
w2229 <= not w2227 and w2228;
w2230 <= not w45 and w717;
w2231 <= w722 and not w2230;
w2232 <= w726 and not w2231;
w2233 <= w730 and not w2232;
w2234 <= w734 and not w2233;
w2235 <= w738 and not w2234;
w2236 <= w742 and not w2235;
w2237 <= w746 and not w2236;
w2238 <= w750 and not w2237;
w2239 <= w754 and not w2238;
w2240 <= w758 and not w2239;
w2241 <= w762 and not w2240;
w2242 <= w766 and not w2241;
w2243 <= w770 and not w2242;
w2244 <= w774 and not w2243;
w2245 <= w778 and not w2244;
w2246 <= w782 and not w2245;
w2247 <= w786 and not w2246;
w2248 <= w790 and not w2247;
w2249 <= w794 and not w2248;
w2250 <= w798 and not w2249;
w2251 <= w802 and not w2250;
w2252 <= w806 and not w2251;
w2253 <= w810 and not w2252;
w2254 <= w814 and not w2253;
w2255 <= w818 and not w2254;
w2256 <= w822 and not w2255;
w2257 <= w826 and not w2256;
w2258 <= w830 and not w2257;
w2259 <= w834 and not w2258;
w2260 <= w838 and not w2259;
w2261 <= w842 and not w2260;
w2262 <= w846 and not w2261;
w2263 <= w850 and not w2262;
w2264 <= w854 and not w2263;
w2265 <= w858 and not w2264;
w2266 <= w862 and not w2265;
w2267 <= w866 and not w2266;
w2268 <= w870 and not w2267;
w2269 <= w874 and not w2268;
w2270 <= w878 and not w2269;
w2271 <= w882 and not w2270;
w2272 <= w886 and not w2271;
w2273 <= w890 and not w2272;
w2274 <= w894 and not w2273;
w2275 <= w898 and not w2274;
w2276 <= w902 and not w2275;
w2277 <= w906 and not w2276;
w2278 <= w910 and not w2277;
w2279 <= w914 and not w2278;
w2280 <= w918 and not w2279;
w2281 <= w922 and not w2280;
w2282 <= w926 and not w2281;
w2283 <= w930 and not w2282;
w2284 <= w934 and not w2283;
w2285 <= w938 and not w2284;
w2286 <= w942 and not w2285;
w2287 <= w946 and not w2286;
w2288 <= w950 and not w2287;
w2289 <= w954 and not w2288;
w2290 <= w958 and not w2289;
w2291 <= w962 and not w2290;
w2292 <= w966 and not w2291;
w2293 <= w970 and not w2292;
w2294 <= w974 and not w2293;
w2295 <= w978 and not w2294;
w2296 <= w982 and not w2295;
w2297 <= w986 and not w2296;
w2298 <= w990 and not w2297;
w2299 <= w994 and not w2298;
w2300 <= w998 and not w2299;
w2301 <= w1002 and not w2300;
w2302 <= w1006 and not w2301;
w2303 <= w1010 and not w2302;
w2304 <= w1277 and not w2303;
w2305 <= w6 and not w2304;
w2306 <= w10 and not w2305;
w2307 <= w14 and not w2306;
w2308 <= w18 and not w2307;
w2309 <= w22 and not w2308;
w2310 <= w26 and not w2309;
w2311 <= w30 and not w2310;
w2312 <= w34 and not w2311;
w2313 <= w38 and not w2312;
w2314 <= req(17) and not w40;
w2315 <= not w2313 and w2314;
w2316 <= w49 and not w384;
w2317 <= w54 and not w2316;
w2318 <= w58 and not w2317;
w2319 <= w62 and not w2318;
w2320 <= w66 and not w2319;
w2321 <= w70 and not w2320;
w2322 <= w74 and not w2321;
w2323 <= w78 and not w2322;
w2324 <= w82 and not w2323;
w2325 <= w86 and not w2324;
w2326 <= w90 and not w2325;
w2327 <= w94 and not w2326;
w2328 <= w98 and not w2327;
w2329 <= w102 and not w2328;
w2330 <= w106 and not w2329;
w2331 <= w110 and not w2330;
w2332 <= w114 and not w2331;
w2333 <= w118 and not w2332;
w2334 <= w122 and not w2333;
w2335 <= w126 and not w2334;
w2336 <= w130 and not w2335;
w2337 <= w134 and not w2336;
w2338 <= w138 and not w2337;
w2339 <= w142 and not w2338;
w2340 <= w146 and not w2339;
w2341 <= w150 and not w2340;
w2342 <= w154 and not w2341;
w2343 <= w158 and not w2342;
w2344 <= w162 and not w2343;
w2345 <= w166 and not w2344;
w2346 <= w170 and not w2345;
w2347 <= w174 and not w2346;
w2348 <= w178 and not w2347;
w2349 <= w182 and not w2348;
w2350 <= w186 and not w2349;
w2351 <= w190 and not w2350;
w2352 <= w194 and not w2351;
w2353 <= w198 and not w2352;
w2354 <= w202 and not w2353;
w2355 <= w206 and not w2354;
w2356 <= w210 and not w2355;
w2357 <= w214 and not w2356;
w2358 <= w218 and not w2357;
w2359 <= w222 and not w2358;
w2360 <= w226 and not w2359;
w2361 <= w230 and not w2360;
w2362 <= w234 and not w2361;
w2363 <= w238 and not w2362;
w2364 <= w242 and not w2363;
w2365 <= w246 and not w2364;
w2366 <= w250 and not w2365;
w2367 <= w254 and not w2366;
w2368 <= w258 and not w2367;
w2369 <= w262 and not w2368;
w2370 <= w266 and not w2369;
w2371 <= w270 and not w2370;
w2372 <= w274 and not w2371;
w2373 <= w278 and not w2372;
w2374 <= w282 and not w2373;
w2375 <= w286 and not w2374;
w2376 <= w290 and not w2375;
w2377 <= w294 and not w2376;
w2378 <= w298 and not w2377;
w2379 <= w302 and not w2378;
w2380 <= w306 and not w2379;
w2381 <= w310 and not w2380;
w2382 <= w314 and not w2381;
w2383 <= w318 and not w2382;
w2384 <= w322 and not w2383;
w2385 <= w326 and not w2384;
w2386 <= w330 and not w2385;
w2387 <= w334 and not w2386;
w2388 <= w1098 and not w2387;
w2389 <= w1100 and not w2388;
w2390 <= w1364 and not w2389;
w2391 <= w345 and not w2390;
w2392 <= w349 and not w2391;
w2393 <= w353 and not w2392;
w2394 <= w357 and not w2393;
w2395 <= w361 and not w2394;
w2396 <= w365 and not w2395;
w2397 <= w369 and not w2396;
w2398 <= w373 and not w2397;
w2399 <= w377 and not w2398;
w2400 <= req(18) and not w379;
w2401 <= not w2399 and w2400;
w2402 <= w388 and not w721;
w2403 <= w393 and not w2402;
w2404 <= w397 and not w2403;
w2405 <= w401 and not w2404;
w2406 <= w405 and not w2405;
w2407 <= w409 and not w2406;
w2408 <= w413 and not w2407;
w2409 <= w417 and not w2408;
w2410 <= w421 and not w2409;
w2411 <= w425 and not w2410;
w2412 <= w429 and not w2411;
w2413 <= w433 and not w2412;
w2414 <= w437 and not w2413;
w2415 <= w441 and not w2414;
w2416 <= w445 and not w2415;
w2417 <= w449 and not w2416;
w2418 <= w453 and not w2417;
w2419 <= w457 and not w2418;
w2420 <= w461 and not w2419;
w2421 <= w465 and not w2420;
w2422 <= w469 and not w2421;
w2423 <= w473 and not w2422;
w2424 <= w477 and not w2423;
w2425 <= w481 and not w2424;
w2426 <= w485 and not w2425;
w2427 <= w489 and not w2426;
w2428 <= w493 and not w2427;
w2429 <= w497 and not w2428;
w2430 <= w501 and not w2429;
w2431 <= w505 and not w2430;
w2432 <= w509 and not w2431;
w2433 <= w513 and not w2432;
w2434 <= w517 and not w2433;
w2435 <= w521 and not w2434;
w2436 <= w525 and not w2435;
w2437 <= w529 and not w2436;
w2438 <= w533 and not w2437;
w2439 <= w537 and not w2438;
w2440 <= w541 and not w2439;
w2441 <= w545 and not w2440;
w2442 <= w549 and not w2441;
w2443 <= w553 and not w2442;
w2444 <= w557 and not w2443;
w2445 <= w561 and not w2444;
w2446 <= w565 and not w2445;
w2447 <= w569 and not w2446;
w2448 <= w573 and not w2447;
w2449 <= w577 and not w2448;
w2450 <= w581 and not w2449;
w2451 <= w585 and not w2450;
w2452 <= w589 and not w2451;
w2453 <= w593 and not w2452;
w2454 <= w597 and not w2453;
w2455 <= w601 and not w2454;
w2456 <= w605 and not w2455;
w2457 <= w609 and not w2456;
w2458 <= w613 and not w2457;
w2459 <= w617 and not w2458;
w2460 <= w621 and not w2459;
w2461 <= w625 and not w2460;
w2462 <= w629 and not w2461;
w2463 <= w633 and not w2462;
w2464 <= w637 and not w2463;
w2465 <= w641 and not w2464;
w2466 <= w645 and not w2465;
w2467 <= w649 and not w2466;
w2468 <= w653 and not w2467;
w2469 <= w657 and not w2468;
w2470 <= w661 and not w2469;
w2471 <= w665 and not w2470;
w2472 <= w669 and not w2471;
w2473 <= w673 and not w2472;
w2474 <= w1188 and not w2473;
w2475 <= w1190 and not w2474;
w2476 <= w1451 and not w2475;
w2477 <= w682 and not w2476;
w2478 <= w686 and not w2477;
w2479 <= w690 and not w2478;
w2480 <= w694 and not w2479;
w2481 <= w698 and not w2480;
w2482 <= w702 and not w2481;
w2483 <= w706 and not w2482;
w2484 <= w710 and not w2483;
w2485 <= w714 and not w2484;
w2486 <= req(19) and not w716;
w2487 <= not w2485 and w2486;
w2488 <= not w53 and w725;
w2489 <= w730 and not w2488;
w2490 <= w734 and not w2489;
w2491 <= w738 and not w2490;
w2492 <= w742 and not w2491;
w2493 <= w746 and not w2492;
w2494 <= w750 and not w2493;
w2495 <= w754 and not w2494;
w2496 <= w758 and not w2495;
w2497 <= w762 and not w2496;
w2498 <= w766 and not w2497;
w2499 <= w770 and not w2498;
w2500 <= w774 and not w2499;
w2501 <= w778 and not w2500;
w2502 <= w782 and not w2501;
w2503 <= w786 and not w2502;
w2504 <= w790 and not w2503;
w2505 <= w794 and not w2504;
w2506 <= w798 and not w2505;
w2507 <= w802 and not w2506;
w2508 <= w806 and not w2507;
w2509 <= w810 and not w2508;
w2510 <= w814 and not w2509;
w2511 <= w818 and not w2510;
w2512 <= w822 and not w2511;
w2513 <= w826 and not w2512;
w2514 <= w830 and not w2513;
w2515 <= w834 and not w2514;
w2516 <= w838 and not w2515;
w2517 <= w842 and not w2516;
w2518 <= w846 and not w2517;
w2519 <= w850 and not w2518;
w2520 <= w854 and not w2519;
w2521 <= w858 and not w2520;
w2522 <= w862 and not w2521;
w2523 <= w866 and not w2522;
w2524 <= w870 and not w2523;
w2525 <= w874 and not w2524;
w2526 <= w878 and not w2525;
w2527 <= w882 and not w2526;
w2528 <= w886 and not w2527;
w2529 <= w890 and not w2528;
w2530 <= w894 and not w2529;
w2531 <= w898 and not w2530;
w2532 <= w902 and not w2531;
w2533 <= w906 and not w2532;
w2534 <= w910 and not w2533;
w2535 <= w914 and not w2534;
w2536 <= w918 and not w2535;
w2537 <= w922 and not w2536;
w2538 <= w926 and not w2537;
w2539 <= w930 and not w2538;
w2540 <= w934 and not w2539;
w2541 <= w938 and not w2540;
w2542 <= w942 and not w2541;
w2543 <= w946 and not w2542;
w2544 <= w950 and not w2543;
w2545 <= w954 and not w2544;
w2546 <= w958 and not w2545;
w2547 <= w962 and not w2546;
w2548 <= w966 and not w2547;
w2549 <= w970 and not w2548;
w2550 <= w974 and not w2549;
w2551 <= w978 and not w2550;
w2552 <= w982 and not w2551;
w2553 <= w986 and not w2552;
w2554 <= w990 and not w2553;
w2555 <= w994 and not w2554;
w2556 <= w998 and not w2555;
w2557 <= w1002 and not w2556;
w2558 <= w1006 and not w2557;
w2559 <= w1010 and not w2558;
w2560 <= w1277 and not w2559;
w2561 <= w6 and not w2560;
w2562 <= w10 and not w2561;
w2563 <= w14 and not w2562;
w2564 <= w18 and not w2563;
w2565 <= w22 and not w2564;
w2566 <= w26 and not w2565;
w2567 <= w30 and not w2566;
w2568 <= w34 and not w2567;
w2569 <= w38 and not w2568;
w2570 <= w42 and not w2569;
w2571 <= w46 and not w2570;
w2572 <= req(20) and not w48;
w2573 <= not w2571 and w2572;
w2574 <= w57 and not w392;
w2575 <= w62 and not w2574;
w2576 <= w66 and not w2575;
w2577 <= w70 and not w2576;
w2578 <= w74 and not w2577;
w2579 <= w78 and not w2578;
w2580 <= w82 and not w2579;
w2581 <= w86 and not w2580;
w2582 <= w90 and not w2581;
w2583 <= w94 and not w2582;
w2584 <= w98 and not w2583;
w2585 <= w102 and not w2584;
w2586 <= w106 and not w2585;
w2587 <= w110 and not w2586;
w2588 <= w114 and not w2587;
w2589 <= w118 and not w2588;
w2590 <= w122 and not w2589;
w2591 <= w126 and not w2590;
w2592 <= w130 and not w2591;
w2593 <= w134 and not w2592;
w2594 <= w138 and not w2593;
w2595 <= w142 and not w2594;
w2596 <= w146 and not w2595;
w2597 <= w150 and not w2596;
w2598 <= w154 and not w2597;
w2599 <= w158 and not w2598;
w2600 <= w162 and not w2599;
w2601 <= w166 and not w2600;
w2602 <= w170 and not w2601;
w2603 <= w174 and not w2602;
w2604 <= w178 and not w2603;
w2605 <= w182 and not w2604;
w2606 <= w186 and not w2605;
w2607 <= w190 and not w2606;
w2608 <= w194 and not w2607;
w2609 <= w198 and not w2608;
w2610 <= w202 and not w2609;
w2611 <= w206 and not w2610;
w2612 <= w210 and not w2611;
w2613 <= w214 and not w2612;
w2614 <= w218 and not w2613;
w2615 <= w222 and not w2614;
w2616 <= w226 and not w2615;
w2617 <= w230 and not w2616;
w2618 <= w234 and not w2617;
w2619 <= w238 and not w2618;
w2620 <= w242 and not w2619;
w2621 <= w246 and not w2620;
w2622 <= w250 and not w2621;
w2623 <= w254 and not w2622;
w2624 <= w258 and not w2623;
w2625 <= w262 and not w2624;
w2626 <= w266 and not w2625;
w2627 <= w270 and not w2626;
w2628 <= w274 and not w2627;
w2629 <= w278 and not w2628;
w2630 <= w282 and not w2629;
w2631 <= w286 and not w2630;
w2632 <= w290 and not w2631;
w2633 <= w294 and not w2632;
w2634 <= w298 and not w2633;
w2635 <= w302 and not w2634;
w2636 <= w306 and not w2635;
w2637 <= w310 and not w2636;
w2638 <= w314 and not w2637;
w2639 <= w318 and not w2638;
w2640 <= w322 and not w2639;
w2641 <= w326 and not w2640;
w2642 <= w330 and not w2641;
w2643 <= w334 and not w2642;
w2644 <= w1098 and not w2643;
w2645 <= w1100 and not w2644;
w2646 <= w1364 and not w2645;
w2647 <= w345 and not w2646;
w2648 <= w349 and not w2647;
w2649 <= w353 and not w2648;
w2650 <= w357 and not w2649;
w2651 <= w361 and not w2650;
w2652 <= w365 and not w2651;
w2653 <= w369 and not w2652;
w2654 <= w373 and not w2653;
w2655 <= w377 and not w2654;
w2656 <= w381 and not w2655;
w2657 <= w385 and not w2656;
w2658 <= req(21) and not w387;
w2659 <= not w2657 and w2658;
w2660 <= w396 and not w729;
w2661 <= w401 and not w2660;
w2662 <= w405 and not w2661;
w2663 <= w409 and not w2662;
w2664 <= w413 and not w2663;
w2665 <= w417 and not w2664;
w2666 <= w421 and not w2665;
w2667 <= w425 and not w2666;
w2668 <= w429 and not w2667;
w2669 <= w433 and not w2668;
w2670 <= w437 and not w2669;
w2671 <= w441 and not w2670;
w2672 <= w445 and not w2671;
w2673 <= w449 and not w2672;
w2674 <= w453 and not w2673;
w2675 <= w457 and not w2674;
w2676 <= w461 and not w2675;
w2677 <= w465 and not w2676;
w2678 <= w469 and not w2677;
w2679 <= w473 and not w2678;
w2680 <= w477 and not w2679;
w2681 <= w481 and not w2680;
w2682 <= w485 and not w2681;
w2683 <= w489 and not w2682;
w2684 <= w493 and not w2683;
w2685 <= w497 and not w2684;
w2686 <= w501 and not w2685;
w2687 <= w505 and not w2686;
w2688 <= w509 and not w2687;
w2689 <= w513 and not w2688;
w2690 <= w517 and not w2689;
w2691 <= w521 and not w2690;
w2692 <= w525 and not w2691;
w2693 <= w529 and not w2692;
w2694 <= w533 and not w2693;
w2695 <= w537 and not w2694;
w2696 <= w541 and not w2695;
w2697 <= w545 and not w2696;
w2698 <= w549 and not w2697;
w2699 <= w553 and not w2698;
w2700 <= w557 and not w2699;
w2701 <= w561 and not w2700;
w2702 <= w565 and not w2701;
w2703 <= w569 and not w2702;
w2704 <= w573 and not w2703;
w2705 <= w577 and not w2704;
w2706 <= w581 and not w2705;
w2707 <= w585 and not w2706;
w2708 <= w589 and not w2707;
w2709 <= w593 and not w2708;
w2710 <= w597 and not w2709;
w2711 <= w601 and not w2710;
w2712 <= w605 and not w2711;
w2713 <= w609 and not w2712;
w2714 <= w613 and not w2713;
w2715 <= w617 and not w2714;
w2716 <= w621 and not w2715;
w2717 <= w625 and not w2716;
w2718 <= w629 and not w2717;
w2719 <= w633 and not w2718;
w2720 <= w637 and not w2719;
w2721 <= w641 and not w2720;
w2722 <= w645 and not w2721;
w2723 <= w649 and not w2722;
w2724 <= w653 and not w2723;
w2725 <= w657 and not w2724;
w2726 <= w661 and not w2725;
w2727 <= w665 and not w2726;
w2728 <= w669 and not w2727;
w2729 <= w673 and not w2728;
w2730 <= w1188 and not w2729;
w2731 <= w1190 and not w2730;
w2732 <= w1451 and not w2731;
w2733 <= w682 and not w2732;
w2734 <= w686 and not w2733;
w2735 <= w690 and not w2734;
w2736 <= w694 and not w2735;
w2737 <= w698 and not w2736;
w2738 <= w702 and not w2737;
w2739 <= w706 and not w2738;
w2740 <= w710 and not w2739;
w2741 <= w714 and not w2740;
w2742 <= w718 and not w2741;
w2743 <= w722 and not w2742;
w2744 <= req(22) and not w724;
w2745 <= not w2743 and w2744;
w2746 <= not w61 and w733;
w2747 <= w738 and not w2746;
w2748 <= w742 and not w2747;
w2749 <= w746 and not w2748;
w2750 <= w750 and not w2749;
w2751 <= w754 and not w2750;
w2752 <= w758 and not w2751;
w2753 <= w762 and not w2752;
w2754 <= w766 and not w2753;
w2755 <= w770 and not w2754;
w2756 <= w774 and not w2755;
w2757 <= w778 and not w2756;
w2758 <= w782 and not w2757;
w2759 <= w786 and not w2758;
w2760 <= w790 and not w2759;
w2761 <= w794 and not w2760;
w2762 <= w798 and not w2761;
w2763 <= w802 and not w2762;
w2764 <= w806 and not w2763;
w2765 <= w810 and not w2764;
w2766 <= w814 and not w2765;
w2767 <= w818 and not w2766;
w2768 <= w822 and not w2767;
w2769 <= w826 and not w2768;
w2770 <= w830 and not w2769;
w2771 <= w834 and not w2770;
w2772 <= w838 and not w2771;
w2773 <= w842 and not w2772;
w2774 <= w846 and not w2773;
w2775 <= w850 and not w2774;
w2776 <= w854 and not w2775;
w2777 <= w858 and not w2776;
w2778 <= w862 and not w2777;
w2779 <= w866 and not w2778;
w2780 <= w870 and not w2779;
w2781 <= w874 and not w2780;
w2782 <= w878 and not w2781;
w2783 <= w882 and not w2782;
w2784 <= w886 and not w2783;
w2785 <= w890 and not w2784;
w2786 <= w894 and not w2785;
w2787 <= w898 and not w2786;
w2788 <= w902 and not w2787;
w2789 <= w906 and not w2788;
w2790 <= w910 and not w2789;
w2791 <= w914 and not w2790;
w2792 <= w918 and not w2791;
w2793 <= w922 and not w2792;
w2794 <= w926 and not w2793;
w2795 <= w930 and not w2794;
w2796 <= w934 and not w2795;
w2797 <= w938 and not w2796;
w2798 <= w942 and not w2797;
w2799 <= w946 and not w2798;
w2800 <= w950 and not w2799;
w2801 <= w954 and not w2800;
w2802 <= w958 and not w2801;
w2803 <= w962 and not w2802;
w2804 <= w966 and not w2803;
w2805 <= w970 and not w2804;
w2806 <= w974 and not w2805;
w2807 <= w978 and not w2806;
w2808 <= w982 and not w2807;
w2809 <= w986 and not w2808;
w2810 <= w990 and not w2809;
w2811 <= w994 and not w2810;
w2812 <= w998 and not w2811;
w2813 <= w1002 and not w2812;
w2814 <= w1006 and not w2813;
w2815 <= w1010 and not w2814;
w2816 <= w1277 and not w2815;
w2817 <= w6 and not w2816;
w2818 <= w10 and not w2817;
w2819 <= w14 and not w2818;
w2820 <= w18 and not w2819;
w2821 <= w22 and not w2820;
w2822 <= w26 and not w2821;
w2823 <= w30 and not w2822;
w2824 <= w34 and not w2823;
w2825 <= w38 and not w2824;
w2826 <= w42 and not w2825;
w2827 <= w46 and not w2826;
w2828 <= w50 and not w2827;
w2829 <= w54 and not w2828;
w2830 <= req(23) and not w56;
w2831 <= not w2829 and w2830;
w2832 <= w65 and not w400;
w2833 <= w70 and not w2832;
w2834 <= w74 and not w2833;
w2835 <= w78 and not w2834;
w2836 <= w82 and not w2835;
w2837 <= w86 and not w2836;
w2838 <= w90 and not w2837;
w2839 <= w94 and not w2838;
w2840 <= w98 and not w2839;
w2841 <= w102 and not w2840;
w2842 <= w106 and not w2841;
w2843 <= w110 and not w2842;
w2844 <= w114 and not w2843;
w2845 <= w118 and not w2844;
w2846 <= w122 and not w2845;
w2847 <= w126 and not w2846;
w2848 <= w130 and not w2847;
w2849 <= w134 and not w2848;
w2850 <= w138 and not w2849;
w2851 <= w142 and not w2850;
w2852 <= w146 and not w2851;
w2853 <= w150 and not w2852;
w2854 <= w154 and not w2853;
w2855 <= w158 and not w2854;
w2856 <= w162 and not w2855;
w2857 <= w166 and not w2856;
w2858 <= w170 and not w2857;
w2859 <= w174 and not w2858;
w2860 <= w178 and not w2859;
w2861 <= w182 and not w2860;
w2862 <= w186 and not w2861;
w2863 <= w190 and not w2862;
w2864 <= w194 and not w2863;
w2865 <= w198 and not w2864;
w2866 <= w202 and not w2865;
w2867 <= w206 and not w2866;
w2868 <= w210 and not w2867;
w2869 <= w214 and not w2868;
w2870 <= w218 and not w2869;
w2871 <= w222 and not w2870;
w2872 <= w226 and not w2871;
w2873 <= w230 and not w2872;
w2874 <= w234 and not w2873;
w2875 <= w238 and not w2874;
w2876 <= w242 and not w2875;
w2877 <= w246 and not w2876;
w2878 <= w250 and not w2877;
w2879 <= w254 and not w2878;
w2880 <= w258 and not w2879;
w2881 <= w262 and not w2880;
w2882 <= w266 and not w2881;
w2883 <= w270 and not w2882;
w2884 <= w274 and not w2883;
w2885 <= w278 and not w2884;
w2886 <= w282 and not w2885;
w2887 <= w286 and not w2886;
w2888 <= w290 and not w2887;
w2889 <= w294 and not w2888;
w2890 <= w298 and not w2889;
w2891 <= w302 and not w2890;
w2892 <= w306 and not w2891;
w2893 <= w310 and not w2892;
w2894 <= w314 and not w2893;
w2895 <= w318 and not w2894;
w2896 <= w322 and not w2895;
w2897 <= w326 and not w2896;
w2898 <= w330 and not w2897;
w2899 <= w334 and not w2898;
w2900 <= w1098 and not w2899;
w2901 <= w1100 and not w2900;
w2902 <= w1364 and not w2901;
w2903 <= w345 and not w2902;
w2904 <= w349 and not w2903;
w2905 <= w353 and not w2904;
w2906 <= w357 and not w2905;
w2907 <= w361 and not w2906;
w2908 <= w365 and not w2907;
w2909 <= w369 and not w2908;
w2910 <= w373 and not w2909;
w2911 <= w377 and not w2910;
w2912 <= w381 and not w2911;
w2913 <= w385 and not w2912;
w2914 <= w389 and not w2913;
w2915 <= w393 and not w2914;
w2916 <= req(24) and not w395;
w2917 <= not w2915 and w2916;
w2918 <= w404 and not w737;
w2919 <= w409 and not w2918;
w2920 <= w413 and not w2919;
w2921 <= w417 and not w2920;
w2922 <= w421 and not w2921;
w2923 <= w425 and not w2922;
w2924 <= w429 and not w2923;
w2925 <= w433 and not w2924;
w2926 <= w437 and not w2925;
w2927 <= w441 and not w2926;
w2928 <= w445 and not w2927;
w2929 <= w449 and not w2928;
w2930 <= w453 and not w2929;
w2931 <= w457 and not w2930;
w2932 <= w461 and not w2931;
w2933 <= w465 and not w2932;
w2934 <= w469 and not w2933;
w2935 <= w473 and not w2934;
w2936 <= w477 and not w2935;
w2937 <= w481 and not w2936;
w2938 <= w485 and not w2937;
w2939 <= w489 and not w2938;
w2940 <= w493 and not w2939;
w2941 <= w497 and not w2940;
w2942 <= w501 and not w2941;
w2943 <= w505 and not w2942;
w2944 <= w509 and not w2943;
w2945 <= w513 and not w2944;
w2946 <= w517 and not w2945;
w2947 <= w521 and not w2946;
w2948 <= w525 and not w2947;
w2949 <= w529 and not w2948;
w2950 <= w533 and not w2949;
w2951 <= w537 and not w2950;
w2952 <= w541 and not w2951;
w2953 <= w545 and not w2952;
w2954 <= w549 and not w2953;
w2955 <= w553 and not w2954;
w2956 <= w557 and not w2955;
w2957 <= w561 and not w2956;
w2958 <= w565 and not w2957;
w2959 <= w569 and not w2958;
w2960 <= w573 and not w2959;
w2961 <= w577 and not w2960;
w2962 <= w581 and not w2961;
w2963 <= w585 and not w2962;
w2964 <= w589 and not w2963;
w2965 <= w593 and not w2964;
w2966 <= w597 and not w2965;
w2967 <= w601 and not w2966;
w2968 <= w605 and not w2967;
w2969 <= w609 and not w2968;
w2970 <= w613 and not w2969;
w2971 <= w617 and not w2970;
w2972 <= w621 and not w2971;
w2973 <= w625 and not w2972;
w2974 <= w629 and not w2973;
w2975 <= w633 and not w2974;
w2976 <= w637 and not w2975;
w2977 <= w641 and not w2976;
w2978 <= w645 and not w2977;
w2979 <= w649 and not w2978;
w2980 <= w653 and not w2979;
w2981 <= w657 and not w2980;
w2982 <= w661 and not w2981;
w2983 <= w665 and not w2982;
w2984 <= w669 and not w2983;
w2985 <= w673 and not w2984;
w2986 <= w1188 and not w2985;
w2987 <= w1190 and not w2986;
w2988 <= w1451 and not w2987;
w2989 <= w682 and not w2988;
w2990 <= w686 and not w2989;
w2991 <= w690 and not w2990;
w2992 <= w694 and not w2991;
w2993 <= w698 and not w2992;
w2994 <= w702 and not w2993;
w2995 <= w706 and not w2994;
w2996 <= w710 and not w2995;
w2997 <= w714 and not w2996;
w2998 <= w718 and not w2997;
w2999 <= w722 and not w2998;
w3000 <= w726 and not w2999;
w3001 <= w730 and not w3000;
w3002 <= req(25) and not w732;
w3003 <= not w3001 and w3002;
w3004 <= not w69 and w741;
w3005 <= w746 and not w3004;
w3006 <= w750 and not w3005;
w3007 <= w754 and not w3006;
w3008 <= w758 and not w3007;
w3009 <= w762 and not w3008;
w3010 <= w766 and not w3009;
w3011 <= w770 and not w3010;
w3012 <= w774 and not w3011;
w3013 <= w778 and not w3012;
w3014 <= w782 and not w3013;
w3015 <= w786 and not w3014;
w3016 <= w790 and not w3015;
w3017 <= w794 and not w3016;
w3018 <= w798 and not w3017;
w3019 <= w802 and not w3018;
w3020 <= w806 and not w3019;
w3021 <= w810 and not w3020;
w3022 <= w814 and not w3021;
w3023 <= w818 and not w3022;
w3024 <= w822 and not w3023;
w3025 <= w826 and not w3024;
w3026 <= w830 and not w3025;
w3027 <= w834 and not w3026;
w3028 <= w838 and not w3027;
w3029 <= w842 and not w3028;
w3030 <= w846 and not w3029;
w3031 <= w850 and not w3030;
w3032 <= w854 and not w3031;
w3033 <= w858 and not w3032;
w3034 <= w862 and not w3033;
w3035 <= w866 and not w3034;
w3036 <= w870 and not w3035;
w3037 <= w874 and not w3036;
w3038 <= w878 and not w3037;
w3039 <= w882 and not w3038;
w3040 <= w886 and not w3039;
w3041 <= w890 and not w3040;
w3042 <= w894 and not w3041;
w3043 <= w898 and not w3042;
w3044 <= w902 and not w3043;
w3045 <= w906 and not w3044;
w3046 <= w910 and not w3045;
w3047 <= w914 and not w3046;
w3048 <= w918 and not w3047;
w3049 <= w922 and not w3048;
w3050 <= w926 and not w3049;
w3051 <= w930 and not w3050;
w3052 <= w934 and not w3051;
w3053 <= w938 and not w3052;
w3054 <= w942 and not w3053;
w3055 <= w946 and not w3054;
w3056 <= w950 and not w3055;
w3057 <= w954 and not w3056;
w3058 <= w958 and not w3057;
w3059 <= w962 and not w3058;
w3060 <= w966 and not w3059;
w3061 <= w970 and not w3060;
w3062 <= w974 and not w3061;
w3063 <= w978 and not w3062;
w3064 <= w982 and not w3063;
w3065 <= w986 and not w3064;
w3066 <= w990 and not w3065;
w3067 <= w994 and not w3066;
w3068 <= w998 and not w3067;
w3069 <= w1002 and not w3068;
w3070 <= w1006 and not w3069;
w3071 <= w1010 and not w3070;
w3072 <= w1277 and not w3071;
w3073 <= w6 and not w3072;
w3074 <= w10 and not w3073;
w3075 <= w14 and not w3074;
w3076 <= w18 and not w3075;
w3077 <= w22 and not w3076;
w3078 <= w26 and not w3077;
w3079 <= w30 and not w3078;
w3080 <= w34 and not w3079;
w3081 <= w38 and not w3080;
w3082 <= w42 and not w3081;
w3083 <= w46 and not w3082;
w3084 <= w50 and not w3083;
w3085 <= w54 and not w3084;
w3086 <= w58 and not w3085;
w3087 <= w62 and not w3086;
w3088 <= req(26) and not w64;
w3089 <= not w3087 and w3088;
w3090 <= w73 and not w408;
w3091 <= w78 and not w3090;
w3092 <= w82 and not w3091;
w3093 <= w86 and not w3092;
w3094 <= w90 and not w3093;
w3095 <= w94 and not w3094;
w3096 <= w98 and not w3095;
w3097 <= w102 and not w3096;
w3098 <= w106 and not w3097;
w3099 <= w110 and not w3098;
w3100 <= w114 and not w3099;
w3101 <= w118 and not w3100;
w3102 <= w122 and not w3101;
w3103 <= w126 and not w3102;
w3104 <= w130 and not w3103;
w3105 <= w134 and not w3104;
w3106 <= w138 and not w3105;
w3107 <= w142 and not w3106;
w3108 <= w146 and not w3107;
w3109 <= w150 and not w3108;
w3110 <= w154 and not w3109;
w3111 <= w158 and not w3110;
w3112 <= w162 and not w3111;
w3113 <= w166 and not w3112;
w3114 <= w170 and not w3113;
w3115 <= w174 and not w3114;
w3116 <= w178 and not w3115;
w3117 <= w182 and not w3116;
w3118 <= w186 and not w3117;
w3119 <= w190 and not w3118;
w3120 <= w194 and not w3119;
w3121 <= w198 and not w3120;
w3122 <= w202 and not w3121;
w3123 <= w206 and not w3122;
w3124 <= w210 and not w3123;
w3125 <= w214 and not w3124;
w3126 <= w218 and not w3125;
w3127 <= w222 and not w3126;
w3128 <= w226 and not w3127;
w3129 <= w230 and not w3128;
w3130 <= w234 and not w3129;
w3131 <= w238 and not w3130;
w3132 <= w242 and not w3131;
w3133 <= w246 and not w3132;
w3134 <= w250 and not w3133;
w3135 <= w254 and not w3134;
w3136 <= w258 and not w3135;
w3137 <= w262 and not w3136;
w3138 <= w266 and not w3137;
w3139 <= w270 and not w3138;
w3140 <= w274 and not w3139;
w3141 <= w278 and not w3140;
w3142 <= w282 and not w3141;
w3143 <= w286 and not w3142;
w3144 <= w290 and not w3143;
w3145 <= w294 and not w3144;
w3146 <= w298 and not w3145;
w3147 <= w302 and not w3146;
w3148 <= w306 and not w3147;
w3149 <= w310 and not w3148;
w3150 <= w314 and not w3149;
w3151 <= w318 and not w3150;
w3152 <= w322 and not w3151;
w3153 <= w326 and not w3152;
w3154 <= w330 and not w3153;
w3155 <= w334 and not w3154;
w3156 <= w1098 and not w3155;
w3157 <= w1100 and not w3156;
w3158 <= w1364 and not w3157;
w3159 <= w345 and not w3158;
w3160 <= w349 and not w3159;
w3161 <= w353 and not w3160;
w3162 <= w357 and not w3161;
w3163 <= w361 and not w3162;
w3164 <= w365 and not w3163;
w3165 <= w369 and not w3164;
w3166 <= w373 and not w3165;
w3167 <= w377 and not w3166;
w3168 <= w381 and not w3167;
w3169 <= w385 and not w3168;
w3170 <= w389 and not w3169;
w3171 <= w393 and not w3170;
w3172 <= w397 and not w3171;
w3173 <= w401 and not w3172;
w3174 <= req(27) and not w403;
w3175 <= not w3173 and w3174;
w3176 <= w412 and not w745;
w3177 <= w417 and not w3176;
w3178 <= w421 and not w3177;
w3179 <= w425 and not w3178;
w3180 <= w429 and not w3179;
w3181 <= w433 and not w3180;
w3182 <= w437 and not w3181;
w3183 <= w441 and not w3182;
w3184 <= w445 and not w3183;
w3185 <= w449 and not w3184;
w3186 <= w453 and not w3185;
w3187 <= w457 and not w3186;
w3188 <= w461 and not w3187;
w3189 <= w465 and not w3188;
w3190 <= w469 and not w3189;
w3191 <= w473 and not w3190;
w3192 <= w477 and not w3191;
w3193 <= w481 and not w3192;
w3194 <= w485 and not w3193;
w3195 <= w489 and not w3194;
w3196 <= w493 and not w3195;
w3197 <= w497 and not w3196;
w3198 <= w501 and not w3197;
w3199 <= w505 and not w3198;
w3200 <= w509 and not w3199;
w3201 <= w513 and not w3200;
w3202 <= w517 and not w3201;
w3203 <= w521 and not w3202;
w3204 <= w525 and not w3203;
w3205 <= w529 and not w3204;
w3206 <= w533 and not w3205;
w3207 <= w537 and not w3206;
w3208 <= w541 and not w3207;
w3209 <= w545 and not w3208;
w3210 <= w549 and not w3209;
w3211 <= w553 and not w3210;
w3212 <= w557 and not w3211;
w3213 <= w561 and not w3212;
w3214 <= w565 and not w3213;
w3215 <= w569 and not w3214;
w3216 <= w573 and not w3215;
w3217 <= w577 and not w3216;
w3218 <= w581 and not w3217;
w3219 <= w585 and not w3218;
w3220 <= w589 and not w3219;
w3221 <= w593 and not w3220;
w3222 <= w597 and not w3221;
w3223 <= w601 and not w3222;
w3224 <= w605 and not w3223;
w3225 <= w609 and not w3224;
w3226 <= w613 and not w3225;
w3227 <= w617 and not w3226;
w3228 <= w621 and not w3227;
w3229 <= w625 and not w3228;
w3230 <= w629 and not w3229;
w3231 <= w633 and not w3230;
w3232 <= w637 and not w3231;
w3233 <= w641 and not w3232;
w3234 <= w645 and not w3233;
w3235 <= w649 and not w3234;
w3236 <= w653 and not w3235;
w3237 <= w657 and not w3236;
w3238 <= w661 and not w3237;
w3239 <= w665 and not w3238;
w3240 <= w669 and not w3239;
w3241 <= w673 and not w3240;
w3242 <= w1188 and not w3241;
w3243 <= w1190 and not w3242;
w3244 <= w1451 and not w3243;
w3245 <= w682 and not w3244;
w3246 <= w686 and not w3245;
w3247 <= w690 and not w3246;
w3248 <= w694 and not w3247;
w3249 <= w698 and not w3248;
w3250 <= w702 and not w3249;
w3251 <= w706 and not w3250;
w3252 <= w710 and not w3251;
w3253 <= w714 and not w3252;
w3254 <= w718 and not w3253;
w3255 <= w722 and not w3254;
w3256 <= w726 and not w3255;
w3257 <= w730 and not w3256;
w3258 <= w734 and not w3257;
w3259 <= w738 and not w3258;
w3260 <= req(28) and not w740;
w3261 <= not w3259 and w3260;
w3262 <= not w77 and w749;
w3263 <= w754 and not w3262;
w3264 <= w758 and not w3263;
w3265 <= w762 and not w3264;
w3266 <= w766 and not w3265;
w3267 <= w770 and not w3266;
w3268 <= w774 and not w3267;
w3269 <= w778 and not w3268;
w3270 <= w782 and not w3269;
w3271 <= w786 and not w3270;
w3272 <= w790 and not w3271;
w3273 <= w794 and not w3272;
w3274 <= w798 and not w3273;
w3275 <= w802 and not w3274;
w3276 <= w806 and not w3275;
w3277 <= w810 and not w3276;
w3278 <= w814 and not w3277;
w3279 <= w818 and not w3278;
w3280 <= w822 and not w3279;
w3281 <= w826 and not w3280;
w3282 <= w830 and not w3281;
w3283 <= w834 and not w3282;
w3284 <= w838 and not w3283;
w3285 <= w842 and not w3284;
w3286 <= w846 and not w3285;
w3287 <= w850 and not w3286;
w3288 <= w854 and not w3287;
w3289 <= w858 and not w3288;
w3290 <= w862 and not w3289;
w3291 <= w866 and not w3290;
w3292 <= w870 and not w3291;
w3293 <= w874 and not w3292;
w3294 <= w878 and not w3293;
w3295 <= w882 and not w3294;
w3296 <= w886 and not w3295;
w3297 <= w890 and not w3296;
w3298 <= w894 and not w3297;
w3299 <= w898 and not w3298;
w3300 <= w902 and not w3299;
w3301 <= w906 and not w3300;
w3302 <= w910 and not w3301;
w3303 <= w914 and not w3302;
w3304 <= w918 and not w3303;
w3305 <= w922 and not w3304;
w3306 <= w926 and not w3305;
w3307 <= w930 and not w3306;
w3308 <= w934 and not w3307;
w3309 <= w938 and not w3308;
w3310 <= w942 and not w3309;
w3311 <= w946 and not w3310;
w3312 <= w950 and not w3311;
w3313 <= w954 and not w3312;
w3314 <= w958 and not w3313;
w3315 <= w962 and not w3314;
w3316 <= w966 and not w3315;
w3317 <= w970 and not w3316;
w3318 <= w974 and not w3317;
w3319 <= w978 and not w3318;
w3320 <= w982 and not w3319;
w3321 <= w986 and not w3320;
w3322 <= w990 and not w3321;
w3323 <= w994 and not w3322;
w3324 <= w998 and not w3323;
w3325 <= w1002 and not w3324;
w3326 <= w1006 and not w3325;
w3327 <= w1010 and not w3326;
w3328 <= w1277 and not w3327;
w3329 <= w6 and not w3328;
w3330 <= w10 and not w3329;
w3331 <= w14 and not w3330;
w3332 <= w18 and not w3331;
w3333 <= w22 and not w3332;
w3334 <= w26 and not w3333;
w3335 <= w30 and not w3334;
w3336 <= w34 and not w3335;
w3337 <= w38 and not w3336;
w3338 <= w42 and not w3337;
w3339 <= w46 and not w3338;
w3340 <= w50 and not w3339;
w3341 <= w54 and not w3340;
w3342 <= w58 and not w3341;
w3343 <= w62 and not w3342;
w3344 <= w66 and not w3343;
w3345 <= w70 and not w3344;
w3346 <= req(29) and not w72;
w3347 <= not w3345 and w3346;
w3348 <= w81 and not w416;
w3349 <= w86 and not w3348;
w3350 <= w90 and not w3349;
w3351 <= w94 and not w3350;
w3352 <= w98 and not w3351;
w3353 <= w102 and not w3352;
w3354 <= w106 and not w3353;
w3355 <= w110 and not w3354;
w3356 <= w114 and not w3355;
w3357 <= w118 and not w3356;
w3358 <= w122 and not w3357;
w3359 <= w126 and not w3358;
w3360 <= w130 and not w3359;
w3361 <= w134 and not w3360;
w3362 <= w138 and not w3361;
w3363 <= w142 and not w3362;
w3364 <= w146 and not w3363;
w3365 <= w150 and not w3364;
w3366 <= w154 and not w3365;
w3367 <= w158 and not w3366;
w3368 <= w162 and not w3367;
w3369 <= w166 and not w3368;
w3370 <= w170 and not w3369;
w3371 <= w174 and not w3370;
w3372 <= w178 and not w3371;
w3373 <= w182 and not w3372;
w3374 <= w186 and not w3373;
w3375 <= w190 and not w3374;
w3376 <= w194 and not w3375;
w3377 <= w198 and not w3376;
w3378 <= w202 and not w3377;
w3379 <= w206 and not w3378;
w3380 <= w210 and not w3379;
w3381 <= w214 and not w3380;
w3382 <= w218 and not w3381;
w3383 <= w222 and not w3382;
w3384 <= w226 and not w3383;
w3385 <= w230 and not w3384;
w3386 <= w234 and not w3385;
w3387 <= w238 and not w3386;
w3388 <= w242 and not w3387;
w3389 <= w246 and not w3388;
w3390 <= w250 and not w3389;
w3391 <= w254 and not w3390;
w3392 <= w258 and not w3391;
w3393 <= w262 and not w3392;
w3394 <= w266 and not w3393;
w3395 <= w270 and not w3394;
w3396 <= w274 and not w3395;
w3397 <= w278 and not w3396;
w3398 <= w282 and not w3397;
w3399 <= w286 and not w3398;
w3400 <= w290 and not w3399;
w3401 <= w294 and not w3400;
w3402 <= w298 and not w3401;
w3403 <= w302 and not w3402;
w3404 <= w306 and not w3403;
w3405 <= w310 and not w3404;
w3406 <= w314 and not w3405;
w3407 <= w318 and not w3406;
w3408 <= w322 and not w3407;
w3409 <= w326 and not w3408;
w3410 <= w330 and not w3409;
w3411 <= w334 and not w3410;
w3412 <= w1098 and not w3411;
w3413 <= w1100 and not w3412;
w3414 <= w1364 and not w3413;
w3415 <= w345 and not w3414;
w3416 <= w349 and not w3415;
w3417 <= w353 and not w3416;
w3418 <= w357 and not w3417;
w3419 <= w361 and not w3418;
w3420 <= w365 and not w3419;
w3421 <= w369 and not w3420;
w3422 <= w373 and not w3421;
w3423 <= w377 and not w3422;
w3424 <= w381 and not w3423;
w3425 <= w385 and not w3424;
w3426 <= w389 and not w3425;
w3427 <= w393 and not w3426;
w3428 <= w397 and not w3427;
w3429 <= w401 and not w3428;
w3430 <= w405 and not w3429;
w3431 <= w409 and not w3430;
w3432 <= req(30) and not w411;
w3433 <= not w3431 and w3432;
w3434 <= w420 and not w753;
w3435 <= w425 and not w3434;
w3436 <= w429 and not w3435;
w3437 <= w433 and not w3436;
w3438 <= w437 and not w3437;
w3439 <= w441 and not w3438;
w3440 <= w445 and not w3439;
w3441 <= w449 and not w3440;
w3442 <= w453 and not w3441;
w3443 <= w457 and not w3442;
w3444 <= w461 and not w3443;
w3445 <= w465 and not w3444;
w3446 <= w469 and not w3445;
w3447 <= w473 and not w3446;
w3448 <= w477 and not w3447;
w3449 <= w481 and not w3448;
w3450 <= w485 and not w3449;
w3451 <= w489 and not w3450;
w3452 <= w493 and not w3451;
w3453 <= w497 and not w3452;
w3454 <= w501 and not w3453;
w3455 <= w505 and not w3454;
w3456 <= w509 and not w3455;
w3457 <= w513 and not w3456;
w3458 <= w517 and not w3457;
w3459 <= w521 and not w3458;
w3460 <= w525 and not w3459;
w3461 <= w529 and not w3460;
w3462 <= w533 and not w3461;
w3463 <= w537 and not w3462;
w3464 <= w541 and not w3463;
w3465 <= w545 and not w3464;
w3466 <= w549 and not w3465;
w3467 <= w553 and not w3466;
w3468 <= w557 and not w3467;
w3469 <= w561 and not w3468;
w3470 <= w565 and not w3469;
w3471 <= w569 and not w3470;
w3472 <= w573 and not w3471;
w3473 <= w577 and not w3472;
w3474 <= w581 and not w3473;
w3475 <= w585 and not w3474;
w3476 <= w589 and not w3475;
w3477 <= w593 and not w3476;
w3478 <= w597 and not w3477;
w3479 <= w601 and not w3478;
w3480 <= w605 and not w3479;
w3481 <= w609 and not w3480;
w3482 <= w613 and not w3481;
w3483 <= w617 and not w3482;
w3484 <= w621 and not w3483;
w3485 <= w625 and not w3484;
w3486 <= w629 and not w3485;
w3487 <= w633 and not w3486;
w3488 <= w637 and not w3487;
w3489 <= w641 and not w3488;
w3490 <= w645 and not w3489;
w3491 <= w649 and not w3490;
w3492 <= w653 and not w3491;
w3493 <= w657 and not w3492;
w3494 <= w661 and not w3493;
w3495 <= w665 and not w3494;
w3496 <= w669 and not w3495;
w3497 <= w673 and not w3496;
w3498 <= w1188 and not w3497;
w3499 <= w1190 and not w3498;
w3500 <= w1451 and not w3499;
w3501 <= w682 and not w3500;
w3502 <= w686 and not w3501;
w3503 <= w690 and not w3502;
w3504 <= w694 and not w3503;
w3505 <= w698 and not w3504;
w3506 <= w702 and not w3505;
w3507 <= w706 and not w3506;
w3508 <= w710 and not w3507;
w3509 <= w714 and not w3508;
w3510 <= w718 and not w3509;
w3511 <= w722 and not w3510;
w3512 <= w726 and not w3511;
w3513 <= w730 and not w3512;
w3514 <= w734 and not w3513;
w3515 <= w738 and not w3514;
w3516 <= w742 and not w3515;
w3517 <= w746 and not w3516;
w3518 <= req(31) and not w748;
w3519 <= not w3517 and w3518;
w3520 <= not w85 and w757;
w3521 <= w762 and not w3520;
w3522 <= w766 and not w3521;
w3523 <= w770 and not w3522;
w3524 <= w774 and not w3523;
w3525 <= w778 and not w3524;
w3526 <= w782 and not w3525;
w3527 <= w786 and not w3526;
w3528 <= w790 and not w3527;
w3529 <= w794 and not w3528;
w3530 <= w798 and not w3529;
w3531 <= w802 and not w3530;
w3532 <= w806 and not w3531;
w3533 <= w810 and not w3532;
w3534 <= w814 and not w3533;
w3535 <= w818 and not w3534;
w3536 <= w822 and not w3535;
w3537 <= w826 and not w3536;
w3538 <= w830 and not w3537;
w3539 <= w834 and not w3538;
w3540 <= w838 and not w3539;
w3541 <= w842 and not w3540;
w3542 <= w846 and not w3541;
w3543 <= w850 and not w3542;
w3544 <= w854 and not w3543;
w3545 <= w858 and not w3544;
w3546 <= w862 and not w3545;
w3547 <= w866 and not w3546;
w3548 <= w870 and not w3547;
w3549 <= w874 and not w3548;
w3550 <= w878 and not w3549;
w3551 <= w882 and not w3550;
w3552 <= w886 and not w3551;
w3553 <= w890 and not w3552;
w3554 <= w894 and not w3553;
w3555 <= w898 and not w3554;
w3556 <= w902 and not w3555;
w3557 <= w906 and not w3556;
w3558 <= w910 and not w3557;
w3559 <= w914 and not w3558;
w3560 <= w918 and not w3559;
w3561 <= w922 and not w3560;
w3562 <= w926 and not w3561;
w3563 <= w930 and not w3562;
w3564 <= w934 and not w3563;
w3565 <= w938 and not w3564;
w3566 <= w942 and not w3565;
w3567 <= w946 and not w3566;
w3568 <= w950 and not w3567;
w3569 <= w954 and not w3568;
w3570 <= w958 and not w3569;
w3571 <= w962 and not w3570;
w3572 <= w966 and not w3571;
w3573 <= w970 and not w3572;
w3574 <= w974 and not w3573;
w3575 <= w978 and not w3574;
w3576 <= w982 and not w3575;
w3577 <= w986 and not w3576;
w3578 <= w990 and not w3577;
w3579 <= w994 and not w3578;
w3580 <= w998 and not w3579;
w3581 <= w1002 and not w3580;
w3582 <= w1006 and not w3581;
w3583 <= w1010 and not w3582;
w3584 <= w1277 and not w3583;
w3585 <= w6 and not w3584;
w3586 <= w10 and not w3585;
w3587 <= w14 and not w3586;
w3588 <= w18 and not w3587;
w3589 <= w22 and not w3588;
w3590 <= w26 and not w3589;
w3591 <= w30 and not w3590;
w3592 <= w34 and not w3591;
w3593 <= w38 and not w3592;
w3594 <= w42 and not w3593;
w3595 <= w46 and not w3594;
w3596 <= w50 and not w3595;
w3597 <= w54 and not w3596;
w3598 <= w58 and not w3597;
w3599 <= w62 and not w3598;
w3600 <= w66 and not w3599;
w3601 <= w70 and not w3600;
w3602 <= w74 and not w3601;
w3603 <= w78 and not w3602;
w3604 <= req(32) and not w80;
w3605 <= not w3603 and w3604;
w3606 <= w89 and not w424;
w3607 <= w94 and not w3606;
w3608 <= w98 and not w3607;
w3609 <= w102 and not w3608;
w3610 <= w106 and not w3609;
w3611 <= w110 and not w3610;
w3612 <= w114 and not w3611;
w3613 <= w118 and not w3612;
w3614 <= w122 and not w3613;
w3615 <= w126 and not w3614;
w3616 <= w130 and not w3615;
w3617 <= w134 and not w3616;
w3618 <= w138 and not w3617;
w3619 <= w142 and not w3618;
w3620 <= w146 and not w3619;
w3621 <= w150 and not w3620;
w3622 <= w154 and not w3621;
w3623 <= w158 and not w3622;
w3624 <= w162 and not w3623;
w3625 <= w166 and not w3624;
w3626 <= w170 and not w3625;
w3627 <= w174 and not w3626;
w3628 <= w178 and not w3627;
w3629 <= w182 and not w3628;
w3630 <= w186 and not w3629;
w3631 <= w190 and not w3630;
w3632 <= w194 and not w3631;
w3633 <= w198 and not w3632;
w3634 <= w202 and not w3633;
w3635 <= w206 and not w3634;
w3636 <= w210 and not w3635;
w3637 <= w214 and not w3636;
w3638 <= w218 and not w3637;
w3639 <= w222 and not w3638;
w3640 <= w226 and not w3639;
w3641 <= w230 and not w3640;
w3642 <= w234 and not w3641;
w3643 <= w238 and not w3642;
w3644 <= w242 and not w3643;
w3645 <= w246 and not w3644;
w3646 <= w250 and not w3645;
w3647 <= w254 and not w3646;
w3648 <= w258 and not w3647;
w3649 <= w262 and not w3648;
w3650 <= w266 and not w3649;
w3651 <= w270 and not w3650;
w3652 <= w274 and not w3651;
w3653 <= w278 and not w3652;
w3654 <= w282 and not w3653;
w3655 <= w286 and not w3654;
w3656 <= w290 and not w3655;
w3657 <= w294 and not w3656;
w3658 <= w298 and not w3657;
w3659 <= w302 and not w3658;
w3660 <= w306 and not w3659;
w3661 <= w310 and not w3660;
w3662 <= w314 and not w3661;
w3663 <= w318 and not w3662;
w3664 <= w322 and not w3663;
w3665 <= w326 and not w3664;
w3666 <= w330 and not w3665;
w3667 <= w334 and not w3666;
w3668 <= w1098 and not w3667;
w3669 <= w1100 and not w3668;
w3670 <= w1364 and not w3669;
w3671 <= w345 and not w3670;
w3672 <= w349 and not w3671;
w3673 <= w353 and not w3672;
w3674 <= w357 and not w3673;
w3675 <= w361 and not w3674;
w3676 <= w365 and not w3675;
w3677 <= w369 and not w3676;
w3678 <= w373 and not w3677;
w3679 <= w377 and not w3678;
w3680 <= w381 and not w3679;
w3681 <= w385 and not w3680;
w3682 <= w389 and not w3681;
w3683 <= w393 and not w3682;
w3684 <= w397 and not w3683;
w3685 <= w401 and not w3684;
w3686 <= w405 and not w3685;
w3687 <= w409 and not w3686;
w3688 <= w413 and not w3687;
w3689 <= w417 and not w3688;
w3690 <= req(33) and not w419;
w3691 <= not w3689 and w3690;
w3692 <= w428 and not w761;
w3693 <= w433 and not w3692;
w3694 <= w437 and not w3693;
w3695 <= w441 and not w3694;
w3696 <= w445 and not w3695;
w3697 <= w449 and not w3696;
w3698 <= w453 and not w3697;
w3699 <= w457 and not w3698;
w3700 <= w461 and not w3699;
w3701 <= w465 and not w3700;
w3702 <= w469 and not w3701;
w3703 <= w473 and not w3702;
w3704 <= w477 and not w3703;
w3705 <= w481 and not w3704;
w3706 <= w485 and not w3705;
w3707 <= w489 and not w3706;
w3708 <= w493 and not w3707;
w3709 <= w497 and not w3708;
w3710 <= w501 and not w3709;
w3711 <= w505 and not w3710;
w3712 <= w509 and not w3711;
w3713 <= w513 and not w3712;
w3714 <= w517 and not w3713;
w3715 <= w521 and not w3714;
w3716 <= w525 and not w3715;
w3717 <= w529 and not w3716;
w3718 <= w533 and not w3717;
w3719 <= w537 and not w3718;
w3720 <= w541 and not w3719;
w3721 <= w545 and not w3720;
w3722 <= w549 and not w3721;
w3723 <= w553 and not w3722;
w3724 <= w557 and not w3723;
w3725 <= w561 and not w3724;
w3726 <= w565 and not w3725;
w3727 <= w569 and not w3726;
w3728 <= w573 and not w3727;
w3729 <= w577 and not w3728;
w3730 <= w581 and not w3729;
w3731 <= w585 and not w3730;
w3732 <= w589 and not w3731;
w3733 <= w593 and not w3732;
w3734 <= w597 and not w3733;
w3735 <= w601 and not w3734;
w3736 <= w605 and not w3735;
w3737 <= w609 and not w3736;
w3738 <= w613 and not w3737;
w3739 <= w617 and not w3738;
w3740 <= w621 and not w3739;
w3741 <= w625 and not w3740;
w3742 <= w629 and not w3741;
w3743 <= w633 and not w3742;
w3744 <= w637 and not w3743;
w3745 <= w641 and not w3744;
w3746 <= w645 and not w3745;
w3747 <= w649 and not w3746;
w3748 <= w653 and not w3747;
w3749 <= w657 and not w3748;
w3750 <= w661 and not w3749;
w3751 <= w665 and not w3750;
w3752 <= w669 and not w3751;
w3753 <= w673 and not w3752;
w3754 <= w1188 and not w3753;
w3755 <= w1190 and not w3754;
w3756 <= w1451 and not w3755;
w3757 <= w682 and not w3756;
w3758 <= w686 and not w3757;
w3759 <= w690 and not w3758;
w3760 <= w694 and not w3759;
w3761 <= w698 and not w3760;
w3762 <= w702 and not w3761;
w3763 <= w706 and not w3762;
w3764 <= w710 and not w3763;
w3765 <= w714 and not w3764;
w3766 <= w718 and not w3765;
w3767 <= w722 and not w3766;
w3768 <= w726 and not w3767;
w3769 <= w730 and not w3768;
w3770 <= w734 and not w3769;
w3771 <= w738 and not w3770;
w3772 <= w742 and not w3771;
w3773 <= w746 and not w3772;
w3774 <= w750 and not w3773;
w3775 <= w754 and not w3774;
w3776 <= req(34) and not w756;
w3777 <= not w3775 and w3776;
w3778 <= not w93 and w765;
w3779 <= w770 and not w3778;
w3780 <= w774 and not w3779;
w3781 <= w778 and not w3780;
w3782 <= w782 and not w3781;
w3783 <= w786 and not w3782;
w3784 <= w790 and not w3783;
w3785 <= w794 and not w3784;
w3786 <= w798 and not w3785;
w3787 <= w802 and not w3786;
w3788 <= w806 and not w3787;
w3789 <= w810 and not w3788;
w3790 <= w814 and not w3789;
w3791 <= w818 and not w3790;
w3792 <= w822 and not w3791;
w3793 <= w826 and not w3792;
w3794 <= w830 and not w3793;
w3795 <= w834 and not w3794;
w3796 <= w838 and not w3795;
w3797 <= w842 and not w3796;
w3798 <= w846 and not w3797;
w3799 <= w850 and not w3798;
w3800 <= w854 and not w3799;
w3801 <= w858 and not w3800;
w3802 <= w862 and not w3801;
w3803 <= w866 and not w3802;
w3804 <= w870 and not w3803;
w3805 <= w874 and not w3804;
w3806 <= w878 and not w3805;
w3807 <= w882 and not w3806;
w3808 <= w886 and not w3807;
w3809 <= w890 and not w3808;
w3810 <= w894 and not w3809;
w3811 <= w898 and not w3810;
w3812 <= w902 and not w3811;
w3813 <= w906 and not w3812;
w3814 <= w910 and not w3813;
w3815 <= w914 and not w3814;
w3816 <= w918 and not w3815;
w3817 <= w922 and not w3816;
w3818 <= w926 and not w3817;
w3819 <= w930 and not w3818;
w3820 <= w934 and not w3819;
w3821 <= w938 and not w3820;
w3822 <= w942 and not w3821;
w3823 <= w946 and not w3822;
w3824 <= w950 and not w3823;
w3825 <= w954 and not w3824;
w3826 <= w958 and not w3825;
w3827 <= w962 and not w3826;
w3828 <= w966 and not w3827;
w3829 <= w970 and not w3828;
w3830 <= w974 and not w3829;
w3831 <= w978 and not w3830;
w3832 <= w982 and not w3831;
w3833 <= w986 and not w3832;
w3834 <= w990 and not w3833;
w3835 <= w994 and not w3834;
w3836 <= w998 and not w3835;
w3837 <= w1002 and not w3836;
w3838 <= w1006 and not w3837;
w3839 <= w1010 and not w3838;
w3840 <= w1277 and not w3839;
w3841 <= w6 and not w3840;
w3842 <= w10 and not w3841;
w3843 <= w14 and not w3842;
w3844 <= w18 and not w3843;
w3845 <= w22 and not w3844;
w3846 <= w26 and not w3845;
w3847 <= w30 and not w3846;
w3848 <= w34 and not w3847;
w3849 <= w38 and not w3848;
w3850 <= w42 and not w3849;
w3851 <= w46 and not w3850;
w3852 <= w50 and not w3851;
w3853 <= w54 and not w3852;
w3854 <= w58 and not w3853;
w3855 <= w62 and not w3854;
w3856 <= w66 and not w3855;
w3857 <= w70 and not w3856;
w3858 <= w74 and not w3857;
w3859 <= w78 and not w3858;
w3860 <= w82 and not w3859;
w3861 <= w86 and not w3860;
w3862 <= req(35) and not w88;
w3863 <= not w3861 and w3862;
w3864 <= w97 and not w432;
w3865 <= w102 and not w3864;
w3866 <= w106 and not w3865;
w3867 <= w110 and not w3866;
w3868 <= w114 and not w3867;
w3869 <= w118 and not w3868;
w3870 <= w122 and not w3869;
w3871 <= w126 and not w3870;
w3872 <= w130 and not w3871;
w3873 <= w134 and not w3872;
w3874 <= w138 and not w3873;
w3875 <= w142 and not w3874;
w3876 <= w146 and not w3875;
w3877 <= w150 and not w3876;
w3878 <= w154 and not w3877;
w3879 <= w158 and not w3878;
w3880 <= w162 and not w3879;
w3881 <= w166 and not w3880;
w3882 <= w170 and not w3881;
w3883 <= w174 and not w3882;
w3884 <= w178 and not w3883;
w3885 <= w182 and not w3884;
w3886 <= w186 and not w3885;
w3887 <= w190 and not w3886;
w3888 <= w194 and not w3887;
w3889 <= w198 and not w3888;
w3890 <= w202 and not w3889;
w3891 <= w206 and not w3890;
w3892 <= w210 and not w3891;
w3893 <= w214 and not w3892;
w3894 <= w218 and not w3893;
w3895 <= w222 and not w3894;
w3896 <= w226 and not w3895;
w3897 <= w230 and not w3896;
w3898 <= w234 and not w3897;
w3899 <= w238 and not w3898;
w3900 <= w242 and not w3899;
w3901 <= w246 and not w3900;
w3902 <= w250 and not w3901;
w3903 <= w254 and not w3902;
w3904 <= w258 and not w3903;
w3905 <= w262 and not w3904;
w3906 <= w266 and not w3905;
w3907 <= w270 and not w3906;
w3908 <= w274 and not w3907;
w3909 <= w278 and not w3908;
w3910 <= w282 and not w3909;
w3911 <= w286 and not w3910;
w3912 <= w290 and not w3911;
w3913 <= w294 and not w3912;
w3914 <= w298 and not w3913;
w3915 <= w302 and not w3914;
w3916 <= w306 and not w3915;
w3917 <= w310 and not w3916;
w3918 <= w314 and not w3917;
w3919 <= w318 and not w3918;
w3920 <= w322 and not w3919;
w3921 <= w326 and not w3920;
w3922 <= w330 and not w3921;
w3923 <= w334 and not w3922;
w3924 <= w1098 and not w3923;
w3925 <= w1100 and not w3924;
w3926 <= w1364 and not w3925;
w3927 <= w345 and not w3926;
w3928 <= w349 and not w3927;
w3929 <= w353 and not w3928;
w3930 <= w357 and not w3929;
w3931 <= w361 and not w3930;
w3932 <= w365 and not w3931;
w3933 <= w369 and not w3932;
w3934 <= w373 and not w3933;
w3935 <= w377 and not w3934;
w3936 <= w381 and not w3935;
w3937 <= w385 and not w3936;
w3938 <= w389 and not w3937;
w3939 <= w393 and not w3938;
w3940 <= w397 and not w3939;
w3941 <= w401 and not w3940;
w3942 <= w405 and not w3941;
w3943 <= w409 and not w3942;
w3944 <= w413 and not w3943;
w3945 <= w417 and not w3944;
w3946 <= w421 and not w3945;
w3947 <= w425 and not w3946;
w3948 <= req(36) and not w427;
w3949 <= not w3947 and w3948;
w3950 <= w436 and not w769;
w3951 <= w441 and not w3950;
w3952 <= w445 and not w3951;
w3953 <= w449 and not w3952;
w3954 <= w453 and not w3953;
w3955 <= w457 and not w3954;
w3956 <= w461 and not w3955;
w3957 <= w465 and not w3956;
w3958 <= w469 and not w3957;
w3959 <= w473 and not w3958;
w3960 <= w477 and not w3959;
w3961 <= w481 and not w3960;
w3962 <= w485 and not w3961;
w3963 <= w489 and not w3962;
w3964 <= w493 and not w3963;
w3965 <= w497 and not w3964;
w3966 <= w501 and not w3965;
w3967 <= w505 and not w3966;
w3968 <= w509 and not w3967;
w3969 <= w513 and not w3968;
w3970 <= w517 and not w3969;
w3971 <= w521 and not w3970;
w3972 <= w525 and not w3971;
w3973 <= w529 and not w3972;
w3974 <= w533 and not w3973;
w3975 <= w537 and not w3974;
w3976 <= w541 and not w3975;
w3977 <= w545 and not w3976;
w3978 <= w549 and not w3977;
w3979 <= w553 and not w3978;
w3980 <= w557 and not w3979;
w3981 <= w561 and not w3980;
w3982 <= w565 and not w3981;
w3983 <= w569 and not w3982;
w3984 <= w573 and not w3983;
w3985 <= w577 and not w3984;
w3986 <= w581 and not w3985;
w3987 <= w585 and not w3986;
w3988 <= w589 and not w3987;
w3989 <= w593 and not w3988;
w3990 <= w597 and not w3989;
w3991 <= w601 and not w3990;
w3992 <= w605 and not w3991;
w3993 <= w609 and not w3992;
w3994 <= w613 and not w3993;
w3995 <= w617 and not w3994;
w3996 <= w621 and not w3995;
w3997 <= w625 and not w3996;
w3998 <= w629 and not w3997;
w3999 <= w633 and not w3998;
w4000 <= w637 and not w3999;
w4001 <= w641 and not w4000;
w4002 <= w645 and not w4001;
w4003 <= w649 and not w4002;
w4004 <= w653 and not w4003;
w4005 <= w657 and not w4004;
w4006 <= w661 and not w4005;
w4007 <= w665 and not w4006;
w4008 <= w669 and not w4007;
w4009 <= w673 and not w4008;
w4010 <= w1188 and not w4009;
w4011 <= w1190 and not w4010;
w4012 <= w1451 and not w4011;
w4013 <= w682 and not w4012;
w4014 <= w686 and not w4013;
w4015 <= w690 and not w4014;
w4016 <= w694 and not w4015;
w4017 <= w698 and not w4016;
w4018 <= w702 and not w4017;
w4019 <= w706 and not w4018;
w4020 <= w710 and not w4019;
w4021 <= w714 and not w4020;
w4022 <= w718 and not w4021;
w4023 <= w722 and not w4022;
w4024 <= w726 and not w4023;
w4025 <= w730 and not w4024;
w4026 <= w734 and not w4025;
w4027 <= w738 and not w4026;
w4028 <= w742 and not w4027;
w4029 <= w746 and not w4028;
w4030 <= w750 and not w4029;
w4031 <= w754 and not w4030;
w4032 <= w758 and not w4031;
w4033 <= w762 and not w4032;
w4034 <= req(37) and not w764;
w4035 <= not w4033 and w4034;
w4036 <= not w101 and w773;
w4037 <= w778 and not w4036;
w4038 <= w782 and not w4037;
w4039 <= w786 and not w4038;
w4040 <= w790 and not w4039;
w4041 <= w794 and not w4040;
w4042 <= w798 and not w4041;
w4043 <= w802 and not w4042;
w4044 <= w806 and not w4043;
w4045 <= w810 and not w4044;
w4046 <= w814 and not w4045;
w4047 <= w818 and not w4046;
w4048 <= w822 and not w4047;
w4049 <= w826 and not w4048;
w4050 <= w830 and not w4049;
w4051 <= w834 and not w4050;
w4052 <= w838 and not w4051;
w4053 <= w842 and not w4052;
w4054 <= w846 and not w4053;
w4055 <= w850 and not w4054;
w4056 <= w854 and not w4055;
w4057 <= w858 and not w4056;
w4058 <= w862 and not w4057;
w4059 <= w866 and not w4058;
w4060 <= w870 and not w4059;
w4061 <= w874 and not w4060;
w4062 <= w878 and not w4061;
w4063 <= w882 and not w4062;
w4064 <= w886 and not w4063;
w4065 <= w890 and not w4064;
w4066 <= w894 and not w4065;
w4067 <= w898 and not w4066;
w4068 <= w902 and not w4067;
w4069 <= w906 and not w4068;
w4070 <= w910 and not w4069;
w4071 <= w914 and not w4070;
w4072 <= w918 and not w4071;
w4073 <= w922 and not w4072;
w4074 <= w926 and not w4073;
w4075 <= w930 and not w4074;
w4076 <= w934 and not w4075;
w4077 <= w938 and not w4076;
w4078 <= w942 and not w4077;
w4079 <= w946 and not w4078;
w4080 <= w950 and not w4079;
w4081 <= w954 and not w4080;
w4082 <= w958 and not w4081;
w4083 <= w962 and not w4082;
w4084 <= w966 and not w4083;
w4085 <= w970 and not w4084;
w4086 <= w974 and not w4085;
w4087 <= w978 and not w4086;
w4088 <= w982 and not w4087;
w4089 <= w986 and not w4088;
w4090 <= w990 and not w4089;
w4091 <= w994 and not w4090;
w4092 <= w998 and not w4091;
w4093 <= w1002 and not w4092;
w4094 <= w1006 and not w4093;
w4095 <= w1010 and not w4094;
w4096 <= w1277 and not w4095;
w4097 <= w6 and not w4096;
w4098 <= w10 and not w4097;
w4099 <= w14 and not w4098;
w4100 <= w18 and not w4099;
w4101 <= w22 and not w4100;
w4102 <= w26 and not w4101;
w4103 <= w30 and not w4102;
w4104 <= w34 and not w4103;
w4105 <= w38 and not w4104;
w4106 <= w42 and not w4105;
w4107 <= w46 and not w4106;
w4108 <= w50 and not w4107;
w4109 <= w54 and not w4108;
w4110 <= w58 and not w4109;
w4111 <= w62 and not w4110;
w4112 <= w66 and not w4111;
w4113 <= w70 and not w4112;
w4114 <= w74 and not w4113;
w4115 <= w78 and not w4114;
w4116 <= w82 and not w4115;
w4117 <= w86 and not w4116;
w4118 <= w90 and not w4117;
w4119 <= w94 and not w4118;
w4120 <= req(38) and not w96;
w4121 <= not w4119 and w4120;
w4122 <= w105 and not w440;
w4123 <= w110 and not w4122;
w4124 <= w114 and not w4123;
w4125 <= w118 and not w4124;
w4126 <= w122 and not w4125;
w4127 <= w126 and not w4126;
w4128 <= w130 and not w4127;
w4129 <= w134 and not w4128;
w4130 <= w138 and not w4129;
w4131 <= w142 and not w4130;
w4132 <= w146 and not w4131;
w4133 <= w150 and not w4132;
w4134 <= w154 and not w4133;
w4135 <= w158 and not w4134;
w4136 <= w162 and not w4135;
w4137 <= w166 and not w4136;
w4138 <= w170 and not w4137;
w4139 <= w174 and not w4138;
w4140 <= w178 and not w4139;
w4141 <= w182 and not w4140;
w4142 <= w186 and not w4141;
w4143 <= w190 and not w4142;
w4144 <= w194 and not w4143;
w4145 <= w198 and not w4144;
w4146 <= w202 and not w4145;
w4147 <= w206 and not w4146;
w4148 <= w210 and not w4147;
w4149 <= w214 and not w4148;
w4150 <= w218 and not w4149;
w4151 <= w222 and not w4150;
w4152 <= w226 and not w4151;
w4153 <= w230 and not w4152;
w4154 <= w234 and not w4153;
w4155 <= w238 and not w4154;
w4156 <= w242 and not w4155;
w4157 <= w246 and not w4156;
w4158 <= w250 and not w4157;
w4159 <= w254 and not w4158;
w4160 <= w258 and not w4159;
w4161 <= w262 and not w4160;
w4162 <= w266 and not w4161;
w4163 <= w270 and not w4162;
w4164 <= w274 and not w4163;
w4165 <= w278 and not w4164;
w4166 <= w282 and not w4165;
w4167 <= w286 and not w4166;
w4168 <= w290 and not w4167;
w4169 <= w294 and not w4168;
w4170 <= w298 and not w4169;
w4171 <= w302 and not w4170;
w4172 <= w306 and not w4171;
w4173 <= w310 and not w4172;
w4174 <= w314 and not w4173;
w4175 <= w318 and not w4174;
w4176 <= w322 and not w4175;
w4177 <= w326 and not w4176;
w4178 <= w330 and not w4177;
w4179 <= w334 and not w4178;
w4180 <= w1098 and not w4179;
w4181 <= w1100 and not w4180;
w4182 <= w1364 and not w4181;
w4183 <= w345 and not w4182;
w4184 <= w349 and not w4183;
w4185 <= w353 and not w4184;
w4186 <= w357 and not w4185;
w4187 <= w361 and not w4186;
w4188 <= w365 and not w4187;
w4189 <= w369 and not w4188;
w4190 <= w373 and not w4189;
w4191 <= w377 and not w4190;
w4192 <= w381 and not w4191;
w4193 <= w385 and not w4192;
w4194 <= w389 and not w4193;
w4195 <= w393 and not w4194;
w4196 <= w397 and not w4195;
w4197 <= w401 and not w4196;
w4198 <= w405 and not w4197;
w4199 <= w409 and not w4198;
w4200 <= w413 and not w4199;
w4201 <= w417 and not w4200;
w4202 <= w421 and not w4201;
w4203 <= w425 and not w4202;
w4204 <= w429 and not w4203;
w4205 <= w433 and not w4204;
w4206 <= req(39) and not w435;
w4207 <= not w4205 and w4206;
w4208 <= w444 and not w777;
w4209 <= w449 and not w4208;
w4210 <= w453 and not w4209;
w4211 <= w457 and not w4210;
w4212 <= w461 and not w4211;
w4213 <= w465 and not w4212;
w4214 <= w469 and not w4213;
w4215 <= w473 and not w4214;
w4216 <= w477 and not w4215;
w4217 <= w481 and not w4216;
w4218 <= w485 and not w4217;
w4219 <= w489 and not w4218;
w4220 <= w493 and not w4219;
w4221 <= w497 and not w4220;
w4222 <= w501 and not w4221;
w4223 <= w505 and not w4222;
w4224 <= w509 and not w4223;
w4225 <= w513 and not w4224;
w4226 <= w517 and not w4225;
w4227 <= w521 and not w4226;
w4228 <= w525 and not w4227;
w4229 <= w529 and not w4228;
w4230 <= w533 and not w4229;
w4231 <= w537 and not w4230;
w4232 <= w541 and not w4231;
w4233 <= w545 and not w4232;
w4234 <= w549 and not w4233;
w4235 <= w553 and not w4234;
w4236 <= w557 and not w4235;
w4237 <= w561 and not w4236;
w4238 <= w565 and not w4237;
w4239 <= w569 and not w4238;
w4240 <= w573 and not w4239;
w4241 <= w577 and not w4240;
w4242 <= w581 and not w4241;
w4243 <= w585 and not w4242;
w4244 <= w589 and not w4243;
w4245 <= w593 and not w4244;
w4246 <= w597 and not w4245;
w4247 <= w601 and not w4246;
w4248 <= w605 and not w4247;
w4249 <= w609 and not w4248;
w4250 <= w613 and not w4249;
w4251 <= w617 and not w4250;
w4252 <= w621 and not w4251;
w4253 <= w625 and not w4252;
w4254 <= w629 and not w4253;
w4255 <= w633 and not w4254;
w4256 <= w637 and not w4255;
w4257 <= w641 and not w4256;
w4258 <= w645 and not w4257;
w4259 <= w649 and not w4258;
w4260 <= w653 and not w4259;
w4261 <= w657 and not w4260;
w4262 <= w661 and not w4261;
w4263 <= w665 and not w4262;
w4264 <= w669 and not w4263;
w4265 <= w673 and not w4264;
w4266 <= w1188 and not w4265;
w4267 <= w1190 and not w4266;
w4268 <= w1451 and not w4267;
w4269 <= w682 and not w4268;
w4270 <= w686 and not w4269;
w4271 <= w690 and not w4270;
w4272 <= w694 and not w4271;
w4273 <= w698 and not w4272;
w4274 <= w702 and not w4273;
w4275 <= w706 and not w4274;
w4276 <= w710 and not w4275;
w4277 <= w714 and not w4276;
w4278 <= w718 and not w4277;
w4279 <= w722 and not w4278;
w4280 <= w726 and not w4279;
w4281 <= w730 and not w4280;
w4282 <= w734 and not w4281;
w4283 <= w738 and not w4282;
w4284 <= w742 and not w4283;
w4285 <= w746 and not w4284;
w4286 <= w750 and not w4285;
w4287 <= w754 and not w4286;
w4288 <= w758 and not w4287;
w4289 <= w762 and not w4288;
w4290 <= w766 and not w4289;
w4291 <= w770 and not w4290;
w4292 <= req(40) and not w772;
w4293 <= not w4291 and w4292;
w4294 <= not w109 and w781;
w4295 <= w786 and not w4294;
w4296 <= w790 and not w4295;
w4297 <= w794 and not w4296;
w4298 <= w798 and not w4297;
w4299 <= w802 and not w4298;
w4300 <= w806 and not w4299;
w4301 <= w810 and not w4300;
w4302 <= w814 and not w4301;
w4303 <= w818 and not w4302;
w4304 <= w822 and not w4303;
w4305 <= w826 and not w4304;
w4306 <= w830 and not w4305;
w4307 <= w834 and not w4306;
w4308 <= w838 and not w4307;
w4309 <= w842 and not w4308;
w4310 <= w846 and not w4309;
w4311 <= w850 and not w4310;
w4312 <= w854 and not w4311;
w4313 <= w858 and not w4312;
w4314 <= w862 and not w4313;
w4315 <= w866 and not w4314;
w4316 <= w870 and not w4315;
w4317 <= w874 and not w4316;
w4318 <= w878 and not w4317;
w4319 <= w882 and not w4318;
w4320 <= w886 and not w4319;
w4321 <= w890 and not w4320;
w4322 <= w894 and not w4321;
w4323 <= w898 and not w4322;
w4324 <= w902 and not w4323;
w4325 <= w906 and not w4324;
w4326 <= w910 and not w4325;
w4327 <= w914 and not w4326;
w4328 <= w918 and not w4327;
w4329 <= w922 and not w4328;
w4330 <= w926 and not w4329;
w4331 <= w930 and not w4330;
w4332 <= w934 and not w4331;
w4333 <= w938 and not w4332;
w4334 <= w942 and not w4333;
w4335 <= w946 and not w4334;
w4336 <= w950 and not w4335;
w4337 <= w954 and not w4336;
w4338 <= w958 and not w4337;
w4339 <= w962 and not w4338;
w4340 <= w966 and not w4339;
w4341 <= w970 and not w4340;
w4342 <= w974 and not w4341;
w4343 <= w978 and not w4342;
w4344 <= w982 and not w4343;
w4345 <= w986 and not w4344;
w4346 <= w990 and not w4345;
w4347 <= w994 and not w4346;
w4348 <= w998 and not w4347;
w4349 <= w1002 and not w4348;
w4350 <= w1006 and not w4349;
w4351 <= w1010 and not w4350;
w4352 <= w1277 and not w4351;
w4353 <= w6 and not w4352;
w4354 <= w10 and not w4353;
w4355 <= w14 and not w4354;
w4356 <= w18 and not w4355;
w4357 <= w22 and not w4356;
w4358 <= w26 and not w4357;
w4359 <= w30 and not w4358;
w4360 <= w34 and not w4359;
w4361 <= w38 and not w4360;
w4362 <= w42 and not w4361;
w4363 <= w46 and not w4362;
w4364 <= w50 and not w4363;
w4365 <= w54 and not w4364;
w4366 <= w58 and not w4365;
w4367 <= w62 and not w4366;
w4368 <= w66 and not w4367;
w4369 <= w70 and not w4368;
w4370 <= w74 and not w4369;
w4371 <= w78 and not w4370;
w4372 <= w82 and not w4371;
w4373 <= w86 and not w4372;
w4374 <= w90 and not w4373;
w4375 <= w94 and not w4374;
w4376 <= w98 and not w4375;
w4377 <= w102 and not w4376;
w4378 <= req(41) and not w104;
w4379 <= not w4377 and w4378;
w4380 <= w113 and not w448;
w4381 <= w118 and not w4380;
w4382 <= w122 and not w4381;
w4383 <= w126 and not w4382;
w4384 <= w130 and not w4383;
w4385 <= w134 and not w4384;
w4386 <= w138 and not w4385;
w4387 <= w142 and not w4386;
w4388 <= w146 and not w4387;
w4389 <= w150 and not w4388;
w4390 <= w154 and not w4389;
w4391 <= w158 and not w4390;
w4392 <= w162 and not w4391;
w4393 <= w166 and not w4392;
w4394 <= w170 and not w4393;
w4395 <= w174 and not w4394;
w4396 <= w178 and not w4395;
w4397 <= w182 and not w4396;
w4398 <= w186 and not w4397;
w4399 <= w190 and not w4398;
w4400 <= w194 and not w4399;
w4401 <= w198 and not w4400;
w4402 <= w202 and not w4401;
w4403 <= w206 and not w4402;
w4404 <= w210 and not w4403;
w4405 <= w214 and not w4404;
w4406 <= w218 and not w4405;
w4407 <= w222 and not w4406;
w4408 <= w226 and not w4407;
w4409 <= w230 and not w4408;
w4410 <= w234 and not w4409;
w4411 <= w238 and not w4410;
w4412 <= w242 and not w4411;
w4413 <= w246 and not w4412;
w4414 <= w250 and not w4413;
w4415 <= w254 and not w4414;
w4416 <= w258 and not w4415;
w4417 <= w262 and not w4416;
w4418 <= w266 and not w4417;
w4419 <= w270 and not w4418;
w4420 <= w274 and not w4419;
w4421 <= w278 and not w4420;
w4422 <= w282 and not w4421;
w4423 <= w286 and not w4422;
w4424 <= w290 and not w4423;
w4425 <= w294 and not w4424;
w4426 <= w298 and not w4425;
w4427 <= w302 and not w4426;
w4428 <= w306 and not w4427;
w4429 <= w310 and not w4428;
w4430 <= w314 and not w4429;
w4431 <= w318 and not w4430;
w4432 <= w322 and not w4431;
w4433 <= w326 and not w4432;
w4434 <= w330 and not w4433;
w4435 <= w334 and not w4434;
w4436 <= w1098 and not w4435;
w4437 <= w1100 and not w4436;
w4438 <= w1364 and not w4437;
w4439 <= w345 and not w4438;
w4440 <= w349 and not w4439;
w4441 <= w353 and not w4440;
w4442 <= w357 and not w4441;
w4443 <= w361 and not w4442;
w4444 <= w365 and not w4443;
w4445 <= w369 and not w4444;
w4446 <= w373 and not w4445;
w4447 <= w377 and not w4446;
w4448 <= w381 and not w4447;
w4449 <= w385 and not w4448;
w4450 <= w389 and not w4449;
w4451 <= w393 and not w4450;
w4452 <= w397 and not w4451;
w4453 <= w401 and not w4452;
w4454 <= w405 and not w4453;
w4455 <= w409 and not w4454;
w4456 <= w413 and not w4455;
w4457 <= w417 and not w4456;
w4458 <= w421 and not w4457;
w4459 <= w425 and not w4458;
w4460 <= w429 and not w4459;
w4461 <= w433 and not w4460;
w4462 <= w437 and not w4461;
w4463 <= w441 and not w4462;
w4464 <= req(42) and not w443;
w4465 <= not w4463 and w4464;
w4466 <= w452 and not w785;
w4467 <= w457 and not w4466;
w4468 <= w461 and not w4467;
w4469 <= w465 and not w4468;
w4470 <= w469 and not w4469;
w4471 <= w473 and not w4470;
w4472 <= w477 and not w4471;
w4473 <= w481 and not w4472;
w4474 <= w485 and not w4473;
w4475 <= w489 and not w4474;
w4476 <= w493 and not w4475;
w4477 <= w497 and not w4476;
w4478 <= w501 and not w4477;
w4479 <= w505 and not w4478;
w4480 <= w509 and not w4479;
w4481 <= w513 and not w4480;
w4482 <= w517 and not w4481;
w4483 <= w521 and not w4482;
w4484 <= w525 and not w4483;
w4485 <= w529 and not w4484;
w4486 <= w533 and not w4485;
w4487 <= w537 and not w4486;
w4488 <= w541 and not w4487;
w4489 <= w545 and not w4488;
w4490 <= w549 and not w4489;
w4491 <= w553 and not w4490;
w4492 <= w557 and not w4491;
w4493 <= w561 and not w4492;
w4494 <= w565 and not w4493;
w4495 <= w569 and not w4494;
w4496 <= w573 and not w4495;
w4497 <= w577 and not w4496;
w4498 <= w581 and not w4497;
w4499 <= w585 and not w4498;
w4500 <= w589 and not w4499;
w4501 <= w593 and not w4500;
w4502 <= w597 and not w4501;
w4503 <= w601 and not w4502;
w4504 <= w605 and not w4503;
w4505 <= w609 and not w4504;
w4506 <= w613 and not w4505;
w4507 <= w617 and not w4506;
w4508 <= w621 and not w4507;
w4509 <= w625 and not w4508;
w4510 <= w629 and not w4509;
w4511 <= w633 and not w4510;
w4512 <= w637 and not w4511;
w4513 <= w641 and not w4512;
w4514 <= w645 and not w4513;
w4515 <= w649 and not w4514;
w4516 <= w653 and not w4515;
w4517 <= w657 and not w4516;
w4518 <= w661 and not w4517;
w4519 <= w665 and not w4518;
w4520 <= w669 and not w4519;
w4521 <= w673 and not w4520;
w4522 <= w1188 and not w4521;
w4523 <= w1190 and not w4522;
w4524 <= w1451 and not w4523;
w4525 <= w682 and not w4524;
w4526 <= w686 and not w4525;
w4527 <= w690 and not w4526;
w4528 <= w694 and not w4527;
w4529 <= w698 and not w4528;
w4530 <= w702 and not w4529;
w4531 <= w706 and not w4530;
w4532 <= w710 and not w4531;
w4533 <= w714 and not w4532;
w4534 <= w718 and not w4533;
w4535 <= w722 and not w4534;
w4536 <= w726 and not w4535;
w4537 <= w730 and not w4536;
w4538 <= w734 and not w4537;
w4539 <= w738 and not w4538;
w4540 <= w742 and not w4539;
w4541 <= w746 and not w4540;
w4542 <= w750 and not w4541;
w4543 <= w754 and not w4542;
w4544 <= w758 and not w4543;
w4545 <= w762 and not w4544;
w4546 <= w766 and not w4545;
w4547 <= w770 and not w4546;
w4548 <= w774 and not w4547;
w4549 <= w778 and not w4548;
w4550 <= req(43) and not w780;
w4551 <= not w4549 and w4550;
w4552 <= not w117 and w789;
w4553 <= w794 and not w4552;
w4554 <= w798 and not w4553;
w4555 <= w802 and not w4554;
w4556 <= w806 and not w4555;
w4557 <= w810 and not w4556;
w4558 <= w814 and not w4557;
w4559 <= w818 and not w4558;
w4560 <= w822 and not w4559;
w4561 <= w826 and not w4560;
w4562 <= w830 and not w4561;
w4563 <= w834 and not w4562;
w4564 <= w838 and not w4563;
w4565 <= w842 and not w4564;
w4566 <= w846 and not w4565;
w4567 <= w850 and not w4566;
w4568 <= w854 and not w4567;
w4569 <= w858 and not w4568;
w4570 <= w862 and not w4569;
w4571 <= w866 and not w4570;
w4572 <= w870 and not w4571;
w4573 <= w874 and not w4572;
w4574 <= w878 and not w4573;
w4575 <= w882 and not w4574;
w4576 <= w886 and not w4575;
w4577 <= w890 and not w4576;
w4578 <= w894 and not w4577;
w4579 <= w898 and not w4578;
w4580 <= w902 and not w4579;
w4581 <= w906 and not w4580;
w4582 <= w910 and not w4581;
w4583 <= w914 and not w4582;
w4584 <= w918 and not w4583;
w4585 <= w922 and not w4584;
w4586 <= w926 and not w4585;
w4587 <= w930 and not w4586;
w4588 <= w934 and not w4587;
w4589 <= w938 and not w4588;
w4590 <= w942 and not w4589;
w4591 <= w946 and not w4590;
w4592 <= w950 and not w4591;
w4593 <= w954 and not w4592;
w4594 <= w958 and not w4593;
w4595 <= w962 and not w4594;
w4596 <= w966 and not w4595;
w4597 <= w970 and not w4596;
w4598 <= w974 and not w4597;
w4599 <= w978 and not w4598;
w4600 <= w982 and not w4599;
w4601 <= w986 and not w4600;
w4602 <= w990 and not w4601;
w4603 <= w994 and not w4602;
w4604 <= w998 and not w4603;
w4605 <= w1002 and not w4604;
w4606 <= w1006 and not w4605;
w4607 <= w1010 and not w4606;
w4608 <= w1277 and not w4607;
w4609 <= w6 and not w4608;
w4610 <= w10 and not w4609;
w4611 <= w14 and not w4610;
w4612 <= w18 and not w4611;
w4613 <= w22 and not w4612;
w4614 <= w26 and not w4613;
w4615 <= w30 and not w4614;
w4616 <= w34 and not w4615;
w4617 <= w38 and not w4616;
w4618 <= w42 and not w4617;
w4619 <= w46 and not w4618;
w4620 <= w50 and not w4619;
w4621 <= w54 and not w4620;
w4622 <= w58 and not w4621;
w4623 <= w62 and not w4622;
w4624 <= w66 and not w4623;
w4625 <= w70 and not w4624;
w4626 <= w74 and not w4625;
w4627 <= w78 and not w4626;
w4628 <= w82 and not w4627;
w4629 <= w86 and not w4628;
w4630 <= w90 and not w4629;
w4631 <= w94 and not w4630;
w4632 <= w98 and not w4631;
w4633 <= w102 and not w4632;
w4634 <= w106 and not w4633;
w4635 <= w110 and not w4634;
w4636 <= req(44) and not w112;
w4637 <= not w4635 and w4636;
w4638 <= w121 and not w456;
w4639 <= w126 and not w4638;
w4640 <= w130 and not w4639;
w4641 <= w134 and not w4640;
w4642 <= w138 and not w4641;
w4643 <= w142 and not w4642;
w4644 <= w146 and not w4643;
w4645 <= w150 and not w4644;
w4646 <= w154 and not w4645;
w4647 <= w158 and not w4646;
w4648 <= w162 and not w4647;
w4649 <= w166 and not w4648;
w4650 <= w170 and not w4649;
w4651 <= w174 and not w4650;
w4652 <= w178 and not w4651;
w4653 <= w182 and not w4652;
w4654 <= w186 and not w4653;
w4655 <= w190 and not w4654;
w4656 <= w194 and not w4655;
w4657 <= w198 and not w4656;
w4658 <= w202 and not w4657;
w4659 <= w206 and not w4658;
w4660 <= w210 and not w4659;
w4661 <= w214 and not w4660;
w4662 <= w218 and not w4661;
w4663 <= w222 and not w4662;
w4664 <= w226 and not w4663;
w4665 <= w230 and not w4664;
w4666 <= w234 and not w4665;
w4667 <= w238 and not w4666;
w4668 <= w242 and not w4667;
w4669 <= w246 and not w4668;
w4670 <= w250 and not w4669;
w4671 <= w254 and not w4670;
w4672 <= w258 and not w4671;
w4673 <= w262 and not w4672;
w4674 <= w266 and not w4673;
w4675 <= w270 and not w4674;
w4676 <= w274 and not w4675;
w4677 <= w278 and not w4676;
w4678 <= w282 and not w4677;
w4679 <= w286 and not w4678;
w4680 <= w290 and not w4679;
w4681 <= w294 and not w4680;
w4682 <= w298 and not w4681;
w4683 <= w302 and not w4682;
w4684 <= w306 and not w4683;
w4685 <= w310 and not w4684;
w4686 <= w314 and not w4685;
w4687 <= w318 and not w4686;
w4688 <= w322 and not w4687;
w4689 <= w326 and not w4688;
w4690 <= w330 and not w4689;
w4691 <= w334 and not w4690;
w4692 <= w1098 and not w4691;
w4693 <= w1100 and not w4692;
w4694 <= w1364 and not w4693;
w4695 <= w345 and not w4694;
w4696 <= w349 and not w4695;
w4697 <= w353 and not w4696;
w4698 <= w357 and not w4697;
w4699 <= w361 and not w4698;
w4700 <= w365 and not w4699;
w4701 <= w369 and not w4700;
w4702 <= w373 and not w4701;
w4703 <= w377 and not w4702;
w4704 <= w381 and not w4703;
w4705 <= w385 and not w4704;
w4706 <= w389 and not w4705;
w4707 <= w393 and not w4706;
w4708 <= w397 and not w4707;
w4709 <= w401 and not w4708;
w4710 <= w405 and not w4709;
w4711 <= w409 and not w4710;
w4712 <= w413 and not w4711;
w4713 <= w417 and not w4712;
w4714 <= w421 and not w4713;
w4715 <= w425 and not w4714;
w4716 <= w429 and not w4715;
w4717 <= w433 and not w4716;
w4718 <= w437 and not w4717;
w4719 <= w441 and not w4718;
w4720 <= w445 and not w4719;
w4721 <= w449 and not w4720;
w4722 <= req(45) and not w451;
w4723 <= not w4721 and w4722;
w4724 <= w460 and not w793;
w4725 <= w465 and not w4724;
w4726 <= w469 and not w4725;
w4727 <= w473 and not w4726;
w4728 <= w477 and not w4727;
w4729 <= w481 and not w4728;
w4730 <= w485 and not w4729;
w4731 <= w489 and not w4730;
w4732 <= w493 and not w4731;
w4733 <= w497 and not w4732;
w4734 <= w501 and not w4733;
w4735 <= w505 and not w4734;
w4736 <= w509 and not w4735;
w4737 <= w513 and not w4736;
w4738 <= w517 and not w4737;
w4739 <= w521 and not w4738;
w4740 <= w525 and not w4739;
w4741 <= w529 and not w4740;
w4742 <= w533 and not w4741;
w4743 <= w537 and not w4742;
w4744 <= w541 and not w4743;
w4745 <= w545 and not w4744;
w4746 <= w549 and not w4745;
w4747 <= w553 and not w4746;
w4748 <= w557 and not w4747;
w4749 <= w561 and not w4748;
w4750 <= w565 and not w4749;
w4751 <= w569 and not w4750;
w4752 <= w573 and not w4751;
w4753 <= w577 and not w4752;
w4754 <= w581 and not w4753;
w4755 <= w585 and not w4754;
w4756 <= w589 and not w4755;
w4757 <= w593 and not w4756;
w4758 <= w597 and not w4757;
w4759 <= w601 and not w4758;
w4760 <= w605 and not w4759;
w4761 <= w609 and not w4760;
w4762 <= w613 and not w4761;
w4763 <= w617 and not w4762;
w4764 <= w621 and not w4763;
w4765 <= w625 and not w4764;
w4766 <= w629 and not w4765;
w4767 <= w633 and not w4766;
w4768 <= w637 and not w4767;
w4769 <= w641 and not w4768;
w4770 <= w645 and not w4769;
w4771 <= w649 and not w4770;
w4772 <= w653 and not w4771;
w4773 <= w657 and not w4772;
w4774 <= w661 and not w4773;
w4775 <= w665 and not w4774;
w4776 <= w669 and not w4775;
w4777 <= w673 and not w4776;
w4778 <= w1188 and not w4777;
w4779 <= w1190 and not w4778;
w4780 <= w1451 and not w4779;
w4781 <= w682 and not w4780;
w4782 <= w686 and not w4781;
w4783 <= w690 and not w4782;
w4784 <= w694 and not w4783;
w4785 <= w698 and not w4784;
w4786 <= w702 and not w4785;
w4787 <= w706 and not w4786;
w4788 <= w710 and not w4787;
w4789 <= w714 and not w4788;
w4790 <= w718 and not w4789;
w4791 <= w722 and not w4790;
w4792 <= w726 and not w4791;
w4793 <= w730 and not w4792;
w4794 <= w734 and not w4793;
w4795 <= w738 and not w4794;
w4796 <= w742 and not w4795;
w4797 <= w746 and not w4796;
w4798 <= w750 and not w4797;
w4799 <= w754 and not w4798;
w4800 <= w758 and not w4799;
w4801 <= w762 and not w4800;
w4802 <= w766 and not w4801;
w4803 <= w770 and not w4802;
w4804 <= w774 and not w4803;
w4805 <= w778 and not w4804;
w4806 <= w782 and not w4805;
w4807 <= w786 and not w4806;
w4808 <= req(46) and not w788;
w4809 <= not w4807 and w4808;
w4810 <= not w125 and w797;
w4811 <= w802 and not w4810;
w4812 <= w806 and not w4811;
w4813 <= w810 and not w4812;
w4814 <= w814 and not w4813;
w4815 <= w818 and not w4814;
w4816 <= w822 and not w4815;
w4817 <= w826 and not w4816;
w4818 <= w830 and not w4817;
w4819 <= w834 and not w4818;
w4820 <= w838 and not w4819;
w4821 <= w842 and not w4820;
w4822 <= w846 and not w4821;
w4823 <= w850 and not w4822;
w4824 <= w854 and not w4823;
w4825 <= w858 and not w4824;
w4826 <= w862 and not w4825;
w4827 <= w866 and not w4826;
w4828 <= w870 and not w4827;
w4829 <= w874 and not w4828;
w4830 <= w878 and not w4829;
w4831 <= w882 and not w4830;
w4832 <= w886 and not w4831;
w4833 <= w890 and not w4832;
w4834 <= w894 and not w4833;
w4835 <= w898 and not w4834;
w4836 <= w902 and not w4835;
w4837 <= w906 and not w4836;
w4838 <= w910 and not w4837;
w4839 <= w914 and not w4838;
w4840 <= w918 and not w4839;
w4841 <= w922 and not w4840;
w4842 <= w926 and not w4841;
w4843 <= w930 and not w4842;
w4844 <= w934 and not w4843;
w4845 <= w938 and not w4844;
w4846 <= w942 and not w4845;
w4847 <= w946 and not w4846;
w4848 <= w950 and not w4847;
w4849 <= w954 and not w4848;
w4850 <= w958 and not w4849;
w4851 <= w962 and not w4850;
w4852 <= w966 and not w4851;
w4853 <= w970 and not w4852;
w4854 <= w974 and not w4853;
w4855 <= w978 and not w4854;
w4856 <= w982 and not w4855;
w4857 <= w986 and not w4856;
w4858 <= w990 and not w4857;
w4859 <= w994 and not w4858;
w4860 <= w998 and not w4859;
w4861 <= w1002 and not w4860;
w4862 <= w1006 and not w4861;
w4863 <= w1010 and not w4862;
w4864 <= w1277 and not w4863;
w4865 <= w6 and not w4864;
w4866 <= w10 and not w4865;
w4867 <= w14 and not w4866;
w4868 <= w18 and not w4867;
w4869 <= w22 and not w4868;
w4870 <= w26 and not w4869;
w4871 <= w30 and not w4870;
w4872 <= w34 and not w4871;
w4873 <= w38 and not w4872;
w4874 <= w42 and not w4873;
w4875 <= w46 and not w4874;
w4876 <= w50 and not w4875;
w4877 <= w54 and not w4876;
w4878 <= w58 and not w4877;
w4879 <= w62 and not w4878;
w4880 <= w66 and not w4879;
w4881 <= w70 and not w4880;
w4882 <= w74 and not w4881;
w4883 <= w78 and not w4882;
w4884 <= w82 and not w4883;
w4885 <= w86 and not w4884;
w4886 <= w90 and not w4885;
w4887 <= w94 and not w4886;
w4888 <= w98 and not w4887;
w4889 <= w102 and not w4888;
w4890 <= w106 and not w4889;
w4891 <= w110 and not w4890;
w4892 <= w114 and not w4891;
w4893 <= w118 and not w4892;
w4894 <= req(47) and not w120;
w4895 <= not w4893 and w4894;
w4896 <= w129 and not w464;
w4897 <= w134 and not w4896;
w4898 <= w138 and not w4897;
w4899 <= w142 and not w4898;
w4900 <= w146 and not w4899;
w4901 <= w150 and not w4900;
w4902 <= w154 and not w4901;
w4903 <= w158 and not w4902;
w4904 <= w162 and not w4903;
w4905 <= w166 and not w4904;
w4906 <= w170 and not w4905;
w4907 <= w174 and not w4906;
w4908 <= w178 and not w4907;
w4909 <= w182 and not w4908;
w4910 <= w186 and not w4909;
w4911 <= w190 and not w4910;
w4912 <= w194 and not w4911;
w4913 <= w198 and not w4912;
w4914 <= w202 and not w4913;
w4915 <= w206 and not w4914;
w4916 <= w210 and not w4915;
w4917 <= w214 and not w4916;
w4918 <= w218 and not w4917;
w4919 <= w222 and not w4918;
w4920 <= w226 and not w4919;
w4921 <= w230 and not w4920;
w4922 <= w234 and not w4921;
w4923 <= w238 and not w4922;
w4924 <= w242 and not w4923;
w4925 <= w246 and not w4924;
w4926 <= w250 and not w4925;
w4927 <= w254 and not w4926;
w4928 <= w258 and not w4927;
w4929 <= w262 and not w4928;
w4930 <= w266 and not w4929;
w4931 <= w270 and not w4930;
w4932 <= w274 and not w4931;
w4933 <= w278 and not w4932;
w4934 <= w282 and not w4933;
w4935 <= w286 and not w4934;
w4936 <= w290 and not w4935;
w4937 <= w294 and not w4936;
w4938 <= w298 and not w4937;
w4939 <= w302 and not w4938;
w4940 <= w306 and not w4939;
w4941 <= w310 and not w4940;
w4942 <= w314 and not w4941;
w4943 <= w318 and not w4942;
w4944 <= w322 and not w4943;
w4945 <= w326 and not w4944;
w4946 <= w330 and not w4945;
w4947 <= w334 and not w4946;
w4948 <= w1098 and not w4947;
w4949 <= w1100 and not w4948;
w4950 <= w1364 and not w4949;
w4951 <= w345 and not w4950;
w4952 <= w349 and not w4951;
w4953 <= w353 and not w4952;
w4954 <= w357 and not w4953;
w4955 <= w361 and not w4954;
w4956 <= w365 and not w4955;
w4957 <= w369 and not w4956;
w4958 <= w373 and not w4957;
w4959 <= w377 and not w4958;
w4960 <= w381 and not w4959;
w4961 <= w385 and not w4960;
w4962 <= w389 and not w4961;
w4963 <= w393 and not w4962;
w4964 <= w397 and not w4963;
w4965 <= w401 and not w4964;
w4966 <= w405 and not w4965;
w4967 <= w409 and not w4966;
w4968 <= w413 and not w4967;
w4969 <= w417 and not w4968;
w4970 <= w421 and not w4969;
w4971 <= w425 and not w4970;
w4972 <= w429 and not w4971;
w4973 <= w433 and not w4972;
w4974 <= w437 and not w4973;
w4975 <= w441 and not w4974;
w4976 <= w445 and not w4975;
w4977 <= w449 and not w4976;
w4978 <= w453 and not w4977;
w4979 <= w457 and not w4978;
w4980 <= req(48) and not w459;
w4981 <= not w4979 and w4980;
w4982 <= w468 and not w801;
w4983 <= w473 and not w4982;
w4984 <= w477 and not w4983;
w4985 <= w481 and not w4984;
w4986 <= w485 and not w4985;
w4987 <= w489 and not w4986;
w4988 <= w493 and not w4987;
w4989 <= w497 and not w4988;
w4990 <= w501 and not w4989;
w4991 <= w505 and not w4990;
w4992 <= w509 and not w4991;
w4993 <= w513 and not w4992;
w4994 <= w517 and not w4993;
w4995 <= w521 and not w4994;
w4996 <= w525 and not w4995;
w4997 <= w529 and not w4996;
w4998 <= w533 and not w4997;
w4999 <= w537 and not w4998;
w5000 <= w541 and not w4999;
w5001 <= w545 and not w5000;
w5002 <= w549 and not w5001;
w5003 <= w553 and not w5002;
w5004 <= w557 and not w5003;
w5005 <= w561 and not w5004;
w5006 <= w565 and not w5005;
w5007 <= w569 and not w5006;
w5008 <= w573 and not w5007;
w5009 <= w577 and not w5008;
w5010 <= w581 and not w5009;
w5011 <= w585 and not w5010;
w5012 <= w589 and not w5011;
w5013 <= w593 and not w5012;
w5014 <= w597 and not w5013;
w5015 <= w601 and not w5014;
w5016 <= w605 and not w5015;
w5017 <= w609 and not w5016;
w5018 <= w613 and not w5017;
w5019 <= w617 and not w5018;
w5020 <= w621 and not w5019;
w5021 <= w625 and not w5020;
w5022 <= w629 and not w5021;
w5023 <= w633 and not w5022;
w5024 <= w637 and not w5023;
w5025 <= w641 and not w5024;
w5026 <= w645 and not w5025;
w5027 <= w649 and not w5026;
w5028 <= w653 and not w5027;
w5029 <= w657 and not w5028;
w5030 <= w661 and not w5029;
w5031 <= w665 and not w5030;
w5032 <= w669 and not w5031;
w5033 <= w673 and not w5032;
w5034 <= w1188 and not w5033;
w5035 <= w1190 and not w5034;
w5036 <= w1451 and not w5035;
w5037 <= w682 and not w5036;
w5038 <= w686 and not w5037;
w5039 <= w690 and not w5038;
w5040 <= w694 and not w5039;
w5041 <= w698 and not w5040;
w5042 <= w702 and not w5041;
w5043 <= w706 and not w5042;
w5044 <= w710 and not w5043;
w5045 <= w714 and not w5044;
w5046 <= w718 and not w5045;
w5047 <= w722 and not w5046;
w5048 <= w726 and not w5047;
w5049 <= w730 and not w5048;
w5050 <= w734 and not w5049;
w5051 <= w738 and not w5050;
w5052 <= w742 and not w5051;
w5053 <= w746 and not w5052;
w5054 <= w750 and not w5053;
w5055 <= w754 and not w5054;
w5056 <= w758 and not w5055;
w5057 <= w762 and not w5056;
w5058 <= w766 and not w5057;
w5059 <= w770 and not w5058;
w5060 <= w774 and not w5059;
w5061 <= w778 and not w5060;
w5062 <= w782 and not w5061;
w5063 <= w786 and not w5062;
w5064 <= w790 and not w5063;
w5065 <= w794 and not w5064;
w5066 <= req(49) and not w796;
w5067 <= not w5065 and w5066;
w5068 <= not w133 and w805;
w5069 <= w810 and not w5068;
w5070 <= w814 and not w5069;
w5071 <= w818 and not w5070;
w5072 <= w822 and not w5071;
w5073 <= w826 and not w5072;
w5074 <= w830 and not w5073;
w5075 <= w834 and not w5074;
w5076 <= w838 and not w5075;
w5077 <= w842 and not w5076;
w5078 <= w846 and not w5077;
w5079 <= w850 and not w5078;
w5080 <= w854 and not w5079;
w5081 <= w858 and not w5080;
w5082 <= w862 and not w5081;
w5083 <= w866 and not w5082;
w5084 <= w870 and not w5083;
w5085 <= w874 and not w5084;
w5086 <= w878 and not w5085;
w5087 <= w882 and not w5086;
w5088 <= w886 and not w5087;
w5089 <= w890 and not w5088;
w5090 <= w894 and not w5089;
w5091 <= w898 and not w5090;
w5092 <= w902 and not w5091;
w5093 <= w906 and not w5092;
w5094 <= w910 and not w5093;
w5095 <= w914 and not w5094;
w5096 <= w918 and not w5095;
w5097 <= w922 and not w5096;
w5098 <= w926 and not w5097;
w5099 <= w930 and not w5098;
w5100 <= w934 and not w5099;
w5101 <= w938 and not w5100;
w5102 <= w942 and not w5101;
w5103 <= w946 and not w5102;
w5104 <= w950 and not w5103;
w5105 <= w954 and not w5104;
w5106 <= w958 and not w5105;
w5107 <= w962 and not w5106;
w5108 <= w966 and not w5107;
w5109 <= w970 and not w5108;
w5110 <= w974 and not w5109;
w5111 <= w978 and not w5110;
w5112 <= w982 and not w5111;
w5113 <= w986 and not w5112;
w5114 <= w990 and not w5113;
w5115 <= w994 and not w5114;
w5116 <= w998 and not w5115;
w5117 <= w1002 and not w5116;
w5118 <= w1006 and not w5117;
w5119 <= w1010 and not w5118;
w5120 <= w1277 and not w5119;
w5121 <= w6 and not w5120;
w5122 <= w10 and not w5121;
w5123 <= w14 and not w5122;
w5124 <= w18 and not w5123;
w5125 <= w22 and not w5124;
w5126 <= w26 and not w5125;
w5127 <= w30 and not w5126;
w5128 <= w34 and not w5127;
w5129 <= w38 and not w5128;
w5130 <= w42 and not w5129;
w5131 <= w46 and not w5130;
w5132 <= w50 and not w5131;
w5133 <= w54 and not w5132;
w5134 <= w58 and not w5133;
w5135 <= w62 and not w5134;
w5136 <= w66 and not w5135;
w5137 <= w70 and not w5136;
w5138 <= w74 and not w5137;
w5139 <= w78 and not w5138;
w5140 <= w82 and not w5139;
w5141 <= w86 and not w5140;
w5142 <= w90 and not w5141;
w5143 <= w94 and not w5142;
w5144 <= w98 and not w5143;
w5145 <= w102 and not w5144;
w5146 <= w106 and not w5145;
w5147 <= w110 and not w5146;
w5148 <= w114 and not w5147;
w5149 <= w118 and not w5148;
w5150 <= w122 and not w5149;
w5151 <= w126 and not w5150;
w5152 <= req(50) and not w128;
w5153 <= not w5151 and w5152;
w5154 <= w137 and not w472;
w5155 <= w142 and not w5154;
w5156 <= w146 and not w5155;
w5157 <= w150 and not w5156;
w5158 <= w154 and not w5157;
w5159 <= w158 and not w5158;
w5160 <= w162 and not w5159;
w5161 <= w166 and not w5160;
w5162 <= w170 and not w5161;
w5163 <= w174 and not w5162;
w5164 <= w178 and not w5163;
w5165 <= w182 and not w5164;
w5166 <= w186 and not w5165;
w5167 <= w190 and not w5166;
w5168 <= w194 and not w5167;
w5169 <= w198 and not w5168;
w5170 <= w202 and not w5169;
w5171 <= w206 and not w5170;
w5172 <= w210 and not w5171;
w5173 <= w214 and not w5172;
w5174 <= w218 and not w5173;
w5175 <= w222 and not w5174;
w5176 <= w226 and not w5175;
w5177 <= w230 and not w5176;
w5178 <= w234 and not w5177;
w5179 <= w238 and not w5178;
w5180 <= w242 and not w5179;
w5181 <= w246 and not w5180;
w5182 <= w250 and not w5181;
w5183 <= w254 and not w5182;
w5184 <= w258 and not w5183;
w5185 <= w262 and not w5184;
w5186 <= w266 and not w5185;
w5187 <= w270 and not w5186;
w5188 <= w274 and not w5187;
w5189 <= w278 and not w5188;
w5190 <= w282 and not w5189;
w5191 <= w286 and not w5190;
w5192 <= w290 and not w5191;
w5193 <= w294 and not w5192;
w5194 <= w298 and not w5193;
w5195 <= w302 and not w5194;
w5196 <= w306 and not w5195;
w5197 <= w310 and not w5196;
w5198 <= w314 and not w5197;
w5199 <= w318 and not w5198;
w5200 <= w322 and not w5199;
w5201 <= w326 and not w5200;
w5202 <= w330 and not w5201;
w5203 <= w334 and not w5202;
w5204 <= w1098 and not w5203;
w5205 <= w1100 and not w5204;
w5206 <= w1364 and not w5205;
w5207 <= w345 and not w5206;
w5208 <= w349 and not w5207;
w5209 <= w353 and not w5208;
w5210 <= w357 and not w5209;
w5211 <= w361 and not w5210;
w5212 <= w365 and not w5211;
w5213 <= w369 and not w5212;
w5214 <= w373 and not w5213;
w5215 <= w377 and not w5214;
w5216 <= w381 and not w5215;
w5217 <= w385 and not w5216;
w5218 <= w389 and not w5217;
w5219 <= w393 and not w5218;
w5220 <= w397 and not w5219;
w5221 <= w401 and not w5220;
w5222 <= w405 and not w5221;
w5223 <= w409 and not w5222;
w5224 <= w413 and not w5223;
w5225 <= w417 and not w5224;
w5226 <= w421 and not w5225;
w5227 <= w425 and not w5226;
w5228 <= w429 and not w5227;
w5229 <= w433 and not w5228;
w5230 <= w437 and not w5229;
w5231 <= w441 and not w5230;
w5232 <= w445 and not w5231;
w5233 <= w449 and not w5232;
w5234 <= w453 and not w5233;
w5235 <= w457 and not w5234;
w5236 <= w461 and not w5235;
w5237 <= w465 and not w5236;
w5238 <= req(51) and not w467;
w5239 <= not w5237 and w5238;
w5240 <= w476 and not w809;
w5241 <= w481 and not w5240;
w5242 <= w485 and not w5241;
w5243 <= w489 and not w5242;
w5244 <= w493 and not w5243;
w5245 <= w497 and not w5244;
w5246 <= w501 and not w5245;
w5247 <= w505 and not w5246;
w5248 <= w509 and not w5247;
w5249 <= w513 and not w5248;
w5250 <= w517 and not w5249;
w5251 <= w521 and not w5250;
w5252 <= w525 and not w5251;
w5253 <= w529 and not w5252;
w5254 <= w533 and not w5253;
w5255 <= w537 and not w5254;
w5256 <= w541 and not w5255;
w5257 <= w545 and not w5256;
w5258 <= w549 and not w5257;
w5259 <= w553 and not w5258;
w5260 <= w557 and not w5259;
w5261 <= w561 and not w5260;
w5262 <= w565 and not w5261;
w5263 <= w569 and not w5262;
w5264 <= w573 and not w5263;
w5265 <= w577 and not w5264;
w5266 <= w581 and not w5265;
w5267 <= w585 and not w5266;
w5268 <= w589 and not w5267;
w5269 <= w593 and not w5268;
w5270 <= w597 and not w5269;
w5271 <= w601 and not w5270;
w5272 <= w605 and not w5271;
w5273 <= w609 and not w5272;
w5274 <= w613 and not w5273;
w5275 <= w617 and not w5274;
w5276 <= w621 and not w5275;
w5277 <= w625 and not w5276;
w5278 <= w629 and not w5277;
w5279 <= w633 and not w5278;
w5280 <= w637 and not w5279;
w5281 <= w641 and not w5280;
w5282 <= w645 and not w5281;
w5283 <= w649 and not w5282;
w5284 <= w653 and not w5283;
w5285 <= w657 and not w5284;
w5286 <= w661 and not w5285;
w5287 <= w665 and not w5286;
w5288 <= w669 and not w5287;
w5289 <= w673 and not w5288;
w5290 <= w1188 and not w5289;
w5291 <= w1190 and not w5290;
w5292 <= w1451 and not w5291;
w5293 <= w682 and not w5292;
w5294 <= w686 and not w5293;
w5295 <= w690 and not w5294;
w5296 <= w694 and not w5295;
w5297 <= w698 and not w5296;
w5298 <= w702 and not w5297;
w5299 <= w706 and not w5298;
w5300 <= w710 and not w5299;
w5301 <= w714 and not w5300;
w5302 <= w718 and not w5301;
w5303 <= w722 and not w5302;
w5304 <= w726 and not w5303;
w5305 <= w730 and not w5304;
w5306 <= w734 and not w5305;
w5307 <= w738 and not w5306;
w5308 <= w742 and not w5307;
w5309 <= w746 and not w5308;
w5310 <= w750 and not w5309;
w5311 <= w754 and not w5310;
w5312 <= w758 and not w5311;
w5313 <= w762 and not w5312;
w5314 <= w766 and not w5313;
w5315 <= w770 and not w5314;
w5316 <= w774 and not w5315;
w5317 <= w778 and not w5316;
w5318 <= w782 and not w5317;
w5319 <= w786 and not w5318;
w5320 <= w790 and not w5319;
w5321 <= w794 and not w5320;
w5322 <= w798 and not w5321;
w5323 <= w802 and not w5322;
w5324 <= req(52) and not w804;
w5325 <= not w5323 and w5324;
w5326 <= not w141 and w813;
w5327 <= w818 and not w5326;
w5328 <= w822 and not w5327;
w5329 <= w826 and not w5328;
w5330 <= w830 and not w5329;
w5331 <= w834 and not w5330;
w5332 <= w838 and not w5331;
w5333 <= w842 and not w5332;
w5334 <= w846 and not w5333;
w5335 <= w850 and not w5334;
w5336 <= w854 and not w5335;
w5337 <= w858 and not w5336;
w5338 <= w862 and not w5337;
w5339 <= w866 and not w5338;
w5340 <= w870 and not w5339;
w5341 <= w874 and not w5340;
w5342 <= w878 and not w5341;
w5343 <= w882 and not w5342;
w5344 <= w886 and not w5343;
w5345 <= w890 and not w5344;
w5346 <= w894 and not w5345;
w5347 <= w898 and not w5346;
w5348 <= w902 and not w5347;
w5349 <= w906 and not w5348;
w5350 <= w910 and not w5349;
w5351 <= w914 and not w5350;
w5352 <= w918 and not w5351;
w5353 <= w922 and not w5352;
w5354 <= w926 and not w5353;
w5355 <= w930 and not w5354;
w5356 <= w934 and not w5355;
w5357 <= w938 and not w5356;
w5358 <= w942 and not w5357;
w5359 <= w946 and not w5358;
w5360 <= w950 and not w5359;
w5361 <= w954 and not w5360;
w5362 <= w958 and not w5361;
w5363 <= w962 and not w5362;
w5364 <= w966 and not w5363;
w5365 <= w970 and not w5364;
w5366 <= w974 and not w5365;
w5367 <= w978 and not w5366;
w5368 <= w982 and not w5367;
w5369 <= w986 and not w5368;
w5370 <= w990 and not w5369;
w5371 <= w994 and not w5370;
w5372 <= w998 and not w5371;
w5373 <= w1002 and not w5372;
w5374 <= w1006 and not w5373;
w5375 <= w1010 and not w5374;
w5376 <= w1277 and not w5375;
w5377 <= w6 and not w5376;
w5378 <= w10 and not w5377;
w5379 <= w14 and not w5378;
w5380 <= w18 and not w5379;
w5381 <= w22 and not w5380;
w5382 <= w26 and not w5381;
w5383 <= w30 and not w5382;
w5384 <= w34 and not w5383;
w5385 <= w38 and not w5384;
w5386 <= w42 and not w5385;
w5387 <= w46 and not w5386;
w5388 <= w50 and not w5387;
w5389 <= w54 and not w5388;
w5390 <= w58 and not w5389;
w5391 <= w62 and not w5390;
w5392 <= w66 and not w5391;
w5393 <= w70 and not w5392;
w5394 <= w74 and not w5393;
w5395 <= w78 and not w5394;
w5396 <= w82 and not w5395;
w5397 <= w86 and not w5396;
w5398 <= w90 and not w5397;
w5399 <= w94 and not w5398;
w5400 <= w98 and not w5399;
w5401 <= w102 and not w5400;
w5402 <= w106 and not w5401;
w5403 <= w110 and not w5402;
w5404 <= w114 and not w5403;
w5405 <= w118 and not w5404;
w5406 <= w122 and not w5405;
w5407 <= w126 and not w5406;
w5408 <= w130 and not w5407;
w5409 <= w134 and not w5408;
w5410 <= req(53) and not w136;
w5411 <= not w5409 and w5410;
w5412 <= w145 and not w480;
w5413 <= w150 and not w5412;
w5414 <= w154 and not w5413;
w5415 <= w158 and not w5414;
w5416 <= w162 and not w5415;
w5417 <= w166 and not w5416;
w5418 <= w170 and not w5417;
w5419 <= w174 and not w5418;
w5420 <= w178 and not w5419;
w5421 <= w182 and not w5420;
w5422 <= w186 and not w5421;
w5423 <= w190 and not w5422;
w5424 <= w194 and not w5423;
w5425 <= w198 and not w5424;
w5426 <= w202 and not w5425;
w5427 <= w206 and not w5426;
w5428 <= w210 and not w5427;
w5429 <= w214 and not w5428;
w5430 <= w218 and not w5429;
w5431 <= w222 and not w5430;
w5432 <= w226 and not w5431;
w5433 <= w230 and not w5432;
w5434 <= w234 and not w5433;
w5435 <= w238 and not w5434;
w5436 <= w242 and not w5435;
w5437 <= w246 and not w5436;
w5438 <= w250 and not w5437;
w5439 <= w254 and not w5438;
w5440 <= w258 and not w5439;
w5441 <= w262 and not w5440;
w5442 <= w266 and not w5441;
w5443 <= w270 and not w5442;
w5444 <= w274 and not w5443;
w5445 <= w278 and not w5444;
w5446 <= w282 and not w5445;
w5447 <= w286 and not w5446;
w5448 <= w290 and not w5447;
w5449 <= w294 and not w5448;
w5450 <= w298 and not w5449;
w5451 <= w302 and not w5450;
w5452 <= w306 and not w5451;
w5453 <= w310 and not w5452;
w5454 <= w314 and not w5453;
w5455 <= w318 and not w5454;
w5456 <= w322 and not w5455;
w5457 <= w326 and not w5456;
w5458 <= w330 and not w5457;
w5459 <= w334 and not w5458;
w5460 <= w1098 and not w5459;
w5461 <= w1100 and not w5460;
w5462 <= w1364 and not w5461;
w5463 <= w345 and not w5462;
w5464 <= w349 and not w5463;
w5465 <= w353 and not w5464;
w5466 <= w357 and not w5465;
w5467 <= w361 and not w5466;
w5468 <= w365 and not w5467;
w5469 <= w369 and not w5468;
w5470 <= w373 and not w5469;
w5471 <= w377 and not w5470;
w5472 <= w381 and not w5471;
w5473 <= w385 and not w5472;
w5474 <= w389 and not w5473;
w5475 <= w393 and not w5474;
w5476 <= w397 and not w5475;
w5477 <= w401 and not w5476;
w5478 <= w405 and not w5477;
w5479 <= w409 and not w5478;
w5480 <= w413 and not w5479;
w5481 <= w417 and not w5480;
w5482 <= w421 and not w5481;
w5483 <= w425 and not w5482;
w5484 <= w429 and not w5483;
w5485 <= w433 and not w5484;
w5486 <= w437 and not w5485;
w5487 <= w441 and not w5486;
w5488 <= w445 and not w5487;
w5489 <= w449 and not w5488;
w5490 <= w453 and not w5489;
w5491 <= w457 and not w5490;
w5492 <= w461 and not w5491;
w5493 <= w465 and not w5492;
w5494 <= w469 and not w5493;
w5495 <= w473 and not w5494;
w5496 <= req(54) and not w475;
w5497 <= not w5495 and w5496;
w5498 <= w484 and not w817;
w5499 <= w489 and not w5498;
w5500 <= w493 and not w5499;
w5501 <= w497 and not w5500;
w5502 <= w501 and not w5501;
w5503 <= w505 and not w5502;
w5504 <= w509 and not w5503;
w5505 <= w513 and not w5504;
w5506 <= w517 and not w5505;
w5507 <= w521 and not w5506;
w5508 <= w525 and not w5507;
w5509 <= w529 and not w5508;
w5510 <= w533 and not w5509;
w5511 <= w537 and not w5510;
w5512 <= w541 and not w5511;
w5513 <= w545 and not w5512;
w5514 <= w549 and not w5513;
w5515 <= w553 and not w5514;
w5516 <= w557 and not w5515;
w5517 <= w561 and not w5516;
w5518 <= w565 and not w5517;
w5519 <= w569 and not w5518;
w5520 <= w573 and not w5519;
w5521 <= w577 and not w5520;
w5522 <= w581 and not w5521;
w5523 <= w585 and not w5522;
w5524 <= w589 and not w5523;
w5525 <= w593 and not w5524;
w5526 <= w597 and not w5525;
w5527 <= w601 and not w5526;
w5528 <= w605 and not w5527;
w5529 <= w609 and not w5528;
w5530 <= w613 and not w5529;
w5531 <= w617 and not w5530;
w5532 <= w621 and not w5531;
w5533 <= w625 and not w5532;
w5534 <= w629 and not w5533;
w5535 <= w633 and not w5534;
w5536 <= w637 and not w5535;
w5537 <= w641 and not w5536;
w5538 <= w645 and not w5537;
w5539 <= w649 and not w5538;
w5540 <= w653 and not w5539;
w5541 <= w657 and not w5540;
w5542 <= w661 and not w5541;
w5543 <= w665 and not w5542;
w5544 <= w669 and not w5543;
w5545 <= w673 and not w5544;
w5546 <= w1188 and not w5545;
w5547 <= w1190 and not w5546;
w5548 <= w1451 and not w5547;
w5549 <= w682 and not w5548;
w5550 <= w686 and not w5549;
w5551 <= w690 and not w5550;
w5552 <= w694 and not w5551;
w5553 <= w698 and not w5552;
w5554 <= w702 and not w5553;
w5555 <= w706 and not w5554;
w5556 <= w710 and not w5555;
w5557 <= w714 and not w5556;
w5558 <= w718 and not w5557;
w5559 <= w722 and not w5558;
w5560 <= w726 and not w5559;
w5561 <= w730 and not w5560;
w5562 <= w734 and not w5561;
w5563 <= w738 and not w5562;
w5564 <= w742 and not w5563;
w5565 <= w746 and not w5564;
w5566 <= w750 and not w5565;
w5567 <= w754 and not w5566;
w5568 <= w758 and not w5567;
w5569 <= w762 and not w5568;
w5570 <= w766 and not w5569;
w5571 <= w770 and not w5570;
w5572 <= w774 and not w5571;
w5573 <= w778 and not w5572;
w5574 <= w782 and not w5573;
w5575 <= w786 and not w5574;
w5576 <= w790 and not w5575;
w5577 <= w794 and not w5576;
w5578 <= w798 and not w5577;
w5579 <= w802 and not w5578;
w5580 <= w806 and not w5579;
w5581 <= w810 and not w5580;
w5582 <= req(55) and not w812;
w5583 <= not w5581 and w5582;
w5584 <= not w149 and w821;
w5585 <= w826 and not w5584;
w5586 <= w830 and not w5585;
w5587 <= w834 and not w5586;
w5588 <= w838 and not w5587;
w5589 <= w842 and not w5588;
w5590 <= w846 and not w5589;
w5591 <= w850 and not w5590;
w5592 <= w854 and not w5591;
w5593 <= w858 and not w5592;
w5594 <= w862 and not w5593;
w5595 <= w866 and not w5594;
w5596 <= w870 and not w5595;
w5597 <= w874 and not w5596;
w5598 <= w878 and not w5597;
w5599 <= w882 and not w5598;
w5600 <= w886 and not w5599;
w5601 <= w890 and not w5600;
w5602 <= w894 and not w5601;
w5603 <= w898 and not w5602;
w5604 <= w902 and not w5603;
w5605 <= w906 and not w5604;
w5606 <= w910 and not w5605;
w5607 <= w914 and not w5606;
w5608 <= w918 and not w5607;
w5609 <= w922 and not w5608;
w5610 <= w926 and not w5609;
w5611 <= w930 and not w5610;
w5612 <= w934 and not w5611;
w5613 <= w938 and not w5612;
w5614 <= w942 and not w5613;
w5615 <= w946 and not w5614;
w5616 <= w950 and not w5615;
w5617 <= w954 and not w5616;
w5618 <= w958 and not w5617;
w5619 <= w962 and not w5618;
w5620 <= w966 and not w5619;
w5621 <= w970 and not w5620;
w5622 <= w974 and not w5621;
w5623 <= w978 and not w5622;
w5624 <= w982 and not w5623;
w5625 <= w986 and not w5624;
w5626 <= w990 and not w5625;
w5627 <= w994 and not w5626;
w5628 <= w998 and not w5627;
w5629 <= w1002 and not w5628;
w5630 <= w1006 and not w5629;
w5631 <= w1010 and not w5630;
w5632 <= w1277 and not w5631;
w5633 <= w6 and not w5632;
w5634 <= w10 and not w5633;
w5635 <= w14 and not w5634;
w5636 <= w18 and not w5635;
w5637 <= w22 and not w5636;
w5638 <= w26 and not w5637;
w5639 <= w30 and not w5638;
w5640 <= w34 and not w5639;
w5641 <= w38 and not w5640;
w5642 <= w42 and not w5641;
w5643 <= w46 and not w5642;
w5644 <= w50 and not w5643;
w5645 <= w54 and not w5644;
w5646 <= w58 and not w5645;
w5647 <= w62 and not w5646;
w5648 <= w66 and not w5647;
w5649 <= w70 and not w5648;
w5650 <= w74 and not w5649;
w5651 <= w78 and not w5650;
w5652 <= w82 and not w5651;
w5653 <= w86 and not w5652;
w5654 <= w90 and not w5653;
w5655 <= w94 and not w5654;
w5656 <= w98 and not w5655;
w5657 <= w102 and not w5656;
w5658 <= w106 and not w5657;
w5659 <= w110 and not w5658;
w5660 <= w114 and not w5659;
w5661 <= w118 and not w5660;
w5662 <= w122 and not w5661;
w5663 <= w126 and not w5662;
w5664 <= w130 and not w5663;
w5665 <= w134 and not w5664;
w5666 <= w138 and not w5665;
w5667 <= w142 and not w5666;
w5668 <= req(56) and not w144;
w5669 <= not w5667 and w5668;
w5670 <= w153 and not w488;
w5671 <= w158 and not w5670;
w5672 <= w162 and not w5671;
w5673 <= w166 and not w5672;
w5674 <= w170 and not w5673;
w5675 <= w174 and not w5674;
w5676 <= w178 and not w5675;
w5677 <= w182 and not w5676;
w5678 <= w186 and not w5677;
w5679 <= w190 and not w5678;
w5680 <= w194 and not w5679;
w5681 <= w198 and not w5680;
w5682 <= w202 and not w5681;
w5683 <= w206 and not w5682;
w5684 <= w210 and not w5683;
w5685 <= w214 and not w5684;
w5686 <= w218 and not w5685;
w5687 <= w222 and not w5686;
w5688 <= w226 and not w5687;
w5689 <= w230 and not w5688;
w5690 <= w234 and not w5689;
w5691 <= w238 and not w5690;
w5692 <= w242 and not w5691;
w5693 <= w246 and not w5692;
w5694 <= w250 and not w5693;
w5695 <= w254 and not w5694;
w5696 <= w258 and not w5695;
w5697 <= w262 and not w5696;
w5698 <= w266 and not w5697;
w5699 <= w270 and not w5698;
w5700 <= w274 and not w5699;
w5701 <= w278 and not w5700;
w5702 <= w282 and not w5701;
w5703 <= w286 and not w5702;
w5704 <= w290 and not w5703;
w5705 <= w294 and not w5704;
w5706 <= w298 and not w5705;
w5707 <= w302 and not w5706;
w5708 <= w306 and not w5707;
w5709 <= w310 and not w5708;
w5710 <= w314 and not w5709;
w5711 <= w318 and not w5710;
w5712 <= w322 and not w5711;
w5713 <= w326 and not w5712;
w5714 <= w330 and not w5713;
w5715 <= w334 and not w5714;
w5716 <= w1098 and not w5715;
w5717 <= w1100 and not w5716;
w5718 <= w1364 and not w5717;
w5719 <= w345 and not w5718;
w5720 <= w349 and not w5719;
w5721 <= w353 and not w5720;
w5722 <= w357 and not w5721;
w5723 <= w361 and not w5722;
w5724 <= w365 and not w5723;
w5725 <= w369 and not w5724;
w5726 <= w373 and not w5725;
w5727 <= w377 and not w5726;
w5728 <= w381 and not w5727;
w5729 <= w385 and not w5728;
w5730 <= w389 and not w5729;
w5731 <= w393 and not w5730;
w5732 <= w397 and not w5731;
w5733 <= w401 and not w5732;
w5734 <= w405 and not w5733;
w5735 <= w409 and not w5734;
w5736 <= w413 and not w5735;
w5737 <= w417 and not w5736;
w5738 <= w421 and not w5737;
w5739 <= w425 and not w5738;
w5740 <= w429 and not w5739;
w5741 <= w433 and not w5740;
w5742 <= w437 and not w5741;
w5743 <= w441 and not w5742;
w5744 <= w445 and not w5743;
w5745 <= w449 and not w5744;
w5746 <= w453 and not w5745;
w5747 <= w457 and not w5746;
w5748 <= w461 and not w5747;
w5749 <= w465 and not w5748;
w5750 <= w469 and not w5749;
w5751 <= w473 and not w5750;
w5752 <= w477 and not w5751;
w5753 <= w481 and not w5752;
w5754 <= req(57) and not w483;
w5755 <= not w5753 and w5754;
w5756 <= w492 and not w825;
w5757 <= w497 and not w5756;
w5758 <= w501 and not w5757;
w5759 <= w505 and not w5758;
w5760 <= w509 and not w5759;
w5761 <= w513 and not w5760;
w5762 <= w517 and not w5761;
w5763 <= w521 and not w5762;
w5764 <= w525 and not w5763;
w5765 <= w529 and not w5764;
w5766 <= w533 and not w5765;
w5767 <= w537 and not w5766;
w5768 <= w541 and not w5767;
w5769 <= w545 and not w5768;
w5770 <= w549 and not w5769;
w5771 <= w553 and not w5770;
w5772 <= w557 and not w5771;
w5773 <= w561 and not w5772;
w5774 <= w565 and not w5773;
w5775 <= w569 and not w5774;
w5776 <= w573 and not w5775;
w5777 <= w577 and not w5776;
w5778 <= w581 and not w5777;
w5779 <= w585 and not w5778;
w5780 <= w589 and not w5779;
w5781 <= w593 and not w5780;
w5782 <= w597 and not w5781;
w5783 <= w601 and not w5782;
w5784 <= w605 and not w5783;
w5785 <= w609 and not w5784;
w5786 <= w613 and not w5785;
w5787 <= w617 and not w5786;
w5788 <= w621 and not w5787;
w5789 <= w625 and not w5788;
w5790 <= w629 and not w5789;
w5791 <= w633 and not w5790;
w5792 <= w637 and not w5791;
w5793 <= w641 and not w5792;
w5794 <= w645 and not w5793;
w5795 <= w649 and not w5794;
w5796 <= w653 and not w5795;
w5797 <= w657 and not w5796;
w5798 <= w661 and not w5797;
w5799 <= w665 and not w5798;
w5800 <= w669 and not w5799;
w5801 <= w673 and not w5800;
w5802 <= w1188 and not w5801;
w5803 <= w1190 and not w5802;
w5804 <= w1451 and not w5803;
w5805 <= w682 and not w5804;
w5806 <= w686 and not w5805;
w5807 <= w690 and not w5806;
w5808 <= w694 and not w5807;
w5809 <= w698 and not w5808;
w5810 <= w702 and not w5809;
w5811 <= w706 and not w5810;
w5812 <= w710 and not w5811;
w5813 <= w714 and not w5812;
w5814 <= w718 and not w5813;
w5815 <= w722 and not w5814;
w5816 <= w726 and not w5815;
w5817 <= w730 and not w5816;
w5818 <= w734 and not w5817;
w5819 <= w738 and not w5818;
w5820 <= w742 and not w5819;
w5821 <= w746 and not w5820;
w5822 <= w750 and not w5821;
w5823 <= w754 and not w5822;
w5824 <= w758 and not w5823;
w5825 <= w762 and not w5824;
w5826 <= w766 and not w5825;
w5827 <= w770 and not w5826;
w5828 <= w774 and not w5827;
w5829 <= w778 and not w5828;
w5830 <= w782 and not w5829;
w5831 <= w786 and not w5830;
w5832 <= w790 and not w5831;
w5833 <= w794 and not w5832;
w5834 <= w798 and not w5833;
w5835 <= w802 and not w5834;
w5836 <= w806 and not w5835;
w5837 <= w810 and not w5836;
w5838 <= w814 and not w5837;
w5839 <= w818 and not w5838;
w5840 <= req(58) and not w820;
w5841 <= not w5839 and w5840;
w5842 <= not w157 and w829;
w5843 <= w834 and not w5842;
w5844 <= w838 and not w5843;
w5845 <= w842 and not w5844;
w5846 <= w846 and not w5845;
w5847 <= w850 and not w5846;
w5848 <= w854 and not w5847;
w5849 <= w858 and not w5848;
w5850 <= w862 and not w5849;
w5851 <= w866 and not w5850;
w5852 <= w870 and not w5851;
w5853 <= w874 and not w5852;
w5854 <= w878 and not w5853;
w5855 <= w882 and not w5854;
w5856 <= w886 and not w5855;
w5857 <= w890 and not w5856;
w5858 <= w894 and not w5857;
w5859 <= w898 and not w5858;
w5860 <= w902 and not w5859;
w5861 <= w906 and not w5860;
w5862 <= w910 and not w5861;
w5863 <= w914 and not w5862;
w5864 <= w918 and not w5863;
w5865 <= w922 and not w5864;
w5866 <= w926 and not w5865;
w5867 <= w930 and not w5866;
w5868 <= w934 and not w5867;
w5869 <= w938 and not w5868;
w5870 <= w942 and not w5869;
w5871 <= w946 and not w5870;
w5872 <= w950 and not w5871;
w5873 <= w954 and not w5872;
w5874 <= w958 and not w5873;
w5875 <= w962 and not w5874;
w5876 <= w966 and not w5875;
w5877 <= w970 and not w5876;
w5878 <= w974 and not w5877;
w5879 <= w978 and not w5878;
w5880 <= w982 and not w5879;
w5881 <= w986 and not w5880;
w5882 <= w990 and not w5881;
w5883 <= w994 and not w5882;
w5884 <= w998 and not w5883;
w5885 <= w1002 and not w5884;
w5886 <= w1006 and not w5885;
w5887 <= w1010 and not w5886;
w5888 <= w1277 and not w5887;
w5889 <= w6 and not w5888;
w5890 <= w10 and not w5889;
w5891 <= w14 and not w5890;
w5892 <= w18 and not w5891;
w5893 <= w22 and not w5892;
w5894 <= w26 and not w5893;
w5895 <= w30 and not w5894;
w5896 <= w34 and not w5895;
w5897 <= w38 and not w5896;
w5898 <= w42 and not w5897;
w5899 <= w46 and not w5898;
w5900 <= w50 and not w5899;
w5901 <= w54 and not w5900;
w5902 <= w58 and not w5901;
w5903 <= w62 and not w5902;
w5904 <= w66 and not w5903;
w5905 <= w70 and not w5904;
w5906 <= w74 and not w5905;
w5907 <= w78 and not w5906;
w5908 <= w82 and not w5907;
w5909 <= w86 and not w5908;
w5910 <= w90 and not w5909;
w5911 <= w94 and not w5910;
w5912 <= w98 and not w5911;
w5913 <= w102 and not w5912;
w5914 <= w106 and not w5913;
w5915 <= w110 and not w5914;
w5916 <= w114 and not w5915;
w5917 <= w118 and not w5916;
w5918 <= w122 and not w5917;
w5919 <= w126 and not w5918;
w5920 <= w130 and not w5919;
w5921 <= w134 and not w5920;
w5922 <= w138 and not w5921;
w5923 <= w142 and not w5922;
w5924 <= w146 and not w5923;
w5925 <= w150 and not w5924;
w5926 <= req(59) and not w152;
w5927 <= not w5925 and w5926;
w5928 <= w161 and not w496;
w5929 <= w166 and not w5928;
w5930 <= w170 and not w5929;
w5931 <= w174 and not w5930;
w5932 <= w178 and not w5931;
w5933 <= w182 and not w5932;
w5934 <= w186 and not w5933;
w5935 <= w190 and not w5934;
w5936 <= w194 and not w5935;
w5937 <= w198 and not w5936;
w5938 <= w202 and not w5937;
w5939 <= w206 and not w5938;
w5940 <= w210 and not w5939;
w5941 <= w214 and not w5940;
w5942 <= w218 and not w5941;
w5943 <= w222 and not w5942;
w5944 <= w226 and not w5943;
w5945 <= w230 and not w5944;
w5946 <= w234 and not w5945;
w5947 <= w238 and not w5946;
w5948 <= w242 and not w5947;
w5949 <= w246 and not w5948;
w5950 <= w250 and not w5949;
w5951 <= w254 and not w5950;
w5952 <= w258 and not w5951;
w5953 <= w262 and not w5952;
w5954 <= w266 and not w5953;
w5955 <= w270 and not w5954;
w5956 <= w274 and not w5955;
w5957 <= w278 and not w5956;
w5958 <= w282 and not w5957;
w5959 <= w286 and not w5958;
w5960 <= w290 and not w5959;
w5961 <= w294 and not w5960;
w5962 <= w298 and not w5961;
w5963 <= w302 and not w5962;
w5964 <= w306 and not w5963;
w5965 <= w310 and not w5964;
w5966 <= w314 and not w5965;
w5967 <= w318 and not w5966;
w5968 <= w322 and not w5967;
w5969 <= w326 and not w5968;
w5970 <= w330 and not w5969;
w5971 <= w334 and not w5970;
w5972 <= w1098 and not w5971;
w5973 <= w1100 and not w5972;
w5974 <= w1364 and not w5973;
w5975 <= w345 and not w5974;
w5976 <= w349 and not w5975;
w5977 <= w353 and not w5976;
w5978 <= w357 and not w5977;
w5979 <= w361 and not w5978;
w5980 <= w365 and not w5979;
w5981 <= w369 and not w5980;
w5982 <= w373 and not w5981;
w5983 <= w377 and not w5982;
w5984 <= w381 and not w5983;
w5985 <= w385 and not w5984;
w5986 <= w389 and not w5985;
w5987 <= w393 and not w5986;
w5988 <= w397 and not w5987;
w5989 <= w401 and not w5988;
w5990 <= w405 and not w5989;
w5991 <= w409 and not w5990;
w5992 <= w413 and not w5991;
w5993 <= w417 and not w5992;
w5994 <= w421 and not w5993;
w5995 <= w425 and not w5994;
w5996 <= w429 and not w5995;
w5997 <= w433 and not w5996;
w5998 <= w437 and not w5997;
w5999 <= w441 and not w5998;
w6000 <= w445 and not w5999;
w6001 <= w449 and not w6000;
w6002 <= w453 and not w6001;
w6003 <= w457 and not w6002;
w6004 <= w461 and not w6003;
w6005 <= w465 and not w6004;
w6006 <= w469 and not w6005;
w6007 <= w473 and not w6006;
w6008 <= w477 and not w6007;
w6009 <= w481 and not w6008;
w6010 <= w485 and not w6009;
w6011 <= w489 and not w6010;
w6012 <= req(60) and not w491;
w6013 <= not w6011 and w6012;
w6014 <= w500 and not w833;
w6015 <= w505 and not w6014;
w6016 <= w509 and not w6015;
w6017 <= w513 and not w6016;
w6018 <= w517 and not w6017;
w6019 <= w521 and not w6018;
w6020 <= w525 and not w6019;
w6021 <= w529 and not w6020;
w6022 <= w533 and not w6021;
w6023 <= w537 and not w6022;
w6024 <= w541 and not w6023;
w6025 <= w545 and not w6024;
w6026 <= w549 and not w6025;
w6027 <= w553 and not w6026;
w6028 <= w557 and not w6027;
w6029 <= w561 and not w6028;
w6030 <= w565 and not w6029;
w6031 <= w569 and not w6030;
w6032 <= w573 and not w6031;
w6033 <= w577 and not w6032;
w6034 <= w581 and not w6033;
w6035 <= w585 and not w6034;
w6036 <= w589 and not w6035;
w6037 <= w593 and not w6036;
w6038 <= w597 and not w6037;
w6039 <= w601 and not w6038;
w6040 <= w605 and not w6039;
w6041 <= w609 and not w6040;
w6042 <= w613 and not w6041;
w6043 <= w617 and not w6042;
w6044 <= w621 and not w6043;
w6045 <= w625 and not w6044;
w6046 <= w629 and not w6045;
w6047 <= w633 and not w6046;
w6048 <= w637 and not w6047;
w6049 <= w641 and not w6048;
w6050 <= w645 and not w6049;
w6051 <= w649 and not w6050;
w6052 <= w653 and not w6051;
w6053 <= w657 and not w6052;
w6054 <= w661 and not w6053;
w6055 <= w665 and not w6054;
w6056 <= w669 and not w6055;
w6057 <= w673 and not w6056;
w6058 <= w1188 and not w6057;
w6059 <= w1190 and not w6058;
w6060 <= w1451 and not w6059;
w6061 <= w682 and not w6060;
w6062 <= w686 and not w6061;
w6063 <= w690 and not w6062;
w6064 <= w694 and not w6063;
w6065 <= w698 and not w6064;
w6066 <= w702 and not w6065;
w6067 <= w706 and not w6066;
w6068 <= w710 and not w6067;
w6069 <= w714 and not w6068;
w6070 <= w718 and not w6069;
w6071 <= w722 and not w6070;
w6072 <= w726 and not w6071;
w6073 <= w730 and not w6072;
w6074 <= w734 and not w6073;
w6075 <= w738 and not w6074;
w6076 <= w742 and not w6075;
w6077 <= w746 and not w6076;
w6078 <= w750 and not w6077;
w6079 <= w754 and not w6078;
w6080 <= w758 and not w6079;
w6081 <= w762 and not w6080;
w6082 <= w766 and not w6081;
w6083 <= w770 and not w6082;
w6084 <= w774 and not w6083;
w6085 <= w778 and not w6084;
w6086 <= w782 and not w6085;
w6087 <= w786 and not w6086;
w6088 <= w790 and not w6087;
w6089 <= w794 and not w6088;
w6090 <= w798 and not w6089;
w6091 <= w802 and not w6090;
w6092 <= w806 and not w6091;
w6093 <= w810 and not w6092;
w6094 <= w814 and not w6093;
w6095 <= w818 and not w6094;
w6096 <= w822 and not w6095;
w6097 <= w826 and not w6096;
w6098 <= req(61) and not w828;
w6099 <= not w6097 and w6098;
w6100 <= not w165 and w837;
w6101 <= w842 and not w6100;
w6102 <= w846 and not w6101;
w6103 <= w850 and not w6102;
w6104 <= w854 and not w6103;
w6105 <= w858 and not w6104;
w6106 <= w862 and not w6105;
w6107 <= w866 and not w6106;
w6108 <= w870 and not w6107;
w6109 <= w874 and not w6108;
w6110 <= w878 and not w6109;
w6111 <= w882 and not w6110;
w6112 <= w886 and not w6111;
w6113 <= w890 and not w6112;
w6114 <= w894 and not w6113;
w6115 <= w898 and not w6114;
w6116 <= w902 and not w6115;
w6117 <= w906 and not w6116;
w6118 <= w910 and not w6117;
w6119 <= w914 and not w6118;
w6120 <= w918 and not w6119;
w6121 <= w922 and not w6120;
w6122 <= w926 and not w6121;
w6123 <= w930 and not w6122;
w6124 <= w934 and not w6123;
w6125 <= w938 and not w6124;
w6126 <= w942 and not w6125;
w6127 <= w946 and not w6126;
w6128 <= w950 and not w6127;
w6129 <= w954 and not w6128;
w6130 <= w958 and not w6129;
w6131 <= w962 and not w6130;
w6132 <= w966 and not w6131;
w6133 <= w970 and not w6132;
w6134 <= w974 and not w6133;
w6135 <= w978 and not w6134;
w6136 <= w982 and not w6135;
w6137 <= w986 and not w6136;
w6138 <= w990 and not w6137;
w6139 <= w994 and not w6138;
w6140 <= w998 and not w6139;
w6141 <= w1002 and not w6140;
w6142 <= w1006 and not w6141;
w6143 <= w1010 and not w6142;
w6144 <= w1277 and not w6143;
w6145 <= w6 and not w6144;
w6146 <= w10 and not w6145;
w6147 <= w14 and not w6146;
w6148 <= w18 and not w6147;
w6149 <= w22 and not w6148;
w6150 <= w26 and not w6149;
w6151 <= w30 and not w6150;
w6152 <= w34 and not w6151;
w6153 <= w38 and not w6152;
w6154 <= w42 and not w6153;
w6155 <= w46 and not w6154;
w6156 <= w50 and not w6155;
w6157 <= w54 and not w6156;
w6158 <= w58 and not w6157;
w6159 <= w62 and not w6158;
w6160 <= w66 and not w6159;
w6161 <= w70 and not w6160;
w6162 <= w74 and not w6161;
w6163 <= w78 and not w6162;
w6164 <= w82 and not w6163;
w6165 <= w86 and not w6164;
w6166 <= w90 and not w6165;
w6167 <= w94 and not w6166;
w6168 <= w98 and not w6167;
w6169 <= w102 and not w6168;
w6170 <= w106 and not w6169;
w6171 <= w110 and not w6170;
w6172 <= w114 and not w6171;
w6173 <= w118 and not w6172;
w6174 <= w122 and not w6173;
w6175 <= w126 and not w6174;
w6176 <= w130 and not w6175;
w6177 <= w134 and not w6176;
w6178 <= w138 and not w6177;
w6179 <= w142 and not w6178;
w6180 <= w146 and not w6179;
w6181 <= w150 and not w6180;
w6182 <= w154 and not w6181;
w6183 <= w158 and not w6182;
w6184 <= req(62) and not w160;
w6185 <= not w6183 and w6184;
w6186 <= w169 and not w504;
w6187 <= w174 and not w6186;
w6188 <= w178 and not w6187;
w6189 <= w182 and not w6188;
w6190 <= w186 and not w6189;
w6191 <= w190 and not w6190;
w6192 <= w194 and not w6191;
w6193 <= w198 and not w6192;
w6194 <= w202 and not w6193;
w6195 <= w206 and not w6194;
w6196 <= w210 and not w6195;
w6197 <= w214 and not w6196;
w6198 <= w218 and not w6197;
w6199 <= w222 and not w6198;
w6200 <= w226 and not w6199;
w6201 <= w230 and not w6200;
w6202 <= w234 and not w6201;
w6203 <= w238 and not w6202;
w6204 <= w242 and not w6203;
w6205 <= w246 and not w6204;
w6206 <= w250 and not w6205;
w6207 <= w254 and not w6206;
w6208 <= w258 and not w6207;
w6209 <= w262 and not w6208;
w6210 <= w266 and not w6209;
w6211 <= w270 and not w6210;
w6212 <= w274 and not w6211;
w6213 <= w278 and not w6212;
w6214 <= w282 and not w6213;
w6215 <= w286 and not w6214;
w6216 <= w290 and not w6215;
w6217 <= w294 and not w6216;
w6218 <= w298 and not w6217;
w6219 <= w302 and not w6218;
w6220 <= w306 and not w6219;
w6221 <= w310 and not w6220;
w6222 <= w314 and not w6221;
w6223 <= w318 and not w6222;
w6224 <= w322 and not w6223;
w6225 <= w326 and not w6224;
w6226 <= w330 and not w6225;
w6227 <= w334 and not w6226;
w6228 <= w1098 and not w6227;
w6229 <= w1100 and not w6228;
w6230 <= w1364 and not w6229;
w6231 <= w345 and not w6230;
w6232 <= w349 and not w6231;
w6233 <= w353 and not w6232;
w6234 <= w357 and not w6233;
w6235 <= w361 and not w6234;
w6236 <= w365 and not w6235;
w6237 <= w369 and not w6236;
w6238 <= w373 and not w6237;
w6239 <= w377 and not w6238;
w6240 <= w381 and not w6239;
w6241 <= w385 and not w6240;
w6242 <= w389 and not w6241;
w6243 <= w393 and not w6242;
w6244 <= w397 and not w6243;
w6245 <= w401 and not w6244;
w6246 <= w405 and not w6245;
w6247 <= w409 and not w6246;
w6248 <= w413 and not w6247;
w6249 <= w417 and not w6248;
w6250 <= w421 and not w6249;
w6251 <= w425 and not w6250;
w6252 <= w429 and not w6251;
w6253 <= w433 and not w6252;
w6254 <= w437 and not w6253;
w6255 <= w441 and not w6254;
w6256 <= w445 and not w6255;
w6257 <= w449 and not w6256;
w6258 <= w453 and not w6257;
w6259 <= w457 and not w6258;
w6260 <= w461 and not w6259;
w6261 <= w465 and not w6260;
w6262 <= w469 and not w6261;
w6263 <= w473 and not w6262;
w6264 <= w477 and not w6263;
w6265 <= w481 and not w6264;
w6266 <= w485 and not w6265;
w6267 <= w489 and not w6266;
w6268 <= w493 and not w6267;
w6269 <= w497 and not w6268;
w6270 <= req(63) and not w499;
w6271 <= not w6269 and w6270;
w6272 <= w508 and not w841;
w6273 <= w513 and not w6272;
w6274 <= w517 and not w6273;
w6275 <= w521 and not w6274;
w6276 <= w525 and not w6275;
w6277 <= w529 and not w6276;
w6278 <= w533 and not w6277;
w6279 <= w537 and not w6278;
w6280 <= w541 and not w6279;
w6281 <= w545 and not w6280;
w6282 <= w549 and not w6281;
w6283 <= w553 and not w6282;
w6284 <= w557 and not w6283;
w6285 <= w561 and not w6284;
w6286 <= w565 and not w6285;
w6287 <= w569 and not w6286;
w6288 <= w573 and not w6287;
w6289 <= w577 and not w6288;
w6290 <= w581 and not w6289;
w6291 <= w585 and not w6290;
w6292 <= w589 and not w6291;
w6293 <= w593 and not w6292;
w6294 <= w597 and not w6293;
w6295 <= w601 and not w6294;
w6296 <= w605 and not w6295;
w6297 <= w609 and not w6296;
w6298 <= w613 and not w6297;
w6299 <= w617 and not w6298;
w6300 <= w621 and not w6299;
w6301 <= w625 and not w6300;
w6302 <= w629 and not w6301;
w6303 <= w633 and not w6302;
w6304 <= w637 and not w6303;
w6305 <= w641 and not w6304;
w6306 <= w645 and not w6305;
w6307 <= w649 and not w6306;
w6308 <= w653 and not w6307;
w6309 <= w657 and not w6308;
w6310 <= w661 and not w6309;
w6311 <= w665 and not w6310;
w6312 <= w669 and not w6311;
w6313 <= w673 and not w6312;
w6314 <= w1188 and not w6313;
w6315 <= w1190 and not w6314;
w6316 <= w1451 and not w6315;
w6317 <= w682 and not w6316;
w6318 <= w686 and not w6317;
w6319 <= w690 and not w6318;
w6320 <= w694 and not w6319;
w6321 <= w698 and not w6320;
w6322 <= w702 and not w6321;
w6323 <= w706 and not w6322;
w6324 <= w710 and not w6323;
w6325 <= w714 and not w6324;
w6326 <= w718 and not w6325;
w6327 <= w722 and not w6326;
w6328 <= w726 and not w6327;
w6329 <= w730 and not w6328;
w6330 <= w734 and not w6329;
w6331 <= w738 and not w6330;
w6332 <= w742 and not w6331;
w6333 <= w746 and not w6332;
w6334 <= w750 and not w6333;
w6335 <= w754 and not w6334;
w6336 <= w758 and not w6335;
w6337 <= w762 and not w6336;
w6338 <= w766 and not w6337;
w6339 <= w770 and not w6338;
w6340 <= w774 and not w6339;
w6341 <= w778 and not w6340;
w6342 <= w782 and not w6341;
w6343 <= w786 and not w6342;
w6344 <= w790 and not w6343;
w6345 <= w794 and not w6344;
w6346 <= w798 and not w6345;
w6347 <= w802 and not w6346;
w6348 <= w806 and not w6347;
w6349 <= w810 and not w6348;
w6350 <= w814 and not w6349;
w6351 <= w818 and not w6350;
w6352 <= w822 and not w6351;
w6353 <= w826 and not w6352;
w6354 <= w830 and not w6353;
w6355 <= w834 and not w6354;
w6356 <= req(64) and not w836;
w6357 <= not w6355 and w6356;
w6358 <= not w173 and w845;
w6359 <= w850 and not w6358;
w6360 <= w854 and not w6359;
w6361 <= w858 and not w6360;
w6362 <= w862 and not w6361;
w6363 <= w866 and not w6362;
w6364 <= w870 and not w6363;
w6365 <= w874 and not w6364;
w6366 <= w878 and not w6365;
w6367 <= w882 and not w6366;
w6368 <= w886 and not w6367;
w6369 <= w890 and not w6368;
w6370 <= w894 and not w6369;
w6371 <= w898 and not w6370;
w6372 <= w902 and not w6371;
w6373 <= w906 and not w6372;
w6374 <= w910 and not w6373;
w6375 <= w914 and not w6374;
w6376 <= w918 and not w6375;
w6377 <= w922 and not w6376;
w6378 <= w926 and not w6377;
w6379 <= w930 and not w6378;
w6380 <= w934 and not w6379;
w6381 <= w938 and not w6380;
w6382 <= w942 and not w6381;
w6383 <= w946 and not w6382;
w6384 <= w950 and not w6383;
w6385 <= w954 and not w6384;
w6386 <= w958 and not w6385;
w6387 <= w962 and not w6386;
w6388 <= w966 and not w6387;
w6389 <= w970 and not w6388;
w6390 <= w974 and not w6389;
w6391 <= w978 and not w6390;
w6392 <= w982 and not w6391;
w6393 <= w986 and not w6392;
w6394 <= w990 and not w6393;
w6395 <= w994 and not w6394;
w6396 <= w998 and not w6395;
w6397 <= w1002 and not w6396;
w6398 <= w1006 and not w6397;
w6399 <= w1010 and not w6398;
w6400 <= w1277 and not w6399;
w6401 <= w6 and not w6400;
w6402 <= w10 and not w6401;
w6403 <= w14 and not w6402;
w6404 <= w18 and not w6403;
w6405 <= w22 and not w6404;
w6406 <= w26 and not w6405;
w6407 <= w30 and not w6406;
w6408 <= w34 and not w6407;
w6409 <= w38 and not w6408;
w6410 <= w42 and not w6409;
w6411 <= w46 and not w6410;
w6412 <= w50 and not w6411;
w6413 <= w54 and not w6412;
w6414 <= w58 and not w6413;
w6415 <= w62 and not w6414;
w6416 <= w66 and not w6415;
w6417 <= w70 and not w6416;
w6418 <= w74 and not w6417;
w6419 <= w78 and not w6418;
w6420 <= w82 and not w6419;
w6421 <= w86 and not w6420;
w6422 <= w90 and not w6421;
w6423 <= w94 and not w6422;
w6424 <= w98 and not w6423;
w6425 <= w102 and not w6424;
w6426 <= w106 and not w6425;
w6427 <= w110 and not w6426;
w6428 <= w114 and not w6427;
w6429 <= w118 and not w6428;
w6430 <= w122 and not w6429;
w6431 <= w126 and not w6430;
w6432 <= w130 and not w6431;
w6433 <= w134 and not w6432;
w6434 <= w138 and not w6433;
w6435 <= w142 and not w6434;
w6436 <= w146 and not w6435;
w6437 <= w150 and not w6436;
w6438 <= w154 and not w6437;
w6439 <= w158 and not w6438;
w6440 <= w162 and not w6439;
w6441 <= w166 and not w6440;
w6442 <= req(65) and not w168;
w6443 <= not w6441 and w6442;
w6444 <= w177 and not w512;
w6445 <= w182 and not w6444;
w6446 <= w186 and not w6445;
w6447 <= w190 and not w6446;
w6448 <= w194 and not w6447;
w6449 <= w198 and not w6448;
w6450 <= w202 and not w6449;
w6451 <= w206 and not w6450;
w6452 <= w210 and not w6451;
w6453 <= w214 and not w6452;
w6454 <= w218 and not w6453;
w6455 <= w222 and not w6454;
w6456 <= w226 and not w6455;
w6457 <= w230 and not w6456;
w6458 <= w234 and not w6457;
w6459 <= w238 and not w6458;
w6460 <= w242 and not w6459;
w6461 <= w246 and not w6460;
w6462 <= w250 and not w6461;
w6463 <= w254 and not w6462;
w6464 <= w258 and not w6463;
w6465 <= w262 and not w6464;
w6466 <= w266 and not w6465;
w6467 <= w270 and not w6466;
w6468 <= w274 and not w6467;
w6469 <= w278 and not w6468;
w6470 <= w282 and not w6469;
w6471 <= w286 and not w6470;
w6472 <= w290 and not w6471;
w6473 <= w294 and not w6472;
w6474 <= w298 and not w6473;
w6475 <= w302 and not w6474;
w6476 <= w306 and not w6475;
w6477 <= w310 and not w6476;
w6478 <= w314 and not w6477;
w6479 <= w318 and not w6478;
w6480 <= w322 and not w6479;
w6481 <= w326 and not w6480;
w6482 <= w330 and not w6481;
w6483 <= w334 and not w6482;
w6484 <= w1098 and not w6483;
w6485 <= w1100 and not w6484;
w6486 <= w1364 and not w6485;
w6487 <= w345 and not w6486;
w6488 <= w349 and not w6487;
w6489 <= w353 and not w6488;
w6490 <= w357 and not w6489;
w6491 <= w361 and not w6490;
w6492 <= w365 and not w6491;
w6493 <= w369 and not w6492;
w6494 <= w373 and not w6493;
w6495 <= w377 and not w6494;
w6496 <= w381 and not w6495;
w6497 <= w385 and not w6496;
w6498 <= w389 and not w6497;
w6499 <= w393 and not w6498;
w6500 <= w397 and not w6499;
w6501 <= w401 and not w6500;
w6502 <= w405 and not w6501;
w6503 <= w409 and not w6502;
w6504 <= w413 and not w6503;
w6505 <= w417 and not w6504;
w6506 <= w421 and not w6505;
w6507 <= w425 and not w6506;
w6508 <= w429 and not w6507;
w6509 <= w433 and not w6508;
w6510 <= w437 and not w6509;
w6511 <= w441 and not w6510;
w6512 <= w445 and not w6511;
w6513 <= w449 and not w6512;
w6514 <= w453 and not w6513;
w6515 <= w457 and not w6514;
w6516 <= w461 and not w6515;
w6517 <= w465 and not w6516;
w6518 <= w469 and not w6517;
w6519 <= w473 and not w6518;
w6520 <= w477 and not w6519;
w6521 <= w481 and not w6520;
w6522 <= w485 and not w6521;
w6523 <= w489 and not w6522;
w6524 <= w493 and not w6523;
w6525 <= w497 and not w6524;
w6526 <= w501 and not w6525;
w6527 <= w505 and not w6526;
w6528 <= req(66) and not w507;
w6529 <= not w6527 and w6528;
w6530 <= w516 and not w849;
w6531 <= w521 and not w6530;
w6532 <= w525 and not w6531;
w6533 <= w529 and not w6532;
w6534 <= w533 and not w6533;
w6535 <= w537 and not w6534;
w6536 <= w541 and not w6535;
w6537 <= w545 and not w6536;
w6538 <= w549 and not w6537;
w6539 <= w553 and not w6538;
w6540 <= w557 and not w6539;
w6541 <= w561 and not w6540;
w6542 <= w565 and not w6541;
w6543 <= w569 and not w6542;
w6544 <= w573 and not w6543;
w6545 <= w577 and not w6544;
w6546 <= w581 and not w6545;
w6547 <= w585 and not w6546;
w6548 <= w589 and not w6547;
w6549 <= w593 and not w6548;
w6550 <= w597 and not w6549;
w6551 <= w601 and not w6550;
w6552 <= w605 and not w6551;
w6553 <= w609 and not w6552;
w6554 <= w613 and not w6553;
w6555 <= w617 and not w6554;
w6556 <= w621 and not w6555;
w6557 <= w625 and not w6556;
w6558 <= w629 and not w6557;
w6559 <= w633 and not w6558;
w6560 <= w637 and not w6559;
w6561 <= w641 and not w6560;
w6562 <= w645 and not w6561;
w6563 <= w649 and not w6562;
w6564 <= w653 and not w6563;
w6565 <= w657 and not w6564;
w6566 <= w661 and not w6565;
w6567 <= w665 and not w6566;
w6568 <= w669 and not w6567;
w6569 <= w673 and not w6568;
w6570 <= w1188 and not w6569;
w6571 <= w1190 and not w6570;
w6572 <= w1451 and not w6571;
w6573 <= w682 and not w6572;
w6574 <= w686 and not w6573;
w6575 <= w690 and not w6574;
w6576 <= w694 and not w6575;
w6577 <= w698 and not w6576;
w6578 <= w702 and not w6577;
w6579 <= w706 and not w6578;
w6580 <= w710 and not w6579;
w6581 <= w714 and not w6580;
w6582 <= w718 and not w6581;
w6583 <= w722 and not w6582;
w6584 <= w726 and not w6583;
w6585 <= w730 and not w6584;
w6586 <= w734 and not w6585;
w6587 <= w738 and not w6586;
w6588 <= w742 and not w6587;
w6589 <= w746 and not w6588;
w6590 <= w750 and not w6589;
w6591 <= w754 and not w6590;
w6592 <= w758 and not w6591;
w6593 <= w762 and not w6592;
w6594 <= w766 and not w6593;
w6595 <= w770 and not w6594;
w6596 <= w774 and not w6595;
w6597 <= w778 and not w6596;
w6598 <= w782 and not w6597;
w6599 <= w786 and not w6598;
w6600 <= w790 and not w6599;
w6601 <= w794 and not w6600;
w6602 <= w798 and not w6601;
w6603 <= w802 and not w6602;
w6604 <= w806 and not w6603;
w6605 <= w810 and not w6604;
w6606 <= w814 and not w6605;
w6607 <= w818 and not w6606;
w6608 <= w822 and not w6607;
w6609 <= w826 and not w6608;
w6610 <= w830 and not w6609;
w6611 <= w834 and not w6610;
w6612 <= w838 and not w6611;
w6613 <= w842 and not w6612;
w6614 <= req(67) and not w844;
w6615 <= not w6613 and w6614;
w6616 <= not w181 and w853;
w6617 <= w858 and not w6616;
w6618 <= w862 and not w6617;
w6619 <= w866 and not w6618;
w6620 <= w870 and not w6619;
w6621 <= w874 and not w6620;
w6622 <= w878 and not w6621;
w6623 <= w882 and not w6622;
w6624 <= w886 and not w6623;
w6625 <= w890 and not w6624;
w6626 <= w894 and not w6625;
w6627 <= w898 and not w6626;
w6628 <= w902 and not w6627;
w6629 <= w906 and not w6628;
w6630 <= w910 and not w6629;
w6631 <= w914 and not w6630;
w6632 <= w918 and not w6631;
w6633 <= w922 and not w6632;
w6634 <= w926 and not w6633;
w6635 <= w930 and not w6634;
w6636 <= w934 and not w6635;
w6637 <= w938 and not w6636;
w6638 <= w942 and not w6637;
w6639 <= w946 and not w6638;
w6640 <= w950 and not w6639;
w6641 <= w954 and not w6640;
w6642 <= w958 and not w6641;
w6643 <= w962 and not w6642;
w6644 <= w966 and not w6643;
w6645 <= w970 and not w6644;
w6646 <= w974 and not w6645;
w6647 <= w978 and not w6646;
w6648 <= w982 and not w6647;
w6649 <= w986 and not w6648;
w6650 <= w990 and not w6649;
w6651 <= w994 and not w6650;
w6652 <= w998 and not w6651;
w6653 <= w1002 and not w6652;
w6654 <= w1006 and not w6653;
w6655 <= w1010 and not w6654;
w6656 <= w1277 and not w6655;
w6657 <= w6 and not w6656;
w6658 <= w10 and not w6657;
w6659 <= w14 and not w6658;
w6660 <= w18 and not w6659;
w6661 <= w22 and not w6660;
w6662 <= w26 and not w6661;
w6663 <= w30 and not w6662;
w6664 <= w34 and not w6663;
w6665 <= w38 and not w6664;
w6666 <= w42 and not w6665;
w6667 <= w46 and not w6666;
w6668 <= w50 and not w6667;
w6669 <= w54 and not w6668;
w6670 <= w58 and not w6669;
w6671 <= w62 and not w6670;
w6672 <= w66 and not w6671;
w6673 <= w70 and not w6672;
w6674 <= w74 and not w6673;
w6675 <= w78 and not w6674;
w6676 <= w82 and not w6675;
w6677 <= w86 and not w6676;
w6678 <= w90 and not w6677;
w6679 <= w94 and not w6678;
w6680 <= w98 and not w6679;
w6681 <= w102 and not w6680;
w6682 <= w106 and not w6681;
w6683 <= w110 and not w6682;
w6684 <= w114 and not w6683;
w6685 <= w118 and not w6684;
w6686 <= w122 and not w6685;
w6687 <= w126 and not w6686;
w6688 <= w130 and not w6687;
w6689 <= w134 and not w6688;
w6690 <= w138 and not w6689;
w6691 <= w142 and not w6690;
w6692 <= w146 and not w6691;
w6693 <= w150 and not w6692;
w6694 <= w154 and not w6693;
w6695 <= w158 and not w6694;
w6696 <= w162 and not w6695;
w6697 <= w166 and not w6696;
w6698 <= w170 and not w6697;
w6699 <= w174 and not w6698;
w6700 <= req(68) and not w176;
w6701 <= not w6699 and w6700;
w6702 <= w185 and not w520;
w6703 <= w190 and not w6702;
w6704 <= w194 and not w6703;
w6705 <= w198 and not w6704;
w6706 <= w202 and not w6705;
w6707 <= w206 and not w6706;
w6708 <= w210 and not w6707;
w6709 <= w214 and not w6708;
w6710 <= w218 and not w6709;
w6711 <= w222 and not w6710;
w6712 <= w226 and not w6711;
w6713 <= w230 and not w6712;
w6714 <= w234 and not w6713;
w6715 <= w238 and not w6714;
w6716 <= w242 and not w6715;
w6717 <= w246 and not w6716;
w6718 <= w250 and not w6717;
w6719 <= w254 and not w6718;
w6720 <= w258 and not w6719;
w6721 <= w262 and not w6720;
w6722 <= w266 and not w6721;
w6723 <= w270 and not w6722;
w6724 <= w274 and not w6723;
w6725 <= w278 and not w6724;
w6726 <= w282 and not w6725;
w6727 <= w286 and not w6726;
w6728 <= w290 and not w6727;
w6729 <= w294 and not w6728;
w6730 <= w298 and not w6729;
w6731 <= w302 and not w6730;
w6732 <= w306 and not w6731;
w6733 <= w310 and not w6732;
w6734 <= w314 and not w6733;
w6735 <= w318 and not w6734;
w6736 <= w322 and not w6735;
w6737 <= w326 and not w6736;
w6738 <= w330 and not w6737;
w6739 <= w334 and not w6738;
w6740 <= w1098 and not w6739;
w6741 <= w1100 and not w6740;
w6742 <= w1364 and not w6741;
w6743 <= w345 and not w6742;
w6744 <= w349 and not w6743;
w6745 <= w353 and not w6744;
w6746 <= w357 and not w6745;
w6747 <= w361 and not w6746;
w6748 <= w365 and not w6747;
w6749 <= w369 and not w6748;
w6750 <= w373 and not w6749;
w6751 <= w377 and not w6750;
w6752 <= w381 and not w6751;
w6753 <= w385 and not w6752;
w6754 <= w389 and not w6753;
w6755 <= w393 and not w6754;
w6756 <= w397 and not w6755;
w6757 <= w401 and not w6756;
w6758 <= w405 and not w6757;
w6759 <= w409 and not w6758;
w6760 <= w413 and not w6759;
w6761 <= w417 and not w6760;
w6762 <= w421 and not w6761;
w6763 <= w425 and not w6762;
w6764 <= w429 and not w6763;
w6765 <= w433 and not w6764;
w6766 <= w437 and not w6765;
w6767 <= w441 and not w6766;
w6768 <= w445 and not w6767;
w6769 <= w449 and not w6768;
w6770 <= w453 and not w6769;
w6771 <= w457 and not w6770;
w6772 <= w461 and not w6771;
w6773 <= w465 and not w6772;
w6774 <= w469 and not w6773;
w6775 <= w473 and not w6774;
w6776 <= w477 and not w6775;
w6777 <= w481 and not w6776;
w6778 <= w485 and not w6777;
w6779 <= w489 and not w6778;
w6780 <= w493 and not w6779;
w6781 <= w497 and not w6780;
w6782 <= w501 and not w6781;
w6783 <= w505 and not w6782;
w6784 <= w509 and not w6783;
w6785 <= w513 and not w6784;
w6786 <= req(69) and not w515;
w6787 <= not w6785 and w6786;
w6788 <= w524 and not w857;
w6789 <= w529 and not w6788;
w6790 <= w533 and not w6789;
w6791 <= w537 and not w6790;
w6792 <= w541 and not w6791;
w6793 <= w545 and not w6792;
w6794 <= w549 and not w6793;
w6795 <= w553 and not w6794;
w6796 <= w557 and not w6795;
w6797 <= w561 and not w6796;
w6798 <= w565 and not w6797;
w6799 <= w569 and not w6798;
w6800 <= w573 and not w6799;
w6801 <= w577 and not w6800;
w6802 <= w581 and not w6801;
w6803 <= w585 and not w6802;
w6804 <= w589 and not w6803;
w6805 <= w593 and not w6804;
w6806 <= w597 and not w6805;
w6807 <= w601 and not w6806;
w6808 <= w605 and not w6807;
w6809 <= w609 and not w6808;
w6810 <= w613 and not w6809;
w6811 <= w617 and not w6810;
w6812 <= w621 and not w6811;
w6813 <= w625 and not w6812;
w6814 <= w629 and not w6813;
w6815 <= w633 and not w6814;
w6816 <= w637 and not w6815;
w6817 <= w641 and not w6816;
w6818 <= w645 and not w6817;
w6819 <= w649 and not w6818;
w6820 <= w653 and not w6819;
w6821 <= w657 and not w6820;
w6822 <= w661 and not w6821;
w6823 <= w665 and not w6822;
w6824 <= w669 and not w6823;
w6825 <= w673 and not w6824;
w6826 <= w1188 and not w6825;
w6827 <= w1190 and not w6826;
w6828 <= w1451 and not w6827;
w6829 <= w682 and not w6828;
w6830 <= w686 and not w6829;
w6831 <= w690 and not w6830;
w6832 <= w694 and not w6831;
w6833 <= w698 and not w6832;
w6834 <= w702 and not w6833;
w6835 <= w706 and not w6834;
w6836 <= w710 and not w6835;
w6837 <= w714 and not w6836;
w6838 <= w718 and not w6837;
w6839 <= w722 and not w6838;
w6840 <= w726 and not w6839;
w6841 <= w730 and not w6840;
w6842 <= w734 and not w6841;
w6843 <= w738 and not w6842;
w6844 <= w742 and not w6843;
w6845 <= w746 and not w6844;
w6846 <= w750 and not w6845;
w6847 <= w754 and not w6846;
w6848 <= w758 and not w6847;
w6849 <= w762 and not w6848;
w6850 <= w766 and not w6849;
w6851 <= w770 and not w6850;
w6852 <= w774 and not w6851;
w6853 <= w778 and not w6852;
w6854 <= w782 and not w6853;
w6855 <= w786 and not w6854;
w6856 <= w790 and not w6855;
w6857 <= w794 and not w6856;
w6858 <= w798 and not w6857;
w6859 <= w802 and not w6858;
w6860 <= w806 and not w6859;
w6861 <= w810 and not w6860;
w6862 <= w814 and not w6861;
w6863 <= w818 and not w6862;
w6864 <= w822 and not w6863;
w6865 <= w826 and not w6864;
w6866 <= w830 and not w6865;
w6867 <= w834 and not w6866;
w6868 <= w838 and not w6867;
w6869 <= w842 and not w6868;
w6870 <= w846 and not w6869;
w6871 <= w850 and not w6870;
w6872 <= req(70) and not w852;
w6873 <= not w6871 and w6872;
w6874 <= not w189 and w861;
w6875 <= w866 and not w6874;
w6876 <= w870 and not w6875;
w6877 <= w874 and not w6876;
w6878 <= w878 and not w6877;
w6879 <= w882 and not w6878;
w6880 <= w886 and not w6879;
w6881 <= w890 and not w6880;
w6882 <= w894 and not w6881;
w6883 <= w898 and not w6882;
w6884 <= w902 and not w6883;
w6885 <= w906 and not w6884;
w6886 <= w910 and not w6885;
w6887 <= w914 and not w6886;
w6888 <= w918 and not w6887;
w6889 <= w922 and not w6888;
w6890 <= w926 and not w6889;
w6891 <= w930 and not w6890;
w6892 <= w934 and not w6891;
w6893 <= w938 and not w6892;
w6894 <= w942 and not w6893;
w6895 <= w946 and not w6894;
w6896 <= w950 and not w6895;
w6897 <= w954 and not w6896;
w6898 <= w958 and not w6897;
w6899 <= w962 and not w6898;
w6900 <= w966 and not w6899;
w6901 <= w970 and not w6900;
w6902 <= w974 and not w6901;
w6903 <= w978 and not w6902;
w6904 <= w982 and not w6903;
w6905 <= w986 and not w6904;
w6906 <= w990 and not w6905;
w6907 <= w994 and not w6906;
w6908 <= w998 and not w6907;
w6909 <= w1002 and not w6908;
w6910 <= w1006 and not w6909;
w6911 <= w1010 and not w6910;
w6912 <= w1277 and not w6911;
w6913 <= w6 and not w6912;
w6914 <= w10 and not w6913;
w6915 <= w14 and not w6914;
w6916 <= w18 and not w6915;
w6917 <= w22 and not w6916;
w6918 <= w26 and not w6917;
w6919 <= w30 and not w6918;
w6920 <= w34 and not w6919;
w6921 <= w38 and not w6920;
w6922 <= w42 and not w6921;
w6923 <= w46 and not w6922;
w6924 <= w50 and not w6923;
w6925 <= w54 and not w6924;
w6926 <= w58 and not w6925;
w6927 <= w62 and not w6926;
w6928 <= w66 and not w6927;
w6929 <= w70 and not w6928;
w6930 <= w74 and not w6929;
w6931 <= w78 and not w6930;
w6932 <= w82 and not w6931;
w6933 <= w86 and not w6932;
w6934 <= w90 and not w6933;
w6935 <= w94 and not w6934;
w6936 <= w98 and not w6935;
w6937 <= w102 and not w6936;
w6938 <= w106 and not w6937;
w6939 <= w110 and not w6938;
w6940 <= w114 and not w6939;
w6941 <= w118 and not w6940;
w6942 <= w122 and not w6941;
w6943 <= w126 and not w6942;
w6944 <= w130 and not w6943;
w6945 <= w134 and not w6944;
w6946 <= w138 and not w6945;
w6947 <= w142 and not w6946;
w6948 <= w146 and not w6947;
w6949 <= w150 and not w6948;
w6950 <= w154 and not w6949;
w6951 <= w158 and not w6950;
w6952 <= w162 and not w6951;
w6953 <= w166 and not w6952;
w6954 <= w170 and not w6953;
w6955 <= w174 and not w6954;
w6956 <= w178 and not w6955;
w6957 <= w182 and not w6956;
w6958 <= req(71) and not w184;
w6959 <= not w6957 and w6958;
w6960 <= w193 and not w528;
w6961 <= w198 and not w6960;
w6962 <= w202 and not w6961;
w6963 <= w206 and not w6962;
w6964 <= w210 and not w6963;
w6965 <= w214 and not w6964;
w6966 <= w218 and not w6965;
w6967 <= w222 and not w6966;
w6968 <= w226 and not w6967;
w6969 <= w230 and not w6968;
w6970 <= w234 and not w6969;
w6971 <= w238 and not w6970;
w6972 <= w242 and not w6971;
w6973 <= w246 and not w6972;
w6974 <= w250 and not w6973;
w6975 <= w254 and not w6974;
w6976 <= w258 and not w6975;
w6977 <= w262 and not w6976;
w6978 <= w266 and not w6977;
w6979 <= w270 and not w6978;
w6980 <= w274 and not w6979;
w6981 <= w278 and not w6980;
w6982 <= w282 and not w6981;
w6983 <= w286 and not w6982;
w6984 <= w290 and not w6983;
w6985 <= w294 and not w6984;
w6986 <= w298 and not w6985;
w6987 <= w302 and not w6986;
w6988 <= w306 and not w6987;
w6989 <= w310 and not w6988;
w6990 <= w314 and not w6989;
w6991 <= w318 and not w6990;
w6992 <= w322 and not w6991;
w6993 <= w326 and not w6992;
w6994 <= w330 and not w6993;
w6995 <= w334 and not w6994;
w6996 <= w1098 and not w6995;
w6997 <= w1100 and not w6996;
w6998 <= w1364 and not w6997;
w6999 <= w345 and not w6998;
w7000 <= w349 and not w6999;
w7001 <= w353 and not w7000;
w7002 <= w357 and not w7001;
w7003 <= w361 and not w7002;
w7004 <= w365 and not w7003;
w7005 <= w369 and not w7004;
w7006 <= w373 and not w7005;
w7007 <= w377 and not w7006;
w7008 <= w381 and not w7007;
w7009 <= w385 and not w7008;
w7010 <= w389 and not w7009;
w7011 <= w393 and not w7010;
w7012 <= w397 and not w7011;
w7013 <= w401 and not w7012;
w7014 <= w405 and not w7013;
w7015 <= w409 and not w7014;
w7016 <= w413 and not w7015;
w7017 <= w417 and not w7016;
w7018 <= w421 and not w7017;
w7019 <= w425 and not w7018;
w7020 <= w429 and not w7019;
w7021 <= w433 and not w7020;
w7022 <= w437 and not w7021;
w7023 <= w441 and not w7022;
w7024 <= w445 and not w7023;
w7025 <= w449 and not w7024;
w7026 <= w453 and not w7025;
w7027 <= w457 and not w7026;
w7028 <= w461 and not w7027;
w7029 <= w465 and not w7028;
w7030 <= w469 and not w7029;
w7031 <= w473 and not w7030;
w7032 <= w477 and not w7031;
w7033 <= w481 and not w7032;
w7034 <= w485 and not w7033;
w7035 <= w489 and not w7034;
w7036 <= w493 and not w7035;
w7037 <= w497 and not w7036;
w7038 <= w501 and not w7037;
w7039 <= w505 and not w7038;
w7040 <= w509 and not w7039;
w7041 <= w513 and not w7040;
w7042 <= w517 and not w7041;
w7043 <= w521 and not w7042;
w7044 <= req(72) and not w523;
w7045 <= not w7043 and w7044;
w7046 <= w532 and not w865;
w7047 <= w537 and not w7046;
w7048 <= w541 and not w7047;
w7049 <= w545 and not w7048;
w7050 <= w549 and not w7049;
w7051 <= w553 and not w7050;
w7052 <= w557 and not w7051;
w7053 <= w561 and not w7052;
w7054 <= w565 and not w7053;
w7055 <= w569 and not w7054;
w7056 <= w573 and not w7055;
w7057 <= w577 and not w7056;
w7058 <= w581 and not w7057;
w7059 <= w585 and not w7058;
w7060 <= w589 and not w7059;
w7061 <= w593 and not w7060;
w7062 <= w597 and not w7061;
w7063 <= w601 and not w7062;
w7064 <= w605 and not w7063;
w7065 <= w609 and not w7064;
w7066 <= w613 and not w7065;
w7067 <= w617 and not w7066;
w7068 <= w621 and not w7067;
w7069 <= w625 and not w7068;
w7070 <= w629 and not w7069;
w7071 <= w633 and not w7070;
w7072 <= w637 and not w7071;
w7073 <= w641 and not w7072;
w7074 <= w645 and not w7073;
w7075 <= w649 and not w7074;
w7076 <= w653 and not w7075;
w7077 <= w657 and not w7076;
w7078 <= w661 and not w7077;
w7079 <= w665 and not w7078;
w7080 <= w669 and not w7079;
w7081 <= w673 and not w7080;
w7082 <= w1188 and not w7081;
w7083 <= w1190 and not w7082;
w7084 <= w1451 and not w7083;
w7085 <= w682 and not w7084;
w7086 <= w686 and not w7085;
w7087 <= w690 and not w7086;
w7088 <= w694 and not w7087;
w7089 <= w698 and not w7088;
w7090 <= w702 and not w7089;
w7091 <= w706 and not w7090;
w7092 <= w710 and not w7091;
w7093 <= w714 and not w7092;
w7094 <= w718 and not w7093;
w7095 <= w722 and not w7094;
w7096 <= w726 and not w7095;
w7097 <= w730 and not w7096;
w7098 <= w734 and not w7097;
w7099 <= w738 and not w7098;
w7100 <= w742 and not w7099;
w7101 <= w746 and not w7100;
w7102 <= w750 and not w7101;
w7103 <= w754 and not w7102;
w7104 <= w758 and not w7103;
w7105 <= w762 and not w7104;
w7106 <= w766 and not w7105;
w7107 <= w770 and not w7106;
w7108 <= w774 and not w7107;
w7109 <= w778 and not w7108;
w7110 <= w782 and not w7109;
w7111 <= w786 and not w7110;
w7112 <= w790 and not w7111;
w7113 <= w794 and not w7112;
w7114 <= w798 and not w7113;
w7115 <= w802 and not w7114;
w7116 <= w806 and not w7115;
w7117 <= w810 and not w7116;
w7118 <= w814 and not w7117;
w7119 <= w818 and not w7118;
w7120 <= w822 and not w7119;
w7121 <= w826 and not w7120;
w7122 <= w830 and not w7121;
w7123 <= w834 and not w7122;
w7124 <= w838 and not w7123;
w7125 <= w842 and not w7124;
w7126 <= w846 and not w7125;
w7127 <= w850 and not w7126;
w7128 <= w854 and not w7127;
w7129 <= w858 and not w7128;
w7130 <= req(73) and not w860;
w7131 <= not w7129 and w7130;
w7132 <= not w197 and w869;
w7133 <= w874 and not w7132;
w7134 <= w878 and not w7133;
w7135 <= w882 and not w7134;
w7136 <= w886 and not w7135;
w7137 <= w890 and not w7136;
w7138 <= w894 and not w7137;
w7139 <= w898 and not w7138;
w7140 <= w902 and not w7139;
w7141 <= w906 and not w7140;
w7142 <= w910 and not w7141;
w7143 <= w914 and not w7142;
w7144 <= w918 and not w7143;
w7145 <= w922 and not w7144;
w7146 <= w926 and not w7145;
w7147 <= w930 and not w7146;
w7148 <= w934 and not w7147;
w7149 <= w938 and not w7148;
w7150 <= w942 and not w7149;
w7151 <= w946 and not w7150;
w7152 <= w950 and not w7151;
w7153 <= w954 and not w7152;
w7154 <= w958 and not w7153;
w7155 <= w962 and not w7154;
w7156 <= w966 and not w7155;
w7157 <= w970 and not w7156;
w7158 <= w974 and not w7157;
w7159 <= w978 and not w7158;
w7160 <= w982 and not w7159;
w7161 <= w986 and not w7160;
w7162 <= w990 and not w7161;
w7163 <= w994 and not w7162;
w7164 <= w998 and not w7163;
w7165 <= w1002 and not w7164;
w7166 <= w1006 and not w7165;
w7167 <= w1010 and not w7166;
w7168 <= w1277 and not w7167;
w7169 <= w6 and not w7168;
w7170 <= w10 and not w7169;
w7171 <= w14 and not w7170;
w7172 <= w18 and not w7171;
w7173 <= w22 and not w7172;
w7174 <= w26 and not w7173;
w7175 <= w30 and not w7174;
w7176 <= w34 and not w7175;
w7177 <= w38 and not w7176;
w7178 <= w42 and not w7177;
w7179 <= w46 and not w7178;
w7180 <= w50 and not w7179;
w7181 <= w54 and not w7180;
w7182 <= w58 and not w7181;
w7183 <= w62 and not w7182;
w7184 <= w66 and not w7183;
w7185 <= w70 and not w7184;
w7186 <= w74 and not w7185;
w7187 <= w78 and not w7186;
w7188 <= w82 and not w7187;
w7189 <= w86 and not w7188;
w7190 <= w90 and not w7189;
w7191 <= w94 and not w7190;
w7192 <= w98 and not w7191;
w7193 <= w102 and not w7192;
w7194 <= w106 and not w7193;
w7195 <= w110 and not w7194;
w7196 <= w114 and not w7195;
w7197 <= w118 and not w7196;
w7198 <= w122 and not w7197;
w7199 <= w126 and not w7198;
w7200 <= w130 and not w7199;
w7201 <= w134 and not w7200;
w7202 <= w138 and not w7201;
w7203 <= w142 and not w7202;
w7204 <= w146 and not w7203;
w7205 <= w150 and not w7204;
w7206 <= w154 and not w7205;
w7207 <= w158 and not w7206;
w7208 <= w162 and not w7207;
w7209 <= w166 and not w7208;
w7210 <= w170 and not w7209;
w7211 <= w174 and not w7210;
w7212 <= w178 and not w7211;
w7213 <= w182 and not w7212;
w7214 <= w186 and not w7213;
w7215 <= w190 and not w7214;
w7216 <= req(74) and not w192;
w7217 <= not w7215 and w7216;
w7218 <= w201 and not w536;
w7219 <= w206 and not w7218;
w7220 <= w210 and not w7219;
w7221 <= w214 and not w7220;
w7222 <= w218 and not w7221;
w7223 <= w222 and not w7222;
w7224 <= w226 and not w7223;
w7225 <= w230 and not w7224;
w7226 <= w234 and not w7225;
w7227 <= w238 and not w7226;
w7228 <= w242 and not w7227;
w7229 <= w246 and not w7228;
w7230 <= w250 and not w7229;
w7231 <= w254 and not w7230;
w7232 <= w258 and not w7231;
w7233 <= w262 and not w7232;
w7234 <= w266 and not w7233;
w7235 <= w270 and not w7234;
w7236 <= w274 and not w7235;
w7237 <= w278 and not w7236;
w7238 <= w282 and not w7237;
w7239 <= w286 and not w7238;
w7240 <= w290 and not w7239;
w7241 <= w294 and not w7240;
w7242 <= w298 and not w7241;
w7243 <= w302 and not w7242;
w7244 <= w306 and not w7243;
w7245 <= w310 and not w7244;
w7246 <= w314 and not w7245;
w7247 <= w318 and not w7246;
w7248 <= w322 and not w7247;
w7249 <= w326 and not w7248;
w7250 <= w330 and not w7249;
w7251 <= w334 and not w7250;
w7252 <= w1098 and not w7251;
w7253 <= w1100 and not w7252;
w7254 <= w1364 and not w7253;
w7255 <= w345 and not w7254;
w7256 <= w349 and not w7255;
w7257 <= w353 and not w7256;
w7258 <= w357 and not w7257;
w7259 <= w361 and not w7258;
w7260 <= w365 and not w7259;
w7261 <= w369 and not w7260;
w7262 <= w373 and not w7261;
w7263 <= w377 and not w7262;
w7264 <= w381 and not w7263;
w7265 <= w385 and not w7264;
w7266 <= w389 and not w7265;
w7267 <= w393 and not w7266;
w7268 <= w397 and not w7267;
w7269 <= w401 and not w7268;
w7270 <= w405 and not w7269;
w7271 <= w409 and not w7270;
w7272 <= w413 and not w7271;
w7273 <= w417 and not w7272;
w7274 <= w421 and not w7273;
w7275 <= w425 and not w7274;
w7276 <= w429 and not w7275;
w7277 <= w433 and not w7276;
w7278 <= w437 and not w7277;
w7279 <= w441 and not w7278;
w7280 <= w445 and not w7279;
w7281 <= w449 and not w7280;
w7282 <= w453 and not w7281;
w7283 <= w457 and not w7282;
w7284 <= w461 and not w7283;
w7285 <= w465 and not w7284;
w7286 <= w469 and not w7285;
w7287 <= w473 and not w7286;
w7288 <= w477 and not w7287;
w7289 <= w481 and not w7288;
w7290 <= w485 and not w7289;
w7291 <= w489 and not w7290;
w7292 <= w493 and not w7291;
w7293 <= w497 and not w7292;
w7294 <= w501 and not w7293;
w7295 <= w505 and not w7294;
w7296 <= w509 and not w7295;
w7297 <= w513 and not w7296;
w7298 <= w517 and not w7297;
w7299 <= w521 and not w7298;
w7300 <= w525 and not w7299;
w7301 <= w529 and not w7300;
w7302 <= req(75) and not w531;
w7303 <= not w7301 and w7302;
w7304 <= w540 and not w873;
w7305 <= w545 and not w7304;
w7306 <= w549 and not w7305;
w7307 <= w553 and not w7306;
w7308 <= w557 and not w7307;
w7309 <= w561 and not w7308;
w7310 <= w565 and not w7309;
w7311 <= w569 and not w7310;
w7312 <= w573 and not w7311;
w7313 <= w577 and not w7312;
w7314 <= w581 and not w7313;
w7315 <= w585 and not w7314;
w7316 <= w589 and not w7315;
w7317 <= w593 and not w7316;
w7318 <= w597 and not w7317;
w7319 <= w601 and not w7318;
w7320 <= w605 and not w7319;
w7321 <= w609 and not w7320;
w7322 <= w613 and not w7321;
w7323 <= w617 and not w7322;
w7324 <= w621 and not w7323;
w7325 <= w625 and not w7324;
w7326 <= w629 and not w7325;
w7327 <= w633 and not w7326;
w7328 <= w637 and not w7327;
w7329 <= w641 and not w7328;
w7330 <= w645 and not w7329;
w7331 <= w649 and not w7330;
w7332 <= w653 and not w7331;
w7333 <= w657 and not w7332;
w7334 <= w661 and not w7333;
w7335 <= w665 and not w7334;
w7336 <= w669 and not w7335;
w7337 <= w673 and not w7336;
w7338 <= w1188 and not w7337;
w7339 <= w1190 and not w7338;
w7340 <= w1451 and not w7339;
w7341 <= w682 and not w7340;
w7342 <= w686 and not w7341;
w7343 <= w690 and not w7342;
w7344 <= w694 and not w7343;
w7345 <= w698 and not w7344;
w7346 <= w702 and not w7345;
w7347 <= w706 and not w7346;
w7348 <= w710 and not w7347;
w7349 <= w714 and not w7348;
w7350 <= w718 and not w7349;
w7351 <= w722 and not w7350;
w7352 <= w726 and not w7351;
w7353 <= w730 and not w7352;
w7354 <= w734 and not w7353;
w7355 <= w738 and not w7354;
w7356 <= w742 and not w7355;
w7357 <= w746 and not w7356;
w7358 <= w750 and not w7357;
w7359 <= w754 and not w7358;
w7360 <= w758 and not w7359;
w7361 <= w762 and not w7360;
w7362 <= w766 and not w7361;
w7363 <= w770 and not w7362;
w7364 <= w774 and not w7363;
w7365 <= w778 and not w7364;
w7366 <= w782 and not w7365;
w7367 <= w786 and not w7366;
w7368 <= w790 and not w7367;
w7369 <= w794 and not w7368;
w7370 <= w798 and not w7369;
w7371 <= w802 and not w7370;
w7372 <= w806 and not w7371;
w7373 <= w810 and not w7372;
w7374 <= w814 and not w7373;
w7375 <= w818 and not w7374;
w7376 <= w822 and not w7375;
w7377 <= w826 and not w7376;
w7378 <= w830 and not w7377;
w7379 <= w834 and not w7378;
w7380 <= w838 and not w7379;
w7381 <= w842 and not w7380;
w7382 <= w846 and not w7381;
w7383 <= w850 and not w7382;
w7384 <= w854 and not w7383;
w7385 <= w858 and not w7384;
w7386 <= w862 and not w7385;
w7387 <= w866 and not w7386;
w7388 <= req(76) and not w868;
w7389 <= not w7387 and w7388;
w7390 <= not w205 and w877;
w7391 <= w882 and not w7390;
w7392 <= w886 and not w7391;
w7393 <= w890 and not w7392;
w7394 <= w894 and not w7393;
w7395 <= w898 and not w7394;
w7396 <= w902 and not w7395;
w7397 <= w906 and not w7396;
w7398 <= w910 and not w7397;
w7399 <= w914 and not w7398;
w7400 <= w918 and not w7399;
w7401 <= w922 and not w7400;
w7402 <= w926 and not w7401;
w7403 <= w930 and not w7402;
w7404 <= w934 and not w7403;
w7405 <= w938 and not w7404;
w7406 <= w942 and not w7405;
w7407 <= w946 and not w7406;
w7408 <= w950 and not w7407;
w7409 <= w954 and not w7408;
w7410 <= w958 and not w7409;
w7411 <= w962 and not w7410;
w7412 <= w966 and not w7411;
w7413 <= w970 and not w7412;
w7414 <= w974 and not w7413;
w7415 <= w978 and not w7414;
w7416 <= w982 and not w7415;
w7417 <= w986 and not w7416;
w7418 <= w990 and not w7417;
w7419 <= w994 and not w7418;
w7420 <= w998 and not w7419;
w7421 <= w1002 and not w7420;
w7422 <= w1006 and not w7421;
w7423 <= w1010 and not w7422;
w7424 <= w1277 and not w7423;
w7425 <= w6 and not w7424;
w7426 <= w10 and not w7425;
w7427 <= w14 and not w7426;
w7428 <= w18 and not w7427;
w7429 <= w22 and not w7428;
w7430 <= w26 and not w7429;
w7431 <= w30 and not w7430;
w7432 <= w34 and not w7431;
w7433 <= w38 and not w7432;
w7434 <= w42 and not w7433;
w7435 <= w46 and not w7434;
w7436 <= w50 and not w7435;
w7437 <= w54 and not w7436;
w7438 <= w58 and not w7437;
w7439 <= w62 and not w7438;
w7440 <= w66 and not w7439;
w7441 <= w70 and not w7440;
w7442 <= w74 and not w7441;
w7443 <= w78 and not w7442;
w7444 <= w82 and not w7443;
w7445 <= w86 and not w7444;
w7446 <= w90 and not w7445;
w7447 <= w94 and not w7446;
w7448 <= w98 and not w7447;
w7449 <= w102 and not w7448;
w7450 <= w106 and not w7449;
w7451 <= w110 and not w7450;
w7452 <= w114 and not w7451;
w7453 <= w118 and not w7452;
w7454 <= w122 and not w7453;
w7455 <= w126 and not w7454;
w7456 <= w130 and not w7455;
w7457 <= w134 and not w7456;
w7458 <= w138 and not w7457;
w7459 <= w142 and not w7458;
w7460 <= w146 and not w7459;
w7461 <= w150 and not w7460;
w7462 <= w154 and not w7461;
w7463 <= w158 and not w7462;
w7464 <= w162 and not w7463;
w7465 <= w166 and not w7464;
w7466 <= w170 and not w7465;
w7467 <= w174 and not w7466;
w7468 <= w178 and not w7467;
w7469 <= w182 and not w7468;
w7470 <= w186 and not w7469;
w7471 <= w190 and not w7470;
w7472 <= w194 and not w7471;
w7473 <= w198 and not w7472;
w7474 <= req(77) and not w200;
w7475 <= not w7473 and w7474;
w7476 <= w209 and not w544;
w7477 <= w214 and not w7476;
w7478 <= w218 and not w7477;
w7479 <= w222 and not w7478;
w7480 <= w226 and not w7479;
w7481 <= w230 and not w7480;
w7482 <= w234 and not w7481;
w7483 <= w238 and not w7482;
w7484 <= w242 and not w7483;
w7485 <= w246 and not w7484;
w7486 <= w250 and not w7485;
w7487 <= w254 and not w7486;
w7488 <= w258 and not w7487;
w7489 <= w262 and not w7488;
w7490 <= w266 and not w7489;
w7491 <= w270 and not w7490;
w7492 <= w274 and not w7491;
w7493 <= w278 and not w7492;
w7494 <= w282 and not w7493;
w7495 <= w286 and not w7494;
w7496 <= w290 and not w7495;
w7497 <= w294 and not w7496;
w7498 <= w298 and not w7497;
w7499 <= w302 and not w7498;
w7500 <= w306 and not w7499;
w7501 <= w310 and not w7500;
w7502 <= w314 and not w7501;
w7503 <= w318 and not w7502;
w7504 <= w322 and not w7503;
w7505 <= w326 and not w7504;
w7506 <= w330 and not w7505;
w7507 <= w334 and not w7506;
w7508 <= w1098 and not w7507;
w7509 <= w1100 and not w7508;
w7510 <= w1364 and not w7509;
w7511 <= w345 and not w7510;
w7512 <= w349 and not w7511;
w7513 <= w353 and not w7512;
w7514 <= w357 and not w7513;
w7515 <= w361 and not w7514;
w7516 <= w365 and not w7515;
w7517 <= w369 and not w7516;
w7518 <= w373 and not w7517;
w7519 <= w377 and not w7518;
w7520 <= w381 and not w7519;
w7521 <= w385 and not w7520;
w7522 <= w389 and not w7521;
w7523 <= w393 and not w7522;
w7524 <= w397 and not w7523;
w7525 <= w401 and not w7524;
w7526 <= w405 and not w7525;
w7527 <= w409 and not w7526;
w7528 <= w413 and not w7527;
w7529 <= w417 and not w7528;
w7530 <= w421 and not w7529;
w7531 <= w425 and not w7530;
w7532 <= w429 and not w7531;
w7533 <= w433 and not w7532;
w7534 <= w437 and not w7533;
w7535 <= w441 and not w7534;
w7536 <= w445 and not w7535;
w7537 <= w449 and not w7536;
w7538 <= w453 and not w7537;
w7539 <= w457 and not w7538;
w7540 <= w461 and not w7539;
w7541 <= w465 and not w7540;
w7542 <= w469 and not w7541;
w7543 <= w473 and not w7542;
w7544 <= w477 and not w7543;
w7545 <= w481 and not w7544;
w7546 <= w485 and not w7545;
w7547 <= w489 and not w7546;
w7548 <= w493 and not w7547;
w7549 <= w497 and not w7548;
w7550 <= w501 and not w7549;
w7551 <= w505 and not w7550;
w7552 <= w509 and not w7551;
w7553 <= w513 and not w7552;
w7554 <= w517 and not w7553;
w7555 <= w521 and not w7554;
w7556 <= w525 and not w7555;
w7557 <= w529 and not w7556;
w7558 <= w533 and not w7557;
w7559 <= w537 and not w7558;
w7560 <= req(78) and not w539;
w7561 <= not w7559 and w7560;
w7562 <= w548 and not w881;
w7563 <= w553 and not w7562;
w7564 <= w557 and not w7563;
w7565 <= w561 and not w7564;
w7566 <= w565 and not w7565;
w7567 <= w569 and not w7566;
w7568 <= w573 and not w7567;
w7569 <= w577 and not w7568;
w7570 <= w581 and not w7569;
w7571 <= w585 and not w7570;
w7572 <= w589 and not w7571;
w7573 <= w593 and not w7572;
w7574 <= w597 and not w7573;
w7575 <= w601 and not w7574;
w7576 <= w605 and not w7575;
w7577 <= w609 and not w7576;
w7578 <= w613 and not w7577;
w7579 <= w617 and not w7578;
w7580 <= w621 and not w7579;
w7581 <= w625 and not w7580;
w7582 <= w629 and not w7581;
w7583 <= w633 and not w7582;
w7584 <= w637 and not w7583;
w7585 <= w641 and not w7584;
w7586 <= w645 and not w7585;
w7587 <= w649 and not w7586;
w7588 <= w653 and not w7587;
w7589 <= w657 and not w7588;
w7590 <= w661 and not w7589;
w7591 <= w665 and not w7590;
w7592 <= w669 and not w7591;
w7593 <= w673 and not w7592;
w7594 <= w1188 and not w7593;
w7595 <= w1190 and not w7594;
w7596 <= w1451 and not w7595;
w7597 <= w682 and not w7596;
w7598 <= w686 and not w7597;
w7599 <= w690 and not w7598;
w7600 <= w694 and not w7599;
w7601 <= w698 and not w7600;
w7602 <= w702 and not w7601;
w7603 <= w706 and not w7602;
w7604 <= w710 and not w7603;
w7605 <= w714 and not w7604;
w7606 <= w718 and not w7605;
w7607 <= w722 and not w7606;
w7608 <= w726 and not w7607;
w7609 <= w730 and not w7608;
w7610 <= w734 and not w7609;
w7611 <= w738 and not w7610;
w7612 <= w742 and not w7611;
w7613 <= w746 and not w7612;
w7614 <= w750 and not w7613;
w7615 <= w754 and not w7614;
w7616 <= w758 and not w7615;
w7617 <= w762 and not w7616;
w7618 <= w766 and not w7617;
w7619 <= w770 and not w7618;
w7620 <= w774 and not w7619;
w7621 <= w778 and not w7620;
w7622 <= w782 and not w7621;
w7623 <= w786 and not w7622;
w7624 <= w790 and not w7623;
w7625 <= w794 and not w7624;
w7626 <= w798 and not w7625;
w7627 <= w802 and not w7626;
w7628 <= w806 and not w7627;
w7629 <= w810 and not w7628;
w7630 <= w814 and not w7629;
w7631 <= w818 and not w7630;
w7632 <= w822 and not w7631;
w7633 <= w826 and not w7632;
w7634 <= w830 and not w7633;
w7635 <= w834 and not w7634;
w7636 <= w838 and not w7635;
w7637 <= w842 and not w7636;
w7638 <= w846 and not w7637;
w7639 <= w850 and not w7638;
w7640 <= w854 and not w7639;
w7641 <= w858 and not w7640;
w7642 <= w862 and not w7641;
w7643 <= w866 and not w7642;
w7644 <= w870 and not w7643;
w7645 <= w874 and not w7644;
w7646 <= req(79) and not w876;
w7647 <= not w7645 and w7646;
w7648 <= not w213 and w885;
w7649 <= w890 and not w7648;
w7650 <= w894 and not w7649;
w7651 <= w898 and not w7650;
w7652 <= w902 and not w7651;
w7653 <= w906 and not w7652;
w7654 <= w910 and not w7653;
w7655 <= w914 and not w7654;
w7656 <= w918 and not w7655;
w7657 <= w922 and not w7656;
w7658 <= w926 and not w7657;
w7659 <= w930 and not w7658;
w7660 <= w934 and not w7659;
w7661 <= w938 and not w7660;
w7662 <= w942 and not w7661;
w7663 <= w946 and not w7662;
w7664 <= w950 and not w7663;
w7665 <= w954 and not w7664;
w7666 <= w958 and not w7665;
w7667 <= w962 and not w7666;
w7668 <= w966 and not w7667;
w7669 <= w970 and not w7668;
w7670 <= w974 and not w7669;
w7671 <= w978 and not w7670;
w7672 <= w982 and not w7671;
w7673 <= w986 and not w7672;
w7674 <= w990 and not w7673;
w7675 <= w994 and not w7674;
w7676 <= w998 and not w7675;
w7677 <= w1002 and not w7676;
w7678 <= w1006 and not w7677;
w7679 <= w1010 and not w7678;
w7680 <= w1277 and not w7679;
w7681 <= w6 and not w7680;
w7682 <= w10 and not w7681;
w7683 <= w14 and not w7682;
w7684 <= w18 and not w7683;
w7685 <= w22 and not w7684;
w7686 <= w26 and not w7685;
w7687 <= w30 and not w7686;
w7688 <= w34 and not w7687;
w7689 <= w38 and not w7688;
w7690 <= w42 and not w7689;
w7691 <= w46 and not w7690;
w7692 <= w50 and not w7691;
w7693 <= w54 and not w7692;
w7694 <= w58 and not w7693;
w7695 <= w62 and not w7694;
w7696 <= w66 and not w7695;
w7697 <= w70 and not w7696;
w7698 <= w74 and not w7697;
w7699 <= w78 and not w7698;
w7700 <= w82 and not w7699;
w7701 <= w86 and not w7700;
w7702 <= w90 and not w7701;
w7703 <= w94 and not w7702;
w7704 <= w98 and not w7703;
w7705 <= w102 and not w7704;
w7706 <= w106 and not w7705;
w7707 <= w110 and not w7706;
w7708 <= w114 and not w7707;
w7709 <= w118 and not w7708;
w7710 <= w122 and not w7709;
w7711 <= w126 and not w7710;
w7712 <= w130 and not w7711;
w7713 <= w134 and not w7712;
w7714 <= w138 and not w7713;
w7715 <= w142 and not w7714;
w7716 <= w146 and not w7715;
w7717 <= w150 and not w7716;
w7718 <= w154 and not w7717;
w7719 <= w158 and not w7718;
w7720 <= w162 and not w7719;
w7721 <= w166 and not w7720;
w7722 <= w170 and not w7721;
w7723 <= w174 and not w7722;
w7724 <= w178 and not w7723;
w7725 <= w182 and not w7724;
w7726 <= w186 and not w7725;
w7727 <= w190 and not w7726;
w7728 <= w194 and not w7727;
w7729 <= w198 and not w7728;
w7730 <= w202 and not w7729;
w7731 <= w206 and not w7730;
w7732 <= req(80) and not w208;
w7733 <= not w7731 and w7732;
w7734 <= w217 and not w552;
w7735 <= w222 and not w7734;
w7736 <= w226 and not w7735;
w7737 <= w230 and not w7736;
w7738 <= w234 and not w7737;
w7739 <= w238 and not w7738;
w7740 <= w242 and not w7739;
w7741 <= w246 and not w7740;
w7742 <= w250 and not w7741;
w7743 <= w254 and not w7742;
w7744 <= w258 and not w7743;
w7745 <= w262 and not w7744;
w7746 <= w266 and not w7745;
w7747 <= w270 and not w7746;
w7748 <= w274 and not w7747;
w7749 <= w278 and not w7748;
w7750 <= w282 and not w7749;
w7751 <= w286 and not w7750;
w7752 <= w290 and not w7751;
w7753 <= w294 and not w7752;
w7754 <= w298 and not w7753;
w7755 <= w302 and not w7754;
w7756 <= w306 and not w7755;
w7757 <= w310 and not w7756;
w7758 <= w314 and not w7757;
w7759 <= w318 and not w7758;
w7760 <= w322 and not w7759;
w7761 <= w326 and not w7760;
w7762 <= w330 and not w7761;
w7763 <= w334 and not w7762;
w7764 <= w1098 and not w7763;
w7765 <= w1100 and not w7764;
w7766 <= w1364 and not w7765;
w7767 <= w345 and not w7766;
w7768 <= w349 and not w7767;
w7769 <= w353 and not w7768;
w7770 <= w357 and not w7769;
w7771 <= w361 and not w7770;
w7772 <= w365 and not w7771;
w7773 <= w369 and not w7772;
w7774 <= w373 and not w7773;
w7775 <= w377 and not w7774;
w7776 <= w381 and not w7775;
w7777 <= w385 and not w7776;
w7778 <= w389 and not w7777;
w7779 <= w393 and not w7778;
w7780 <= w397 and not w7779;
w7781 <= w401 and not w7780;
w7782 <= w405 and not w7781;
w7783 <= w409 and not w7782;
w7784 <= w413 and not w7783;
w7785 <= w417 and not w7784;
w7786 <= w421 and not w7785;
w7787 <= w425 and not w7786;
w7788 <= w429 and not w7787;
w7789 <= w433 and not w7788;
w7790 <= w437 and not w7789;
w7791 <= w441 and not w7790;
w7792 <= w445 and not w7791;
w7793 <= w449 and not w7792;
w7794 <= w453 and not w7793;
w7795 <= w457 and not w7794;
w7796 <= w461 and not w7795;
w7797 <= w465 and not w7796;
w7798 <= w469 and not w7797;
w7799 <= w473 and not w7798;
w7800 <= w477 and not w7799;
w7801 <= w481 and not w7800;
w7802 <= w485 and not w7801;
w7803 <= w489 and not w7802;
w7804 <= w493 and not w7803;
w7805 <= w497 and not w7804;
w7806 <= w501 and not w7805;
w7807 <= w505 and not w7806;
w7808 <= w509 and not w7807;
w7809 <= w513 and not w7808;
w7810 <= w517 and not w7809;
w7811 <= w521 and not w7810;
w7812 <= w525 and not w7811;
w7813 <= w529 and not w7812;
w7814 <= w533 and not w7813;
w7815 <= w537 and not w7814;
w7816 <= w541 and not w7815;
w7817 <= w545 and not w7816;
w7818 <= req(81) and not w547;
w7819 <= not w7817 and w7818;
w7820 <= w556 and not w889;
w7821 <= w561 and not w7820;
w7822 <= w565 and not w7821;
w7823 <= w569 and not w7822;
w7824 <= w573 and not w7823;
w7825 <= w577 and not w7824;
w7826 <= w581 and not w7825;
w7827 <= w585 and not w7826;
w7828 <= w589 and not w7827;
w7829 <= w593 and not w7828;
w7830 <= w597 and not w7829;
w7831 <= w601 and not w7830;
w7832 <= w605 and not w7831;
w7833 <= w609 and not w7832;
w7834 <= w613 and not w7833;
w7835 <= w617 and not w7834;
w7836 <= w621 and not w7835;
w7837 <= w625 and not w7836;
w7838 <= w629 and not w7837;
w7839 <= w633 and not w7838;
w7840 <= w637 and not w7839;
w7841 <= w641 and not w7840;
w7842 <= w645 and not w7841;
w7843 <= w649 and not w7842;
w7844 <= w653 and not w7843;
w7845 <= w657 and not w7844;
w7846 <= w661 and not w7845;
w7847 <= w665 and not w7846;
w7848 <= w669 and not w7847;
w7849 <= w673 and not w7848;
w7850 <= w1188 and not w7849;
w7851 <= w1190 and not w7850;
w7852 <= w1451 and not w7851;
w7853 <= w682 and not w7852;
w7854 <= w686 and not w7853;
w7855 <= w690 and not w7854;
w7856 <= w694 and not w7855;
w7857 <= w698 and not w7856;
w7858 <= w702 and not w7857;
w7859 <= w706 and not w7858;
w7860 <= w710 and not w7859;
w7861 <= w714 and not w7860;
w7862 <= w718 and not w7861;
w7863 <= w722 and not w7862;
w7864 <= w726 and not w7863;
w7865 <= w730 and not w7864;
w7866 <= w734 and not w7865;
w7867 <= w738 and not w7866;
w7868 <= w742 and not w7867;
w7869 <= w746 and not w7868;
w7870 <= w750 and not w7869;
w7871 <= w754 and not w7870;
w7872 <= w758 and not w7871;
w7873 <= w762 and not w7872;
w7874 <= w766 and not w7873;
w7875 <= w770 and not w7874;
w7876 <= w774 and not w7875;
w7877 <= w778 and not w7876;
w7878 <= w782 and not w7877;
w7879 <= w786 and not w7878;
w7880 <= w790 and not w7879;
w7881 <= w794 and not w7880;
w7882 <= w798 and not w7881;
w7883 <= w802 and not w7882;
w7884 <= w806 and not w7883;
w7885 <= w810 and not w7884;
w7886 <= w814 and not w7885;
w7887 <= w818 and not w7886;
w7888 <= w822 and not w7887;
w7889 <= w826 and not w7888;
w7890 <= w830 and not w7889;
w7891 <= w834 and not w7890;
w7892 <= w838 and not w7891;
w7893 <= w842 and not w7892;
w7894 <= w846 and not w7893;
w7895 <= w850 and not w7894;
w7896 <= w854 and not w7895;
w7897 <= w858 and not w7896;
w7898 <= w862 and not w7897;
w7899 <= w866 and not w7898;
w7900 <= w870 and not w7899;
w7901 <= w874 and not w7900;
w7902 <= w878 and not w7901;
w7903 <= w882 and not w7902;
w7904 <= req(82) and not w884;
w7905 <= not w7903 and w7904;
w7906 <= not w221 and w893;
w7907 <= w898 and not w7906;
w7908 <= w902 and not w7907;
w7909 <= w906 and not w7908;
w7910 <= w910 and not w7909;
w7911 <= w914 and not w7910;
w7912 <= w918 and not w7911;
w7913 <= w922 and not w7912;
w7914 <= w926 and not w7913;
w7915 <= w930 and not w7914;
w7916 <= w934 and not w7915;
w7917 <= w938 and not w7916;
w7918 <= w942 and not w7917;
w7919 <= w946 and not w7918;
w7920 <= w950 and not w7919;
w7921 <= w954 and not w7920;
w7922 <= w958 and not w7921;
w7923 <= w962 and not w7922;
w7924 <= w966 and not w7923;
w7925 <= w970 and not w7924;
w7926 <= w974 and not w7925;
w7927 <= w978 and not w7926;
w7928 <= w982 and not w7927;
w7929 <= w986 and not w7928;
w7930 <= w990 and not w7929;
w7931 <= w994 and not w7930;
w7932 <= w998 and not w7931;
w7933 <= w1002 and not w7932;
w7934 <= w1006 and not w7933;
w7935 <= w1010 and not w7934;
w7936 <= w1277 and not w7935;
w7937 <= w6 and not w7936;
w7938 <= w10 and not w7937;
w7939 <= w14 and not w7938;
w7940 <= w18 and not w7939;
w7941 <= w22 and not w7940;
w7942 <= w26 and not w7941;
w7943 <= w30 and not w7942;
w7944 <= w34 and not w7943;
w7945 <= w38 and not w7944;
w7946 <= w42 and not w7945;
w7947 <= w46 and not w7946;
w7948 <= w50 and not w7947;
w7949 <= w54 and not w7948;
w7950 <= w58 and not w7949;
w7951 <= w62 and not w7950;
w7952 <= w66 and not w7951;
w7953 <= w70 and not w7952;
w7954 <= w74 and not w7953;
w7955 <= w78 and not w7954;
w7956 <= w82 and not w7955;
w7957 <= w86 and not w7956;
w7958 <= w90 and not w7957;
w7959 <= w94 and not w7958;
w7960 <= w98 and not w7959;
w7961 <= w102 and not w7960;
w7962 <= w106 and not w7961;
w7963 <= w110 and not w7962;
w7964 <= w114 and not w7963;
w7965 <= w118 and not w7964;
w7966 <= w122 and not w7965;
w7967 <= w126 and not w7966;
w7968 <= w130 and not w7967;
w7969 <= w134 and not w7968;
w7970 <= w138 and not w7969;
w7971 <= w142 and not w7970;
w7972 <= w146 and not w7971;
w7973 <= w150 and not w7972;
w7974 <= w154 and not w7973;
w7975 <= w158 and not w7974;
w7976 <= w162 and not w7975;
w7977 <= w166 and not w7976;
w7978 <= w170 and not w7977;
w7979 <= w174 and not w7978;
w7980 <= w178 and not w7979;
w7981 <= w182 and not w7980;
w7982 <= w186 and not w7981;
w7983 <= w190 and not w7982;
w7984 <= w194 and not w7983;
w7985 <= w198 and not w7984;
w7986 <= w202 and not w7985;
w7987 <= w206 and not w7986;
w7988 <= w210 and not w7987;
w7989 <= w214 and not w7988;
w7990 <= req(83) and not w216;
w7991 <= not w7989 and w7990;
w7992 <= w225 and not w560;
w7993 <= w230 and not w7992;
w7994 <= w234 and not w7993;
w7995 <= w238 and not w7994;
w7996 <= w242 and not w7995;
w7997 <= w246 and not w7996;
w7998 <= w250 and not w7997;
w7999 <= w254 and not w7998;
w8000 <= w258 and not w7999;
w8001 <= w262 and not w8000;
w8002 <= w266 and not w8001;
w8003 <= w270 and not w8002;
w8004 <= w274 and not w8003;
w8005 <= w278 and not w8004;
w8006 <= w282 and not w8005;
w8007 <= w286 and not w8006;
w8008 <= w290 and not w8007;
w8009 <= w294 and not w8008;
w8010 <= w298 and not w8009;
w8011 <= w302 and not w8010;
w8012 <= w306 and not w8011;
w8013 <= w310 and not w8012;
w8014 <= w314 and not w8013;
w8015 <= w318 and not w8014;
w8016 <= w322 and not w8015;
w8017 <= w326 and not w8016;
w8018 <= w330 and not w8017;
w8019 <= w334 and not w8018;
w8020 <= w1098 and not w8019;
w8021 <= w1100 and not w8020;
w8022 <= w1364 and not w8021;
w8023 <= w345 and not w8022;
w8024 <= w349 and not w8023;
w8025 <= w353 and not w8024;
w8026 <= w357 and not w8025;
w8027 <= w361 and not w8026;
w8028 <= w365 and not w8027;
w8029 <= w369 and not w8028;
w8030 <= w373 and not w8029;
w8031 <= w377 and not w8030;
w8032 <= w381 and not w8031;
w8033 <= w385 and not w8032;
w8034 <= w389 and not w8033;
w8035 <= w393 and not w8034;
w8036 <= w397 and not w8035;
w8037 <= w401 and not w8036;
w8038 <= w405 and not w8037;
w8039 <= w409 and not w8038;
w8040 <= w413 and not w8039;
w8041 <= w417 and not w8040;
w8042 <= w421 and not w8041;
w8043 <= w425 and not w8042;
w8044 <= w429 and not w8043;
w8045 <= w433 and not w8044;
w8046 <= w437 and not w8045;
w8047 <= w441 and not w8046;
w8048 <= w445 and not w8047;
w8049 <= w449 and not w8048;
w8050 <= w453 and not w8049;
w8051 <= w457 and not w8050;
w8052 <= w461 and not w8051;
w8053 <= w465 and not w8052;
w8054 <= w469 and not w8053;
w8055 <= w473 and not w8054;
w8056 <= w477 and not w8055;
w8057 <= w481 and not w8056;
w8058 <= w485 and not w8057;
w8059 <= w489 and not w8058;
w8060 <= w493 and not w8059;
w8061 <= w497 and not w8060;
w8062 <= w501 and not w8061;
w8063 <= w505 and not w8062;
w8064 <= w509 and not w8063;
w8065 <= w513 and not w8064;
w8066 <= w517 and not w8065;
w8067 <= w521 and not w8066;
w8068 <= w525 and not w8067;
w8069 <= w529 and not w8068;
w8070 <= w533 and not w8069;
w8071 <= w537 and not w8070;
w8072 <= w541 and not w8071;
w8073 <= w545 and not w8072;
w8074 <= w549 and not w8073;
w8075 <= w553 and not w8074;
w8076 <= req(84) and not w555;
w8077 <= not w8075 and w8076;
w8078 <= w564 and not w897;
w8079 <= w569 and not w8078;
w8080 <= w573 and not w8079;
w8081 <= w577 and not w8080;
w8082 <= w581 and not w8081;
w8083 <= w585 and not w8082;
w8084 <= w589 and not w8083;
w8085 <= w593 and not w8084;
w8086 <= w597 and not w8085;
w8087 <= w601 and not w8086;
w8088 <= w605 and not w8087;
w8089 <= w609 and not w8088;
w8090 <= w613 and not w8089;
w8091 <= w617 and not w8090;
w8092 <= w621 and not w8091;
w8093 <= w625 and not w8092;
w8094 <= w629 and not w8093;
w8095 <= w633 and not w8094;
w8096 <= w637 and not w8095;
w8097 <= w641 and not w8096;
w8098 <= w645 and not w8097;
w8099 <= w649 and not w8098;
w8100 <= w653 and not w8099;
w8101 <= w657 and not w8100;
w8102 <= w661 and not w8101;
w8103 <= w665 and not w8102;
w8104 <= w669 and not w8103;
w8105 <= w673 and not w8104;
w8106 <= w1188 and not w8105;
w8107 <= w1190 and not w8106;
w8108 <= w1451 and not w8107;
w8109 <= w682 and not w8108;
w8110 <= w686 and not w8109;
w8111 <= w690 and not w8110;
w8112 <= w694 and not w8111;
w8113 <= w698 and not w8112;
w8114 <= w702 and not w8113;
w8115 <= w706 and not w8114;
w8116 <= w710 and not w8115;
w8117 <= w714 and not w8116;
w8118 <= w718 and not w8117;
w8119 <= w722 and not w8118;
w8120 <= w726 and not w8119;
w8121 <= w730 and not w8120;
w8122 <= w734 and not w8121;
w8123 <= w738 and not w8122;
w8124 <= w742 and not w8123;
w8125 <= w746 and not w8124;
w8126 <= w750 and not w8125;
w8127 <= w754 and not w8126;
w8128 <= w758 and not w8127;
w8129 <= w762 and not w8128;
w8130 <= w766 and not w8129;
w8131 <= w770 and not w8130;
w8132 <= w774 and not w8131;
w8133 <= w778 and not w8132;
w8134 <= w782 and not w8133;
w8135 <= w786 and not w8134;
w8136 <= w790 and not w8135;
w8137 <= w794 and not w8136;
w8138 <= w798 and not w8137;
w8139 <= w802 and not w8138;
w8140 <= w806 and not w8139;
w8141 <= w810 and not w8140;
w8142 <= w814 and not w8141;
w8143 <= w818 and not w8142;
w8144 <= w822 and not w8143;
w8145 <= w826 and not w8144;
w8146 <= w830 and not w8145;
w8147 <= w834 and not w8146;
w8148 <= w838 and not w8147;
w8149 <= w842 and not w8148;
w8150 <= w846 and not w8149;
w8151 <= w850 and not w8150;
w8152 <= w854 and not w8151;
w8153 <= w858 and not w8152;
w8154 <= w862 and not w8153;
w8155 <= w866 and not w8154;
w8156 <= w870 and not w8155;
w8157 <= w874 and not w8156;
w8158 <= w878 and not w8157;
w8159 <= w882 and not w8158;
w8160 <= w886 and not w8159;
w8161 <= w890 and not w8160;
w8162 <= req(85) and not w892;
w8163 <= not w8161 and w8162;
w8164 <= not w229 and w901;
w8165 <= w906 and not w8164;
w8166 <= w910 and not w8165;
w8167 <= w914 and not w8166;
w8168 <= w918 and not w8167;
w8169 <= w922 and not w8168;
w8170 <= w926 and not w8169;
w8171 <= w930 and not w8170;
w8172 <= w934 and not w8171;
w8173 <= w938 and not w8172;
w8174 <= w942 and not w8173;
w8175 <= w946 and not w8174;
w8176 <= w950 and not w8175;
w8177 <= w954 and not w8176;
w8178 <= w958 and not w8177;
w8179 <= w962 and not w8178;
w8180 <= w966 and not w8179;
w8181 <= w970 and not w8180;
w8182 <= w974 and not w8181;
w8183 <= w978 and not w8182;
w8184 <= w982 and not w8183;
w8185 <= w986 and not w8184;
w8186 <= w990 and not w8185;
w8187 <= w994 and not w8186;
w8188 <= w998 and not w8187;
w8189 <= w1002 and not w8188;
w8190 <= w1006 and not w8189;
w8191 <= w1010 and not w8190;
w8192 <= w1277 and not w8191;
w8193 <= w6 and not w8192;
w8194 <= w10 and not w8193;
w8195 <= w14 and not w8194;
w8196 <= w18 and not w8195;
w8197 <= w22 and not w8196;
w8198 <= w26 and not w8197;
w8199 <= w30 and not w8198;
w8200 <= w34 and not w8199;
w8201 <= w38 and not w8200;
w8202 <= w42 and not w8201;
w8203 <= w46 and not w8202;
w8204 <= w50 and not w8203;
w8205 <= w54 and not w8204;
w8206 <= w58 and not w8205;
w8207 <= w62 and not w8206;
w8208 <= w66 and not w8207;
w8209 <= w70 and not w8208;
w8210 <= w74 and not w8209;
w8211 <= w78 and not w8210;
w8212 <= w82 and not w8211;
w8213 <= w86 and not w8212;
w8214 <= w90 and not w8213;
w8215 <= w94 and not w8214;
w8216 <= w98 and not w8215;
w8217 <= w102 and not w8216;
w8218 <= w106 and not w8217;
w8219 <= w110 and not w8218;
w8220 <= w114 and not w8219;
w8221 <= w118 and not w8220;
w8222 <= w122 and not w8221;
w8223 <= w126 and not w8222;
w8224 <= w130 and not w8223;
w8225 <= w134 and not w8224;
w8226 <= w138 and not w8225;
w8227 <= w142 and not w8226;
w8228 <= w146 and not w8227;
w8229 <= w150 and not w8228;
w8230 <= w154 and not w8229;
w8231 <= w158 and not w8230;
w8232 <= w162 and not w8231;
w8233 <= w166 and not w8232;
w8234 <= w170 and not w8233;
w8235 <= w174 and not w8234;
w8236 <= w178 and not w8235;
w8237 <= w182 and not w8236;
w8238 <= w186 and not w8237;
w8239 <= w190 and not w8238;
w8240 <= w194 and not w8239;
w8241 <= w198 and not w8240;
w8242 <= w202 and not w8241;
w8243 <= w206 and not w8242;
w8244 <= w210 and not w8243;
w8245 <= w214 and not w8244;
w8246 <= w218 and not w8245;
w8247 <= w222 and not w8246;
w8248 <= req(86) and not w224;
w8249 <= not w8247 and w8248;
w8250 <= w233 and not w568;
w8251 <= w238 and not w8250;
w8252 <= w242 and not w8251;
w8253 <= w246 and not w8252;
w8254 <= w250 and not w8253;
w8255 <= w254 and not w8254;
w8256 <= w258 and not w8255;
w8257 <= w262 and not w8256;
w8258 <= w266 and not w8257;
w8259 <= w270 and not w8258;
w8260 <= w274 and not w8259;
w8261 <= w278 and not w8260;
w8262 <= w282 and not w8261;
w8263 <= w286 and not w8262;
w8264 <= w290 and not w8263;
w8265 <= w294 and not w8264;
w8266 <= w298 and not w8265;
w8267 <= w302 and not w8266;
w8268 <= w306 and not w8267;
w8269 <= w310 and not w8268;
w8270 <= w314 and not w8269;
w8271 <= w318 and not w8270;
w8272 <= w322 and not w8271;
w8273 <= w326 and not w8272;
w8274 <= w330 and not w8273;
w8275 <= w334 and not w8274;
w8276 <= w1098 and not w8275;
w8277 <= w1100 and not w8276;
w8278 <= w1364 and not w8277;
w8279 <= w345 and not w8278;
w8280 <= w349 and not w8279;
w8281 <= w353 and not w8280;
w8282 <= w357 and not w8281;
w8283 <= w361 and not w8282;
w8284 <= w365 and not w8283;
w8285 <= w369 and not w8284;
w8286 <= w373 and not w8285;
w8287 <= w377 and not w8286;
w8288 <= w381 and not w8287;
w8289 <= w385 and not w8288;
w8290 <= w389 and not w8289;
w8291 <= w393 and not w8290;
w8292 <= w397 and not w8291;
w8293 <= w401 and not w8292;
w8294 <= w405 and not w8293;
w8295 <= w409 and not w8294;
w8296 <= w413 and not w8295;
w8297 <= w417 and not w8296;
w8298 <= w421 and not w8297;
w8299 <= w425 and not w8298;
w8300 <= w429 and not w8299;
w8301 <= w433 and not w8300;
w8302 <= w437 and not w8301;
w8303 <= w441 and not w8302;
w8304 <= w445 and not w8303;
w8305 <= w449 and not w8304;
w8306 <= w453 and not w8305;
w8307 <= w457 and not w8306;
w8308 <= w461 and not w8307;
w8309 <= w465 and not w8308;
w8310 <= w469 and not w8309;
w8311 <= w473 and not w8310;
w8312 <= w477 and not w8311;
w8313 <= w481 and not w8312;
w8314 <= w485 and not w8313;
w8315 <= w489 and not w8314;
w8316 <= w493 and not w8315;
w8317 <= w497 and not w8316;
w8318 <= w501 and not w8317;
w8319 <= w505 and not w8318;
w8320 <= w509 and not w8319;
w8321 <= w513 and not w8320;
w8322 <= w517 and not w8321;
w8323 <= w521 and not w8322;
w8324 <= w525 and not w8323;
w8325 <= w529 and not w8324;
w8326 <= w533 and not w8325;
w8327 <= w537 and not w8326;
w8328 <= w541 and not w8327;
w8329 <= w545 and not w8328;
w8330 <= w549 and not w8329;
w8331 <= w553 and not w8330;
w8332 <= w557 and not w8331;
w8333 <= w561 and not w8332;
w8334 <= req(87) and not w563;
w8335 <= not w8333 and w8334;
w8336 <= w572 and not w905;
w8337 <= w577 and not w8336;
w8338 <= w581 and not w8337;
w8339 <= w585 and not w8338;
w8340 <= w589 and not w8339;
w8341 <= w593 and not w8340;
w8342 <= w597 and not w8341;
w8343 <= w601 and not w8342;
w8344 <= w605 and not w8343;
w8345 <= w609 and not w8344;
w8346 <= w613 and not w8345;
w8347 <= w617 and not w8346;
w8348 <= w621 and not w8347;
w8349 <= w625 and not w8348;
w8350 <= w629 and not w8349;
w8351 <= w633 and not w8350;
w8352 <= w637 and not w8351;
w8353 <= w641 and not w8352;
w8354 <= w645 and not w8353;
w8355 <= w649 and not w8354;
w8356 <= w653 and not w8355;
w8357 <= w657 and not w8356;
w8358 <= w661 and not w8357;
w8359 <= w665 and not w8358;
w8360 <= w669 and not w8359;
w8361 <= w673 and not w8360;
w8362 <= w1188 and not w8361;
w8363 <= w1190 and not w8362;
w8364 <= w1451 and not w8363;
w8365 <= w682 and not w8364;
w8366 <= w686 and not w8365;
w8367 <= w690 and not w8366;
w8368 <= w694 and not w8367;
w8369 <= w698 and not w8368;
w8370 <= w702 and not w8369;
w8371 <= w706 and not w8370;
w8372 <= w710 and not w8371;
w8373 <= w714 and not w8372;
w8374 <= w718 and not w8373;
w8375 <= w722 and not w8374;
w8376 <= w726 and not w8375;
w8377 <= w730 and not w8376;
w8378 <= w734 and not w8377;
w8379 <= w738 and not w8378;
w8380 <= w742 and not w8379;
w8381 <= w746 and not w8380;
w8382 <= w750 and not w8381;
w8383 <= w754 and not w8382;
w8384 <= w758 and not w8383;
w8385 <= w762 and not w8384;
w8386 <= w766 and not w8385;
w8387 <= w770 and not w8386;
w8388 <= w774 and not w8387;
w8389 <= w778 and not w8388;
w8390 <= w782 and not w8389;
w8391 <= w786 and not w8390;
w8392 <= w790 and not w8391;
w8393 <= w794 and not w8392;
w8394 <= w798 and not w8393;
w8395 <= w802 and not w8394;
w8396 <= w806 and not w8395;
w8397 <= w810 and not w8396;
w8398 <= w814 and not w8397;
w8399 <= w818 and not w8398;
w8400 <= w822 and not w8399;
w8401 <= w826 and not w8400;
w8402 <= w830 and not w8401;
w8403 <= w834 and not w8402;
w8404 <= w838 and not w8403;
w8405 <= w842 and not w8404;
w8406 <= w846 and not w8405;
w8407 <= w850 and not w8406;
w8408 <= w854 and not w8407;
w8409 <= w858 and not w8408;
w8410 <= w862 and not w8409;
w8411 <= w866 and not w8410;
w8412 <= w870 and not w8411;
w8413 <= w874 and not w8412;
w8414 <= w878 and not w8413;
w8415 <= w882 and not w8414;
w8416 <= w886 and not w8415;
w8417 <= w890 and not w8416;
w8418 <= w894 and not w8417;
w8419 <= w898 and not w8418;
w8420 <= req(88) and not w900;
w8421 <= not w8419 and w8420;
w8422 <= not w237 and w909;
w8423 <= w914 and not w8422;
w8424 <= w918 and not w8423;
w8425 <= w922 and not w8424;
w8426 <= w926 and not w8425;
w8427 <= w930 and not w8426;
w8428 <= w934 and not w8427;
w8429 <= w938 and not w8428;
w8430 <= w942 and not w8429;
w8431 <= w946 and not w8430;
w8432 <= w950 and not w8431;
w8433 <= w954 and not w8432;
w8434 <= w958 and not w8433;
w8435 <= w962 and not w8434;
w8436 <= w966 and not w8435;
w8437 <= w970 and not w8436;
w8438 <= w974 and not w8437;
w8439 <= w978 and not w8438;
w8440 <= w982 and not w8439;
w8441 <= w986 and not w8440;
w8442 <= w990 and not w8441;
w8443 <= w994 and not w8442;
w8444 <= w998 and not w8443;
w8445 <= w1002 and not w8444;
w8446 <= w1006 and not w8445;
w8447 <= w1010 and not w8446;
w8448 <= w1277 and not w8447;
w8449 <= w6 and not w8448;
w8450 <= w10 and not w8449;
w8451 <= w14 and not w8450;
w8452 <= w18 and not w8451;
w8453 <= w22 and not w8452;
w8454 <= w26 and not w8453;
w8455 <= w30 and not w8454;
w8456 <= w34 and not w8455;
w8457 <= w38 and not w8456;
w8458 <= w42 and not w8457;
w8459 <= w46 and not w8458;
w8460 <= w50 and not w8459;
w8461 <= w54 and not w8460;
w8462 <= w58 and not w8461;
w8463 <= w62 and not w8462;
w8464 <= w66 and not w8463;
w8465 <= w70 and not w8464;
w8466 <= w74 and not w8465;
w8467 <= w78 and not w8466;
w8468 <= w82 and not w8467;
w8469 <= w86 and not w8468;
w8470 <= w90 and not w8469;
w8471 <= w94 and not w8470;
w8472 <= w98 and not w8471;
w8473 <= w102 and not w8472;
w8474 <= w106 and not w8473;
w8475 <= w110 and not w8474;
w8476 <= w114 and not w8475;
w8477 <= w118 and not w8476;
w8478 <= w122 and not w8477;
w8479 <= w126 and not w8478;
w8480 <= w130 and not w8479;
w8481 <= w134 and not w8480;
w8482 <= w138 and not w8481;
w8483 <= w142 and not w8482;
w8484 <= w146 and not w8483;
w8485 <= w150 and not w8484;
w8486 <= w154 and not w8485;
w8487 <= w158 and not w8486;
w8488 <= w162 and not w8487;
w8489 <= w166 and not w8488;
w8490 <= w170 and not w8489;
w8491 <= w174 and not w8490;
w8492 <= w178 and not w8491;
w8493 <= w182 and not w8492;
w8494 <= w186 and not w8493;
w8495 <= w190 and not w8494;
w8496 <= w194 and not w8495;
w8497 <= w198 and not w8496;
w8498 <= w202 and not w8497;
w8499 <= w206 and not w8498;
w8500 <= w210 and not w8499;
w8501 <= w214 and not w8500;
w8502 <= w218 and not w8501;
w8503 <= w222 and not w8502;
w8504 <= w226 and not w8503;
w8505 <= w230 and not w8504;
w8506 <= req(89) and not w232;
w8507 <= not w8505 and w8506;
w8508 <= w241 and not w576;
w8509 <= w246 and not w8508;
w8510 <= w250 and not w8509;
w8511 <= w254 and not w8510;
w8512 <= w258 and not w8511;
w8513 <= w262 and not w8512;
w8514 <= w266 and not w8513;
w8515 <= w270 and not w8514;
w8516 <= w274 and not w8515;
w8517 <= w278 and not w8516;
w8518 <= w282 and not w8517;
w8519 <= w286 and not w8518;
w8520 <= w290 and not w8519;
w8521 <= w294 and not w8520;
w8522 <= w298 and not w8521;
w8523 <= w302 and not w8522;
w8524 <= w306 and not w8523;
w8525 <= w310 and not w8524;
w8526 <= w314 and not w8525;
w8527 <= w318 and not w8526;
w8528 <= w322 and not w8527;
w8529 <= w326 and not w8528;
w8530 <= w330 and not w8529;
w8531 <= w334 and not w8530;
w8532 <= w1098 and not w8531;
w8533 <= w1100 and not w8532;
w8534 <= w1364 and not w8533;
w8535 <= w345 and not w8534;
w8536 <= w349 and not w8535;
w8537 <= w353 and not w8536;
w8538 <= w357 and not w8537;
w8539 <= w361 and not w8538;
w8540 <= w365 and not w8539;
w8541 <= w369 and not w8540;
w8542 <= w373 and not w8541;
w8543 <= w377 and not w8542;
w8544 <= w381 and not w8543;
w8545 <= w385 and not w8544;
w8546 <= w389 and not w8545;
w8547 <= w393 and not w8546;
w8548 <= w397 and not w8547;
w8549 <= w401 and not w8548;
w8550 <= w405 and not w8549;
w8551 <= w409 and not w8550;
w8552 <= w413 and not w8551;
w8553 <= w417 and not w8552;
w8554 <= w421 and not w8553;
w8555 <= w425 and not w8554;
w8556 <= w429 and not w8555;
w8557 <= w433 and not w8556;
w8558 <= w437 and not w8557;
w8559 <= w441 and not w8558;
w8560 <= w445 and not w8559;
w8561 <= w449 and not w8560;
w8562 <= w453 and not w8561;
w8563 <= w457 and not w8562;
w8564 <= w461 and not w8563;
w8565 <= w465 and not w8564;
w8566 <= w469 and not w8565;
w8567 <= w473 and not w8566;
w8568 <= w477 and not w8567;
w8569 <= w481 and not w8568;
w8570 <= w485 and not w8569;
w8571 <= w489 and not w8570;
w8572 <= w493 and not w8571;
w8573 <= w497 and not w8572;
w8574 <= w501 and not w8573;
w8575 <= w505 and not w8574;
w8576 <= w509 and not w8575;
w8577 <= w513 and not w8576;
w8578 <= w517 and not w8577;
w8579 <= w521 and not w8578;
w8580 <= w525 and not w8579;
w8581 <= w529 and not w8580;
w8582 <= w533 and not w8581;
w8583 <= w537 and not w8582;
w8584 <= w541 and not w8583;
w8585 <= w545 and not w8584;
w8586 <= w549 and not w8585;
w8587 <= w553 and not w8586;
w8588 <= w557 and not w8587;
w8589 <= w561 and not w8588;
w8590 <= w565 and not w8589;
w8591 <= w569 and not w8590;
w8592 <= req(90) and not w571;
w8593 <= not w8591 and w8592;
w8594 <= w580 and not w913;
w8595 <= w585 and not w8594;
w8596 <= w589 and not w8595;
w8597 <= w593 and not w8596;
w8598 <= w597 and not w8597;
w8599 <= w601 and not w8598;
w8600 <= w605 and not w8599;
w8601 <= w609 and not w8600;
w8602 <= w613 and not w8601;
w8603 <= w617 and not w8602;
w8604 <= w621 and not w8603;
w8605 <= w625 and not w8604;
w8606 <= w629 and not w8605;
w8607 <= w633 and not w8606;
w8608 <= w637 and not w8607;
w8609 <= w641 and not w8608;
w8610 <= w645 and not w8609;
w8611 <= w649 and not w8610;
w8612 <= w653 and not w8611;
w8613 <= w657 and not w8612;
w8614 <= w661 and not w8613;
w8615 <= w665 and not w8614;
w8616 <= w669 and not w8615;
w8617 <= w673 and not w8616;
w8618 <= w1188 and not w8617;
w8619 <= w1190 and not w8618;
w8620 <= w1451 and not w8619;
w8621 <= w682 and not w8620;
w8622 <= w686 and not w8621;
w8623 <= w690 and not w8622;
w8624 <= w694 and not w8623;
w8625 <= w698 and not w8624;
w8626 <= w702 and not w8625;
w8627 <= w706 and not w8626;
w8628 <= w710 and not w8627;
w8629 <= w714 and not w8628;
w8630 <= w718 and not w8629;
w8631 <= w722 and not w8630;
w8632 <= w726 and not w8631;
w8633 <= w730 and not w8632;
w8634 <= w734 and not w8633;
w8635 <= w738 and not w8634;
w8636 <= w742 and not w8635;
w8637 <= w746 and not w8636;
w8638 <= w750 and not w8637;
w8639 <= w754 and not w8638;
w8640 <= w758 and not w8639;
w8641 <= w762 and not w8640;
w8642 <= w766 and not w8641;
w8643 <= w770 and not w8642;
w8644 <= w774 and not w8643;
w8645 <= w778 and not w8644;
w8646 <= w782 and not w8645;
w8647 <= w786 and not w8646;
w8648 <= w790 and not w8647;
w8649 <= w794 and not w8648;
w8650 <= w798 and not w8649;
w8651 <= w802 and not w8650;
w8652 <= w806 and not w8651;
w8653 <= w810 and not w8652;
w8654 <= w814 and not w8653;
w8655 <= w818 and not w8654;
w8656 <= w822 and not w8655;
w8657 <= w826 and not w8656;
w8658 <= w830 and not w8657;
w8659 <= w834 and not w8658;
w8660 <= w838 and not w8659;
w8661 <= w842 and not w8660;
w8662 <= w846 and not w8661;
w8663 <= w850 and not w8662;
w8664 <= w854 and not w8663;
w8665 <= w858 and not w8664;
w8666 <= w862 and not w8665;
w8667 <= w866 and not w8666;
w8668 <= w870 and not w8667;
w8669 <= w874 and not w8668;
w8670 <= w878 and not w8669;
w8671 <= w882 and not w8670;
w8672 <= w886 and not w8671;
w8673 <= w890 and not w8672;
w8674 <= w894 and not w8673;
w8675 <= w898 and not w8674;
w8676 <= w902 and not w8675;
w8677 <= w906 and not w8676;
w8678 <= req(91) and not w908;
w8679 <= not w8677 and w8678;
w8680 <= not w245 and w917;
w8681 <= w922 and not w8680;
w8682 <= w926 and not w8681;
w8683 <= w930 and not w8682;
w8684 <= w934 and not w8683;
w8685 <= w938 and not w8684;
w8686 <= w942 and not w8685;
w8687 <= w946 and not w8686;
w8688 <= w950 and not w8687;
w8689 <= w954 and not w8688;
w8690 <= w958 and not w8689;
w8691 <= w962 and not w8690;
w8692 <= w966 and not w8691;
w8693 <= w970 and not w8692;
w8694 <= w974 and not w8693;
w8695 <= w978 and not w8694;
w8696 <= w982 and not w8695;
w8697 <= w986 and not w8696;
w8698 <= w990 and not w8697;
w8699 <= w994 and not w8698;
w8700 <= w998 and not w8699;
w8701 <= w1002 and not w8700;
w8702 <= w1006 and not w8701;
w8703 <= w1010 and not w8702;
w8704 <= w1277 and not w8703;
w8705 <= w6 and not w8704;
w8706 <= w10 and not w8705;
w8707 <= w14 and not w8706;
w8708 <= w18 and not w8707;
w8709 <= w22 and not w8708;
w8710 <= w26 and not w8709;
w8711 <= w30 and not w8710;
w8712 <= w34 and not w8711;
w8713 <= w38 and not w8712;
w8714 <= w42 and not w8713;
w8715 <= w46 and not w8714;
w8716 <= w50 and not w8715;
w8717 <= w54 and not w8716;
w8718 <= w58 and not w8717;
w8719 <= w62 and not w8718;
w8720 <= w66 and not w8719;
w8721 <= w70 and not w8720;
w8722 <= w74 and not w8721;
w8723 <= w78 and not w8722;
w8724 <= w82 and not w8723;
w8725 <= w86 and not w8724;
w8726 <= w90 and not w8725;
w8727 <= w94 and not w8726;
w8728 <= w98 and not w8727;
w8729 <= w102 and not w8728;
w8730 <= w106 and not w8729;
w8731 <= w110 and not w8730;
w8732 <= w114 and not w8731;
w8733 <= w118 and not w8732;
w8734 <= w122 and not w8733;
w8735 <= w126 and not w8734;
w8736 <= w130 and not w8735;
w8737 <= w134 and not w8736;
w8738 <= w138 and not w8737;
w8739 <= w142 and not w8738;
w8740 <= w146 and not w8739;
w8741 <= w150 and not w8740;
w8742 <= w154 and not w8741;
w8743 <= w158 and not w8742;
w8744 <= w162 and not w8743;
w8745 <= w166 and not w8744;
w8746 <= w170 and not w8745;
w8747 <= w174 and not w8746;
w8748 <= w178 and not w8747;
w8749 <= w182 and not w8748;
w8750 <= w186 and not w8749;
w8751 <= w190 and not w8750;
w8752 <= w194 and not w8751;
w8753 <= w198 and not w8752;
w8754 <= w202 and not w8753;
w8755 <= w206 and not w8754;
w8756 <= w210 and not w8755;
w8757 <= w214 and not w8756;
w8758 <= w218 and not w8757;
w8759 <= w222 and not w8758;
w8760 <= w226 and not w8759;
w8761 <= w230 and not w8760;
w8762 <= w234 and not w8761;
w8763 <= w238 and not w8762;
w8764 <= req(92) and not w240;
w8765 <= not w8763 and w8764;
w8766 <= w249 and not w584;
w8767 <= w254 and not w8766;
w8768 <= w258 and not w8767;
w8769 <= w262 and not w8768;
w8770 <= w266 and not w8769;
w8771 <= w270 and not w8770;
w8772 <= w274 and not w8771;
w8773 <= w278 and not w8772;
w8774 <= w282 and not w8773;
w8775 <= w286 and not w8774;
w8776 <= w290 and not w8775;
w8777 <= w294 and not w8776;
w8778 <= w298 and not w8777;
w8779 <= w302 and not w8778;
w8780 <= w306 and not w8779;
w8781 <= w310 and not w8780;
w8782 <= w314 and not w8781;
w8783 <= w318 and not w8782;
w8784 <= w322 and not w8783;
w8785 <= w326 and not w8784;
w8786 <= w330 and not w8785;
w8787 <= w334 and not w8786;
w8788 <= w1098 and not w8787;
w8789 <= w1100 and not w8788;
w8790 <= w1364 and not w8789;
w8791 <= w345 and not w8790;
w8792 <= w349 and not w8791;
w8793 <= w353 and not w8792;
w8794 <= w357 and not w8793;
w8795 <= w361 and not w8794;
w8796 <= w365 and not w8795;
w8797 <= w369 and not w8796;
w8798 <= w373 and not w8797;
w8799 <= w377 and not w8798;
w8800 <= w381 and not w8799;
w8801 <= w385 and not w8800;
w8802 <= w389 and not w8801;
w8803 <= w393 and not w8802;
w8804 <= w397 and not w8803;
w8805 <= w401 and not w8804;
w8806 <= w405 and not w8805;
w8807 <= w409 and not w8806;
w8808 <= w413 and not w8807;
w8809 <= w417 and not w8808;
w8810 <= w421 and not w8809;
w8811 <= w425 and not w8810;
w8812 <= w429 and not w8811;
w8813 <= w433 and not w8812;
w8814 <= w437 and not w8813;
w8815 <= w441 and not w8814;
w8816 <= w445 and not w8815;
w8817 <= w449 and not w8816;
w8818 <= w453 and not w8817;
w8819 <= w457 and not w8818;
w8820 <= w461 and not w8819;
w8821 <= w465 and not w8820;
w8822 <= w469 and not w8821;
w8823 <= w473 and not w8822;
w8824 <= w477 and not w8823;
w8825 <= w481 and not w8824;
w8826 <= w485 and not w8825;
w8827 <= w489 and not w8826;
w8828 <= w493 and not w8827;
w8829 <= w497 and not w8828;
w8830 <= w501 and not w8829;
w8831 <= w505 and not w8830;
w8832 <= w509 and not w8831;
w8833 <= w513 and not w8832;
w8834 <= w517 and not w8833;
w8835 <= w521 and not w8834;
w8836 <= w525 and not w8835;
w8837 <= w529 and not w8836;
w8838 <= w533 and not w8837;
w8839 <= w537 and not w8838;
w8840 <= w541 and not w8839;
w8841 <= w545 and not w8840;
w8842 <= w549 and not w8841;
w8843 <= w553 and not w8842;
w8844 <= w557 and not w8843;
w8845 <= w561 and not w8844;
w8846 <= w565 and not w8845;
w8847 <= w569 and not w8846;
w8848 <= w573 and not w8847;
w8849 <= w577 and not w8848;
w8850 <= req(93) and not w579;
w8851 <= not w8849 and w8850;
w8852 <= w588 and not w921;
w8853 <= w593 and not w8852;
w8854 <= w597 and not w8853;
w8855 <= w601 and not w8854;
w8856 <= w605 and not w8855;
w8857 <= w609 and not w8856;
w8858 <= w613 and not w8857;
w8859 <= w617 and not w8858;
w8860 <= w621 and not w8859;
w8861 <= w625 and not w8860;
w8862 <= w629 and not w8861;
w8863 <= w633 and not w8862;
w8864 <= w637 and not w8863;
w8865 <= w641 and not w8864;
w8866 <= w645 and not w8865;
w8867 <= w649 and not w8866;
w8868 <= w653 and not w8867;
w8869 <= w657 and not w8868;
w8870 <= w661 and not w8869;
w8871 <= w665 and not w8870;
w8872 <= w669 and not w8871;
w8873 <= w673 and not w8872;
w8874 <= w1188 and not w8873;
w8875 <= w1190 and not w8874;
w8876 <= w1451 and not w8875;
w8877 <= w682 and not w8876;
w8878 <= w686 and not w8877;
w8879 <= w690 and not w8878;
w8880 <= w694 and not w8879;
w8881 <= w698 and not w8880;
w8882 <= w702 and not w8881;
w8883 <= w706 and not w8882;
w8884 <= w710 and not w8883;
w8885 <= w714 and not w8884;
w8886 <= w718 and not w8885;
w8887 <= w722 and not w8886;
w8888 <= w726 and not w8887;
w8889 <= w730 and not w8888;
w8890 <= w734 and not w8889;
w8891 <= w738 and not w8890;
w8892 <= w742 and not w8891;
w8893 <= w746 and not w8892;
w8894 <= w750 and not w8893;
w8895 <= w754 and not w8894;
w8896 <= w758 and not w8895;
w8897 <= w762 and not w8896;
w8898 <= w766 and not w8897;
w8899 <= w770 and not w8898;
w8900 <= w774 and not w8899;
w8901 <= w778 and not w8900;
w8902 <= w782 and not w8901;
w8903 <= w786 and not w8902;
w8904 <= w790 and not w8903;
w8905 <= w794 and not w8904;
w8906 <= w798 and not w8905;
w8907 <= w802 and not w8906;
w8908 <= w806 and not w8907;
w8909 <= w810 and not w8908;
w8910 <= w814 and not w8909;
w8911 <= w818 and not w8910;
w8912 <= w822 and not w8911;
w8913 <= w826 and not w8912;
w8914 <= w830 and not w8913;
w8915 <= w834 and not w8914;
w8916 <= w838 and not w8915;
w8917 <= w842 and not w8916;
w8918 <= w846 and not w8917;
w8919 <= w850 and not w8918;
w8920 <= w854 and not w8919;
w8921 <= w858 and not w8920;
w8922 <= w862 and not w8921;
w8923 <= w866 and not w8922;
w8924 <= w870 and not w8923;
w8925 <= w874 and not w8924;
w8926 <= w878 and not w8925;
w8927 <= w882 and not w8926;
w8928 <= w886 and not w8927;
w8929 <= w890 and not w8928;
w8930 <= w894 and not w8929;
w8931 <= w898 and not w8930;
w8932 <= w902 and not w8931;
w8933 <= w906 and not w8932;
w8934 <= w910 and not w8933;
w8935 <= w914 and not w8934;
w8936 <= req(94) and not w916;
w8937 <= not w8935 and w8936;
w8938 <= not w253 and w925;
w8939 <= w930 and not w8938;
w8940 <= w934 and not w8939;
w8941 <= w938 and not w8940;
w8942 <= w942 and not w8941;
w8943 <= w946 and not w8942;
w8944 <= w950 and not w8943;
w8945 <= w954 and not w8944;
w8946 <= w958 and not w8945;
w8947 <= w962 and not w8946;
w8948 <= w966 and not w8947;
w8949 <= w970 and not w8948;
w8950 <= w974 and not w8949;
w8951 <= w978 and not w8950;
w8952 <= w982 and not w8951;
w8953 <= w986 and not w8952;
w8954 <= w990 and not w8953;
w8955 <= w994 and not w8954;
w8956 <= w998 and not w8955;
w8957 <= w1002 and not w8956;
w8958 <= w1006 and not w8957;
w8959 <= w1010 and not w8958;
w8960 <= w1277 and not w8959;
w8961 <= w6 and not w8960;
w8962 <= w10 and not w8961;
w8963 <= w14 and not w8962;
w8964 <= w18 and not w8963;
w8965 <= w22 and not w8964;
w8966 <= w26 and not w8965;
w8967 <= w30 and not w8966;
w8968 <= w34 and not w8967;
w8969 <= w38 and not w8968;
w8970 <= w42 and not w8969;
w8971 <= w46 and not w8970;
w8972 <= w50 and not w8971;
w8973 <= w54 and not w8972;
w8974 <= w58 and not w8973;
w8975 <= w62 and not w8974;
w8976 <= w66 and not w8975;
w8977 <= w70 and not w8976;
w8978 <= w74 and not w8977;
w8979 <= w78 and not w8978;
w8980 <= w82 and not w8979;
w8981 <= w86 and not w8980;
w8982 <= w90 and not w8981;
w8983 <= w94 and not w8982;
w8984 <= w98 and not w8983;
w8985 <= w102 and not w8984;
w8986 <= w106 and not w8985;
w8987 <= w110 and not w8986;
w8988 <= w114 and not w8987;
w8989 <= w118 and not w8988;
w8990 <= w122 and not w8989;
w8991 <= w126 and not w8990;
w8992 <= w130 and not w8991;
w8993 <= w134 and not w8992;
w8994 <= w138 and not w8993;
w8995 <= w142 and not w8994;
w8996 <= w146 and not w8995;
w8997 <= w150 and not w8996;
w8998 <= w154 and not w8997;
w8999 <= w158 and not w8998;
w9000 <= w162 and not w8999;
w9001 <= w166 and not w9000;
w9002 <= w170 and not w9001;
w9003 <= w174 and not w9002;
w9004 <= w178 and not w9003;
w9005 <= w182 and not w9004;
w9006 <= w186 and not w9005;
w9007 <= w190 and not w9006;
w9008 <= w194 and not w9007;
w9009 <= w198 and not w9008;
w9010 <= w202 and not w9009;
w9011 <= w206 and not w9010;
w9012 <= w210 and not w9011;
w9013 <= w214 and not w9012;
w9014 <= w218 and not w9013;
w9015 <= w222 and not w9014;
w9016 <= w226 and not w9015;
w9017 <= w230 and not w9016;
w9018 <= w234 and not w9017;
w9019 <= w238 and not w9018;
w9020 <= w242 and not w9019;
w9021 <= w246 and not w9020;
w9022 <= req(95) and not w248;
w9023 <= not w9021 and w9022;
w9024 <= w257 and not w592;
w9025 <= w262 and not w9024;
w9026 <= w266 and not w9025;
w9027 <= w270 and not w9026;
w9028 <= w274 and not w9027;
w9029 <= w278 and not w9028;
w9030 <= w282 and not w9029;
w9031 <= w286 and not w9030;
w9032 <= w290 and not w9031;
w9033 <= w294 and not w9032;
w9034 <= w298 and not w9033;
w9035 <= w302 and not w9034;
w9036 <= w306 and not w9035;
w9037 <= w310 and not w9036;
w9038 <= w314 and not w9037;
w9039 <= w318 and not w9038;
w9040 <= w322 and not w9039;
w9041 <= w326 and not w9040;
w9042 <= w330 and not w9041;
w9043 <= w334 and not w9042;
w9044 <= w1098 and not w9043;
w9045 <= w1100 and not w9044;
w9046 <= w1364 and not w9045;
w9047 <= w345 and not w9046;
w9048 <= w349 and not w9047;
w9049 <= w353 and not w9048;
w9050 <= w357 and not w9049;
w9051 <= w361 and not w9050;
w9052 <= w365 and not w9051;
w9053 <= w369 and not w9052;
w9054 <= w373 and not w9053;
w9055 <= w377 and not w9054;
w9056 <= w381 and not w9055;
w9057 <= w385 and not w9056;
w9058 <= w389 and not w9057;
w9059 <= w393 and not w9058;
w9060 <= w397 and not w9059;
w9061 <= w401 and not w9060;
w9062 <= w405 and not w9061;
w9063 <= w409 and not w9062;
w9064 <= w413 and not w9063;
w9065 <= w417 and not w9064;
w9066 <= w421 and not w9065;
w9067 <= w425 and not w9066;
w9068 <= w429 and not w9067;
w9069 <= w433 and not w9068;
w9070 <= w437 and not w9069;
w9071 <= w441 and not w9070;
w9072 <= w445 and not w9071;
w9073 <= w449 and not w9072;
w9074 <= w453 and not w9073;
w9075 <= w457 and not w9074;
w9076 <= w461 and not w9075;
w9077 <= w465 and not w9076;
w9078 <= w469 and not w9077;
w9079 <= w473 and not w9078;
w9080 <= w477 and not w9079;
w9081 <= w481 and not w9080;
w9082 <= w485 and not w9081;
w9083 <= w489 and not w9082;
w9084 <= w493 and not w9083;
w9085 <= w497 and not w9084;
w9086 <= w501 and not w9085;
w9087 <= w505 and not w9086;
w9088 <= w509 and not w9087;
w9089 <= w513 and not w9088;
w9090 <= w517 and not w9089;
w9091 <= w521 and not w9090;
w9092 <= w525 and not w9091;
w9093 <= w529 and not w9092;
w9094 <= w533 and not w9093;
w9095 <= w537 and not w9094;
w9096 <= w541 and not w9095;
w9097 <= w545 and not w9096;
w9098 <= w549 and not w9097;
w9099 <= w553 and not w9098;
w9100 <= w557 and not w9099;
w9101 <= w561 and not w9100;
w9102 <= w565 and not w9101;
w9103 <= w569 and not w9102;
w9104 <= w573 and not w9103;
w9105 <= w577 and not w9104;
w9106 <= w581 and not w9105;
w9107 <= w585 and not w9106;
w9108 <= req(96) and not w587;
w9109 <= not w9107 and w9108;
w9110 <= w596 and not w929;
w9111 <= w601 and not w9110;
w9112 <= w605 and not w9111;
w9113 <= w609 and not w9112;
w9114 <= w613 and not w9113;
w9115 <= w617 and not w9114;
w9116 <= w621 and not w9115;
w9117 <= w625 and not w9116;
w9118 <= w629 and not w9117;
w9119 <= w633 and not w9118;
w9120 <= w637 and not w9119;
w9121 <= w641 and not w9120;
w9122 <= w645 and not w9121;
w9123 <= w649 and not w9122;
w9124 <= w653 and not w9123;
w9125 <= w657 and not w9124;
w9126 <= w661 and not w9125;
w9127 <= w665 and not w9126;
w9128 <= w669 and not w9127;
w9129 <= w673 and not w9128;
w9130 <= w1188 and not w9129;
w9131 <= w1190 and not w9130;
w9132 <= w1451 and not w9131;
w9133 <= w682 and not w9132;
w9134 <= w686 and not w9133;
w9135 <= w690 and not w9134;
w9136 <= w694 and not w9135;
w9137 <= w698 and not w9136;
w9138 <= w702 and not w9137;
w9139 <= w706 and not w9138;
w9140 <= w710 and not w9139;
w9141 <= w714 and not w9140;
w9142 <= w718 and not w9141;
w9143 <= w722 and not w9142;
w9144 <= w726 and not w9143;
w9145 <= w730 and not w9144;
w9146 <= w734 and not w9145;
w9147 <= w738 and not w9146;
w9148 <= w742 and not w9147;
w9149 <= w746 and not w9148;
w9150 <= w750 and not w9149;
w9151 <= w754 and not w9150;
w9152 <= w758 and not w9151;
w9153 <= w762 and not w9152;
w9154 <= w766 and not w9153;
w9155 <= w770 and not w9154;
w9156 <= w774 and not w9155;
w9157 <= w778 and not w9156;
w9158 <= w782 and not w9157;
w9159 <= w786 and not w9158;
w9160 <= w790 and not w9159;
w9161 <= w794 and not w9160;
w9162 <= w798 and not w9161;
w9163 <= w802 and not w9162;
w9164 <= w806 and not w9163;
w9165 <= w810 and not w9164;
w9166 <= w814 and not w9165;
w9167 <= w818 and not w9166;
w9168 <= w822 and not w9167;
w9169 <= w826 and not w9168;
w9170 <= w830 and not w9169;
w9171 <= w834 and not w9170;
w9172 <= w838 and not w9171;
w9173 <= w842 and not w9172;
w9174 <= w846 and not w9173;
w9175 <= w850 and not w9174;
w9176 <= w854 and not w9175;
w9177 <= w858 and not w9176;
w9178 <= w862 and not w9177;
w9179 <= w866 and not w9178;
w9180 <= w870 and not w9179;
w9181 <= w874 and not w9180;
w9182 <= w878 and not w9181;
w9183 <= w882 and not w9182;
w9184 <= w886 and not w9183;
w9185 <= w890 and not w9184;
w9186 <= w894 and not w9185;
w9187 <= w898 and not w9186;
w9188 <= w902 and not w9187;
w9189 <= w906 and not w9188;
w9190 <= w910 and not w9189;
w9191 <= w914 and not w9190;
w9192 <= w918 and not w9191;
w9193 <= w922 and not w9192;
w9194 <= req(97) and not w924;
w9195 <= not w9193 and w9194;
w9196 <= not w261 and w933;
w9197 <= w938 and not w9196;
w9198 <= w942 and not w9197;
w9199 <= w946 and not w9198;
w9200 <= w950 and not w9199;
w9201 <= w954 and not w9200;
w9202 <= w958 and not w9201;
w9203 <= w962 and not w9202;
w9204 <= w966 and not w9203;
w9205 <= w970 and not w9204;
w9206 <= w974 and not w9205;
w9207 <= w978 and not w9206;
w9208 <= w982 and not w9207;
w9209 <= w986 and not w9208;
w9210 <= w990 and not w9209;
w9211 <= w994 and not w9210;
w9212 <= w998 and not w9211;
w9213 <= w1002 and not w9212;
w9214 <= w1006 and not w9213;
w9215 <= w1010 and not w9214;
w9216 <= w1277 and not w9215;
w9217 <= w6 and not w9216;
w9218 <= w10 and not w9217;
w9219 <= w14 and not w9218;
w9220 <= w18 and not w9219;
w9221 <= w22 and not w9220;
w9222 <= w26 and not w9221;
w9223 <= w30 and not w9222;
w9224 <= w34 and not w9223;
w9225 <= w38 and not w9224;
w9226 <= w42 and not w9225;
w9227 <= w46 and not w9226;
w9228 <= w50 and not w9227;
w9229 <= w54 and not w9228;
w9230 <= w58 and not w9229;
w9231 <= w62 and not w9230;
w9232 <= w66 and not w9231;
w9233 <= w70 and not w9232;
w9234 <= w74 and not w9233;
w9235 <= w78 and not w9234;
w9236 <= w82 and not w9235;
w9237 <= w86 and not w9236;
w9238 <= w90 and not w9237;
w9239 <= w94 and not w9238;
w9240 <= w98 and not w9239;
w9241 <= w102 and not w9240;
w9242 <= w106 and not w9241;
w9243 <= w110 and not w9242;
w9244 <= w114 and not w9243;
w9245 <= w118 and not w9244;
w9246 <= w122 and not w9245;
w9247 <= w126 and not w9246;
w9248 <= w130 and not w9247;
w9249 <= w134 and not w9248;
w9250 <= w138 and not w9249;
w9251 <= w142 and not w9250;
w9252 <= w146 and not w9251;
w9253 <= w150 and not w9252;
w9254 <= w154 and not w9253;
w9255 <= w158 and not w9254;
w9256 <= w162 and not w9255;
w9257 <= w166 and not w9256;
w9258 <= w170 and not w9257;
w9259 <= w174 and not w9258;
w9260 <= w178 and not w9259;
w9261 <= w182 and not w9260;
w9262 <= w186 and not w9261;
w9263 <= w190 and not w9262;
w9264 <= w194 and not w9263;
w9265 <= w198 and not w9264;
w9266 <= w202 and not w9265;
w9267 <= w206 and not w9266;
w9268 <= w210 and not w9267;
w9269 <= w214 and not w9268;
w9270 <= w218 and not w9269;
w9271 <= w222 and not w9270;
w9272 <= w226 and not w9271;
w9273 <= w230 and not w9272;
w9274 <= w234 and not w9273;
w9275 <= w238 and not w9274;
w9276 <= w242 and not w9275;
w9277 <= w246 and not w9276;
w9278 <= w250 and not w9277;
w9279 <= w254 and not w9278;
w9280 <= req(98) and not w256;
w9281 <= not w9279 and w9280;
w9282 <= w265 and not w600;
w9283 <= w270 and not w9282;
w9284 <= w274 and not w9283;
w9285 <= w278 and not w9284;
w9286 <= w282 and not w9285;
w9287 <= w286 and not w9286;
w9288 <= w290 and not w9287;
w9289 <= w294 and not w9288;
w9290 <= w298 and not w9289;
w9291 <= w302 and not w9290;
w9292 <= w306 and not w9291;
w9293 <= w310 and not w9292;
w9294 <= w314 and not w9293;
w9295 <= w318 and not w9294;
w9296 <= w322 and not w9295;
w9297 <= w326 and not w9296;
w9298 <= w330 and not w9297;
w9299 <= w334 and not w9298;
w9300 <= w1098 and not w9299;
w9301 <= w1100 and not w9300;
w9302 <= w1364 and not w9301;
w9303 <= w345 and not w9302;
w9304 <= w349 and not w9303;
w9305 <= w353 and not w9304;
w9306 <= w357 and not w9305;
w9307 <= w361 and not w9306;
w9308 <= w365 and not w9307;
w9309 <= w369 and not w9308;
w9310 <= w373 and not w9309;
w9311 <= w377 and not w9310;
w9312 <= w381 and not w9311;
w9313 <= w385 and not w9312;
w9314 <= w389 and not w9313;
w9315 <= w393 and not w9314;
w9316 <= w397 and not w9315;
w9317 <= w401 and not w9316;
w9318 <= w405 and not w9317;
w9319 <= w409 and not w9318;
w9320 <= w413 and not w9319;
w9321 <= w417 and not w9320;
w9322 <= w421 and not w9321;
w9323 <= w425 and not w9322;
w9324 <= w429 and not w9323;
w9325 <= w433 and not w9324;
w9326 <= w437 and not w9325;
w9327 <= w441 and not w9326;
w9328 <= w445 and not w9327;
w9329 <= w449 and not w9328;
w9330 <= w453 and not w9329;
w9331 <= w457 and not w9330;
w9332 <= w461 and not w9331;
w9333 <= w465 and not w9332;
w9334 <= w469 and not w9333;
w9335 <= w473 and not w9334;
w9336 <= w477 and not w9335;
w9337 <= w481 and not w9336;
w9338 <= w485 and not w9337;
w9339 <= w489 and not w9338;
w9340 <= w493 and not w9339;
w9341 <= w497 and not w9340;
w9342 <= w501 and not w9341;
w9343 <= w505 and not w9342;
w9344 <= w509 and not w9343;
w9345 <= w513 and not w9344;
w9346 <= w517 and not w9345;
w9347 <= w521 and not w9346;
w9348 <= w525 and not w9347;
w9349 <= w529 and not w9348;
w9350 <= w533 and not w9349;
w9351 <= w537 and not w9350;
w9352 <= w541 and not w9351;
w9353 <= w545 and not w9352;
w9354 <= w549 and not w9353;
w9355 <= w553 and not w9354;
w9356 <= w557 and not w9355;
w9357 <= w561 and not w9356;
w9358 <= w565 and not w9357;
w9359 <= w569 and not w9358;
w9360 <= w573 and not w9359;
w9361 <= w577 and not w9360;
w9362 <= w581 and not w9361;
w9363 <= w585 and not w9362;
w9364 <= w589 and not w9363;
w9365 <= w593 and not w9364;
w9366 <= req(99) and not w595;
w9367 <= not w9365 and w9366;
w9368 <= w604 and not w937;
w9369 <= w609 and not w9368;
w9370 <= w613 and not w9369;
w9371 <= w617 and not w9370;
w9372 <= w621 and not w9371;
w9373 <= w625 and not w9372;
w9374 <= w629 and not w9373;
w9375 <= w633 and not w9374;
w9376 <= w637 and not w9375;
w9377 <= w641 and not w9376;
w9378 <= w645 and not w9377;
w9379 <= w649 and not w9378;
w9380 <= w653 and not w9379;
w9381 <= w657 and not w9380;
w9382 <= w661 and not w9381;
w9383 <= w665 and not w9382;
w9384 <= w669 and not w9383;
w9385 <= w673 and not w9384;
w9386 <= w1188 and not w9385;
w9387 <= w1190 and not w9386;
w9388 <= w1451 and not w9387;
w9389 <= w682 and not w9388;
w9390 <= w686 and not w9389;
w9391 <= w690 and not w9390;
w9392 <= w694 and not w9391;
w9393 <= w698 and not w9392;
w9394 <= w702 and not w9393;
w9395 <= w706 and not w9394;
w9396 <= w710 and not w9395;
w9397 <= w714 and not w9396;
w9398 <= w718 and not w9397;
w9399 <= w722 and not w9398;
w9400 <= w726 and not w9399;
w9401 <= w730 and not w9400;
w9402 <= w734 and not w9401;
w9403 <= w738 and not w9402;
w9404 <= w742 and not w9403;
w9405 <= w746 and not w9404;
w9406 <= w750 and not w9405;
w9407 <= w754 and not w9406;
w9408 <= w758 and not w9407;
w9409 <= w762 and not w9408;
w9410 <= w766 and not w9409;
w9411 <= w770 and not w9410;
w9412 <= w774 and not w9411;
w9413 <= w778 and not w9412;
w9414 <= w782 and not w9413;
w9415 <= w786 and not w9414;
w9416 <= w790 and not w9415;
w9417 <= w794 and not w9416;
w9418 <= w798 and not w9417;
w9419 <= w802 and not w9418;
w9420 <= w806 and not w9419;
w9421 <= w810 and not w9420;
w9422 <= w814 and not w9421;
w9423 <= w818 and not w9422;
w9424 <= w822 and not w9423;
w9425 <= w826 and not w9424;
w9426 <= w830 and not w9425;
w9427 <= w834 and not w9426;
w9428 <= w838 and not w9427;
w9429 <= w842 and not w9428;
w9430 <= w846 and not w9429;
w9431 <= w850 and not w9430;
w9432 <= w854 and not w9431;
w9433 <= w858 and not w9432;
w9434 <= w862 and not w9433;
w9435 <= w866 and not w9434;
w9436 <= w870 and not w9435;
w9437 <= w874 and not w9436;
w9438 <= w878 and not w9437;
w9439 <= w882 and not w9438;
w9440 <= w886 and not w9439;
w9441 <= w890 and not w9440;
w9442 <= w894 and not w9441;
w9443 <= w898 and not w9442;
w9444 <= w902 and not w9443;
w9445 <= w906 and not w9444;
w9446 <= w910 and not w9445;
w9447 <= w914 and not w9446;
w9448 <= w918 and not w9447;
w9449 <= w922 and not w9448;
w9450 <= w926 and not w9449;
w9451 <= w930 and not w9450;
w9452 <= req(100) and not w932;
w9453 <= not w9451 and w9452;
w9454 <= not w269 and w941;
w9455 <= w946 and not w9454;
w9456 <= w950 and not w9455;
w9457 <= w954 and not w9456;
w9458 <= w958 and not w9457;
w9459 <= w962 and not w9458;
w9460 <= w966 and not w9459;
w9461 <= w970 and not w9460;
w9462 <= w974 and not w9461;
w9463 <= w978 and not w9462;
w9464 <= w982 and not w9463;
w9465 <= w986 and not w9464;
w9466 <= w990 and not w9465;
w9467 <= w994 and not w9466;
w9468 <= w998 and not w9467;
w9469 <= w1002 and not w9468;
w9470 <= w1006 and not w9469;
w9471 <= w1010 and not w9470;
w9472 <= w1277 and not w9471;
w9473 <= w6 and not w9472;
w9474 <= w10 and not w9473;
w9475 <= w14 and not w9474;
w9476 <= w18 and not w9475;
w9477 <= w22 and not w9476;
w9478 <= w26 and not w9477;
w9479 <= w30 and not w9478;
w9480 <= w34 and not w9479;
w9481 <= w38 and not w9480;
w9482 <= w42 and not w9481;
w9483 <= w46 and not w9482;
w9484 <= w50 and not w9483;
w9485 <= w54 and not w9484;
w9486 <= w58 and not w9485;
w9487 <= w62 and not w9486;
w9488 <= w66 and not w9487;
w9489 <= w70 and not w9488;
w9490 <= w74 and not w9489;
w9491 <= w78 and not w9490;
w9492 <= w82 and not w9491;
w9493 <= w86 and not w9492;
w9494 <= w90 and not w9493;
w9495 <= w94 and not w9494;
w9496 <= w98 and not w9495;
w9497 <= w102 and not w9496;
w9498 <= w106 and not w9497;
w9499 <= w110 and not w9498;
w9500 <= w114 and not w9499;
w9501 <= w118 and not w9500;
w9502 <= w122 and not w9501;
w9503 <= w126 and not w9502;
w9504 <= w130 and not w9503;
w9505 <= w134 and not w9504;
w9506 <= w138 and not w9505;
w9507 <= w142 and not w9506;
w9508 <= w146 and not w9507;
w9509 <= w150 and not w9508;
w9510 <= w154 and not w9509;
w9511 <= w158 and not w9510;
w9512 <= w162 and not w9511;
w9513 <= w166 and not w9512;
w9514 <= w170 and not w9513;
w9515 <= w174 and not w9514;
w9516 <= w178 and not w9515;
w9517 <= w182 and not w9516;
w9518 <= w186 and not w9517;
w9519 <= w190 and not w9518;
w9520 <= w194 and not w9519;
w9521 <= w198 and not w9520;
w9522 <= w202 and not w9521;
w9523 <= w206 and not w9522;
w9524 <= w210 and not w9523;
w9525 <= w214 and not w9524;
w9526 <= w218 and not w9525;
w9527 <= w222 and not w9526;
w9528 <= w226 and not w9527;
w9529 <= w230 and not w9528;
w9530 <= w234 and not w9529;
w9531 <= w238 and not w9530;
w9532 <= w242 and not w9531;
w9533 <= w246 and not w9532;
w9534 <= w250 and not w9533;
w9535 <= w254 and not w9534;
w9536 <= w258 and not w9535;
w9537 <= w262 and not w9536;
w9538 <= req(101) and not w264;
w9539 <= not w9537 and w9538;
w9540 <= w273 and not w608;
w9541 <= w278 and not w9540;
w9542 <= w282 and not w9541;
w9543 <= w286 and not w9542;
w9544 <= w290 and not w9543;
w9545 <= w294 and not w9544;
w9546 <= w298 and not w9545;
w9547 <= w302 and not w9546;
w9548 <= w306 and not w9547;
w9549 <= w310 and not w9548;
w9550 <= w314 and not w9549;
w9551 <= w318 and not w9550;
w9552 <= w322 and not w9551;
w9553 <= w326 and not w9552;
w9554 <= w330 and not w9553;
w9555 <= w334 and not w9554;
w9556 <= w1098 and not w9555;
w9557 <= w1100 and not w9556;
w9558 <= w1364 and not w9557;
w9559 <= w345 and not w9558;
w9560 <= w349 and not w9559;
w9561 <= w353 and not w9560;
w9562 <= w357 and not w9561;
w9563 <= w361 and not w9562;
w9564 <= w365 and not w9563;
w9565 <= w369 and not w9564;
w9566 <= w373 and not w9565;
w9567 <= w377 and not w9566;
w9568 <= w381 and not w9567;
w9569 <= w385 and not w9568;
w9570 <= w389 and not w9569;
w9571 <= w393 and not w9570;
w9572 <= w397 and not w9571;
w9573 <= w401 and not w9572;
w9574 <= w405 and not w9573;
w9575 <= w409 and not w9574;
w9576 <= w413 and not w9575;
w9577 <= w417 and not w9576;
w9578 <= w421 and not w9577;
w9579 <= w425 and not w9578;
w9580 <= w429 and not w9579;
w9581 <= w433 and not w9580;
w9582 <= w437 and not w9581;
w9583 <= w441 and not w9582;
w9584 <= w445 and not w9583;
w9585 <= w449 and not w9584;
w9586 <= w453 and not w9585;
w9587 <= w457 and not w9586;
w9588 <= w461 and not w9587;
w9589 <= w465 and not w9588;
w9590 <= w469 and not w9589;
w9591 <= w473 and not w9590;
w9592 <= w477 and not w9591;
w9593 <= w481 and not w9592;
w9594 <= w485 and not w9593;
w9595 <= w489 and not w9594;
w9596 <= w493 and not w9595;
w9597 <= w497 and not w9596;
w9598 <= w501 and not w9597;
w9599 <= w505 and not w9598;
w9600 <= w509 and not w9599;
w9601 <= w513 and not w9600;
w9602 <= w517 and not w9601;
w9603 <= w521 and not w9602;
w9604 <= w525 and not w9603;
w9605 <= w529 and not w9604;
w9606 <= w533 and not w9605;
w9607 <= w537 and not w9606;
w9608 <= w541 and not w9607;
w9609 <= w545 and not w9608;
w9610 <= w549 and not w9609;
w9611 <= w553 and not w9610;
w9612 <= w557 and not w9611;
w9613 <= w561 and not w9612;
w9614 <= w565 and not w9613;
w9615 <= w569 and not w9614;
w9616 <= w573 and not w9615;
w9617 <= w577 and not w9616;
w9618 <= w581 and not w9617;
w9619 <= w585 and not w9618;
w9620 <= w589 and not w9619;
w9621 <= w593 and not w9620;
w9622 <= w597 and not w9621;
w9623 <= w601 and not w9622;
w9624 <= req(102) and not w603;
w9625 <= not w9623 and w9624;
w9626 <= w612 and not w945;
w9627 <= w617 and not w9626;
w9628 <= w621 and not w9627;
w9629 <= w625 and not w9628;
w9630 <= w629 and not w9629;
w9631 <= w633 and not w9630;
w9632 <= w637 and not w9631;
w9633 <= w641 and not w9632;
w9634 <= w645 and not w9633;
w9635 <= w649 and not w9634;
w9636 <= w653 and not w9635;
w9637 <= w657 and not w9636;
w9638 <= w661 and not w9637;
w9639 <= w665 and not w9638;
w9640 <= w669 and not w9639;
w9641 <= w673 and not w9640;
w9642 <= w1188 and not w9641;
w9643 <= w1190 and not w9642;
w9644 <= w1451 and not w9643;
w9645 <= w682 and not w9644;
w9646 <= w686 and not w9645;
w9647 <= w690 and not w9646;
w9648 <= w694 and not w9647;
w9649 <= w698 and not w9648;
w9650 <= w702 and not w9649;
w9651 <= w706 and not w9650;
w9652 <= w710 and not w9651;
w9653 <= w714 and not w9652;
w9654 <= w718 and not w9653;
w9655 <= w722 and not w9654;
w9656 <= w726 and not w9655;
w9657 <= w730 and not w9656;
w9658 <= w734 and not w9657;
w9659 <= w738 and not w9658;
w9660 <= w742 and not w9659;
w9661 <= w746 and not w9660;
w9662 <= w750 and not w9661;
w9663 <= w754 and not w9662;
w9664 <= w758 and not w9663;
w9665 <= w762 and not w9664;
w9666 <= w766 and not w9665;
w9667 <= w770 and not w9666;
w9668 <= w774 and not w9667;
w9669 <= w778 and not w9668;
w9670 <= w782 and not w9669;
w9671 <= w786 and not w9670;
w9672 <= w790 and not w9671;
w9673 <= w794 and not w9672;
w9674 <= w798 and not w9673;
w9675 <= w802 and not w9674;
w9676 <= w806 and not w9675;
w9677 <= w810 and not w9676;
w9678 <= w814 and not w9677;
w9679 <= w818 and not w9678;
w9680 <= w822 and not w9679;
w9681 <= w826 and not w9680;
w9682 <= w830 and not w9681;
w9683 <= w834 and not w9682;
w9684 <= w838 and not w9683;
w9685 <= w842 and not w9684;
w9686 <= w846 and not w9685;
w9687 <= w850 and not w9686;
w9688 <= w854 and not w9687;
w9689 <= w858 and not w9688;
w9690 <= w862 and not w9689;
w9691 <= w866 and not w9690;
w9692 <= w870 and not w9691;
w9693 <= w874 and not w9692;
w9694 <= w878 and not w9693;
w9695 <= w882 and not w9694;
w9696 <= w886 and not w9695;
w9697 <= w890 and not w9696;
w9698 <= w894 and not w9697;
w9699 <= w898 and not w9698;
w9700 <= w902 and not w9699;
w9701 <= w906 and not w9700;
w9702 <= w910 and not w9701;
w9703 <= w914 and not w9702;
w9704 <= w918 and not w9703;
w9705 <= w922 and not w9704;
w9706 <= w926 and not w9705;
w9707 <= w930 and not w9706;
w9708 <= w934 and not w9707;
w9709 <= w938 and not w9708;
w9710 <= req(103) and not w940;
w9711 <= not w9709 and w9710;
w9712 <= not w277 and w949;
w9713 <= w954 and not w9712;
w9714 <= w958 and not w9713;
w9715 <= w962 and not w9714;
w9716 <= w966 and not w9715;
w9717 <= w970 and not w9716;
w9718 <= w974 and not w9717;
w9719 <= w978 and not w9718;
w9720 <= w982 and not w9719;
w9721 <= w986 and not w9720;
w9722 <= w990 and not w9721;
w9723 <= w994 and not w9722;
w9724 <= w998 and not w9723;
w9725 <= w1002 and not w9724;
w9726 <= w1006 and not w9725;
w9727 <= w1010 and not w9726;
w9728 <= w1277 and not w9727;
w9729 <= w6 and not w9728;
w9730 <= w10 and not w9729;
w9731 <= w14 and not w9730;
w9732 <= w18 and not w9731;
w9733 <= w22 and not w9732;
w9734 <= w26 and not w9733;
w9735 <= w30 and not w9734;
w9736 <= w34 and not w9735;
w9737 <= w38 and not w9736;
w9738 <= w42 and not w9737;
w9739 <= w46 and not w9738;
w9740 <= w50 and not w9739;
w9741 <= w54 and not w9740;
w9742 <= w58 and not w9741;
w9743 <= w62 and not w9742;
w9744 <= w66 and not w9743;
w9745 <= w70 and not w9744;
w9746 <= w74 and not w9745;
w9747 <= w78 and not w9746;
w9748 <= w82 and not w9747;
w9749 <= w86 and not w9748;
w9750 <= w90 and not w9749;
w9751 <= w94 and not w9750;
w9752 <= w98 and not w9751;
w9753 <= w102 and not w9752;
w9754 <= w106 and not w9753;
w9755 <= w110 and not w9754;
w9756 <= w114 and not w9755;
w9757 <= w118 and not w9756;
w9758 <= w122 and not w9757;
w9759 <= w126 and not w9758;
w9760 <= w130 and not w9759;
w9761 <= w134 and not w9760;
w9762 <= w138 and not w9761;
w9763 <= w142 and not w9762;
w9764 <= w146 and not w9763;
w9765 <= w150 and not w9764;
w9766 <= w154 and not w9765;
w9767 <= w158 and not w9766;
w9768 <= w162 and not w9767;
w9769 <= w166 and not w9768;
w9770 <= w170 and not w9769;
w9771 <= w174 and not w9770;
w9772 <= w178 and not w9771;
w9773 <= w182 and not w9772;
w9774 <= w186 and not w9773;
w9775 <= w190 and not w9774;
w9776 <= w194 and not w9775;
w9777 <= w198 and not w9776;
w9778 <= w202 and not w9777;
w9779 <= w206 and not w9778;
w9780 <= w210 and not w9779;
w9781 <= w214 and not w9780;
w9782 <= w218 and not w9781;
w9783 <= w222 and not w9782;
w9784 <= w226 and not w9783;
w9785 <= w230 and not w9784;
w9786 <= w234 and not w9785;
w9787 <= w238 and not w9786;
w9788 <= w242 and not w9787;
w9789 <= w246 and not w9788;
w9790 <= w250 and not w9789;
w9791 <= w254 and not w9790;
w9792 <= w258 and not w9791;
w9793 <= w262 and not w9792;
w9794 <= w266 and not w9793;
w9795 <= w270 and not w9794;
w9796 <= req(104) and not w272;
w9797 <= not w9795 and w9796;
w9798 <= w281 and not w616;
w9799 <= w286 and not w9798;
w9800 <= w290 and not w9799;
w9801 <= w294 and not w9800;
w9802 <= w298 and not w9801;
w9803 <= w302 and not w9802;
w9804 <= w306 and not w9803;
w9805 <= w310 and not w9804;
w9806 <= w314 and not w9805;
w9807 <= w318 and not w9806;
w9808 <= w322 and not w9807;
w9809 <= w326 and not w9808;
w9810 <= w330 and not w9809;
w9811 <= w334 and not w9810;
w9812 <= w1098 and not w9811;
w9813 <= w1100 and not w9812;
w9814 <= w1364 and not w9813;
w9815 <= w345 and not w9814;
w9816 <= w349 and not w9815;
w9817 <= w353 and not w9816;
w9818 <= w357 and not w9817;
w9819 <= w361 and not w9818;
w9820 <= w365 and not w9819;
w9821 <= w369 and not w9820;
w9822 <= w373 and not w9821;
w9823 <= w377 and not w9822;
w9824 <= w381 and not w9823;
w9825 <= w385 and not w9824;
w9826 <= w389 and not w9825;
w9827 <= w393 and not w9826;
w9828 <= w397 and not w9827;
w9829 <= w401 and not w9828;
w9830 <= w405 and not w9829;
w9831 <= w409 and not w9830;
w9832 <= w413 and not w9831;
w9833 <= w417 and not w9832;
w9834 <= w421 and not w9833;
w9835 <= w425 and not w9834;
w9836 <= w429 and not w9835;
w9837 <= w433 and not w9836;
w9838 <= w437 and not w9837;
w9839 <= w441 and not w9838;
w9840 <= w445 and not w9839;
w9841 <= w449 and not w9840;
w9842 <= w453 and not w9841;
w9843 <= w457 and not w9842;
w9844 <= w461 and not w9843;
w9845 <= w465 and not w9844;
w9846 <= w469 and not w9845;
w9847 <= w473 and not w9846;
w9848 <= w477 and not w9847;
w9849 <= w481 and not w9848;
w9850 <= w485 and not w9849;
w9851 <= w489 and not w9850;
w9852 <= w493 and not w9851;
w9853 <= w497 and not w9852;
w9854 <= w501 and not w9853;
w9855 <= w505 and not w9854;
w9856 <= w509 and not w9855;
w9857 <= w513 and not w9856;
w9858 <= w517 and not w9857;
w9859 <= w521 and not w9858;
w9860 <= w525 and not w9859;
w9861 <= w529 and not w9860;
w9862 <= w533 and not w9861;
w9863 <= w537 and not w9862;
w9864 <= w541 and not w9863;
w9865 <= w545 and not w9864;
w9866 <= w549 and not w9865;
w9867 <= w553 and not w9866;
w9868 <= w557 and not w9867;
w9869 <= w561 and not w9868;
w9870 <= w565 and not w9869;
w9871 <= w569 and not w9870;
w9872 <= w573 and not w9871;
w9873 <= w577 and not w9872;
w9874 <= w581 and not w9873;
w9875 <= w585 and not w9874;
w9876 <= w589 and not w9875;
w9877 <= w593 and not w9876;
w9878 <= w597 and not w9877;
w9879 <= w601 and not w9878;
w9880 <= w605 and not w9879;
w9881 <= w609 and not w9880;
w9882 <= req(105) and not w611;
w9883 <= not w9881 and w9882;
w9884 <= w620 and not w953;
w9885 <= w625 and not w9884;
w9886 <= w629 and not w9885;
w9887 <= w633 and not w9886;
w9888 <= w637 and not w9887;
w9889 <= w641 and not w9888;
w9890 <= w645 and not w9889;
w9891 <= w649 and not w9890;
w9892 <= w653 and not w9891;
w9893 <= w657 and not w9892;
w9894 <= w661 and not w9893;
w9895 <= w665 and not w9894;
w9896 <= w669 and not w9895;
w9897 <= w673 and not w9896;
w9898 <= w1188 and not w9897;
w9899 <= w1190 and not w9898;
w9900 <= w1451 and not w9899;
w9901 <= w682 and not w9900;
w9902 <= w686 and not w9901;
w9903 <= w690 and not w9902;
w9904 <= w694 and not w9903;
w9905 <= w698 and not w9904;
w9906 <= w702 and not w9905;
w9907 <= w706 and not w9906;
w9908 <= w710 and not w9907;
w9909 <= w714 and not w9908;
w9910 <= w718 and not w9909;
w9911 <= w722 and not w9910;
w9912 <= w726 and not w9911;
w9913 <= w730 and not w9912;
w9914 <= w734 and not w9913;
w9915 <= w738 and not w9914;
w9916 <= w742 and not w9915;
w9917 <= w746 and not w9916;
w9918 <= w750 and not w9917;
w9919 <= w754 and not w9918;
w9920 <= w758 and not w9919;
w9921 <= w762 and not w9920;
w9922 <= w766 and not w9921;
w9923 <= w770 and not w9922;
w9924 <= w774 and not w9923;
w9925 <= w778 and not w9924;
w9926 <= w782 and not w9925;
w9927 <= w786 and not w9926;
w9928 <= w790 and not w9927;
w9929 <= w794 and not w9928;
w9930 <= w798 and not w9929;
w9931 <= w802 and not w9930;
w9932 <= w806 and not w9931;
w9933 <= w810 and not w9932;
w9934 <= w814 and not w9933;
w9935 <= w818 and not w9934;
w9936 <= w822 and not w9935;
w9937 <= w826 and not w9936;
w9938 <= w830 and not w9937;
w9939 <= w834 and not w9938;
w9940 <= w838 and not w9939;
w9941 <= w842 and not w9940;
w9942 <= w846 and not w9941;
w9943 <= w850 and not w9942;
w9944 <= w854 and not w9943;
w9945 <= w858 and not w9944;
w9946 <= w862 and not w9945;
w9947 <= w866 and not w9946;
w9948 <= w870 and not w9947;
w9949 <= w874 and not w9948;
w9950 <= w878 and not w9949;
w9951 <= w882 and not w9950;
w9952 <= w886 and not w9951;
w9953 <= w890 and not w9952;
w9954 <= w894 and not w9953;
w9955 <= w898 and not w9954;
w9956 <= w902 and not w9955;
w9957 <= w906 and not w9956;
w9958 <= w910 and not w9957;
w9959 <= w914 and not w9958;
w9960 <= w918 and not w9959;
w9961 <= w922 and not w9960;
w9962 <= w926 and not w9961;
w9963 <= w930 and not w9962;
w9964 <= w934 and not w9963;
w9965 <= w938 and not w9964;
w9966 <= w942 and not w9965;
w9967 <= w946 and not w9966;
w9968 <= req(106) and not w948;
w9969 <= not w9967 and w9968;
w9970 <= not w285 and w957;
w9971 <= w962 and not w9970;
w9972 <= w966 and not w9971;
w9973 <= w970 and not w9972;
w9974 <= w974 and not w9973;
w9975 <= w978 and not w9974;
w9976 <= w982 and not w9975;
w9977 <= w986 and not w9976;
w9978 <= w990 and not w9977;
w9979 <= w994 and not w9978;
w9980 <= w998 and not w9979;
w9981 <= w1002 and not w9980;
w9982 <= w1006 and not w9981;
w9983 <= w1010 and not w9982;
w9984 <= w1277 and not w9983;
w9985 <= w6 and not w9984;
w9986 <= w10 and not w9985;
w9987 <= w14 and not w9986;
w9988 <= w18 and not w9987;
w9989 <= w22 and not w9988;
w9990 <= w26 and not w9989;
w9991 <= w30 and not w9990;
w9992 <= w34 and not w9991;
w9993 <= w38 and not w9992;
w9994 <= w42 and not w9993;
w9995 <= w46 and not w9994;
w9996 <= w50 and not w9995;
w9997 <= w54 and not w9996;
w9998 <= w58 and not w9997;
w9999 <= w62 and not w9998;
w10000 <= w66 and not w9999;
w10001 <= w70 and not w10000;
w10002 <= w74 and not w10001;
w10003 <= w78 and not w10002;
w10004 <= w82 and not w10003;
w10005 <= w86 and not w10004;
w10006 <= w90 and not w10005;
w10007 <= w94 and not w10006;
w10008 <= w98 and not w10007;
w10009 <= w102 and not w10008;
w10010 <= w106 and not w10009;
w10011 <= w110 and not w10010;
w10012 <= w114 and not w10011;
w10013 <= w118 and not w10012;
w10014 <= w122 and not w10013;
w10015 <= w126 and not w10014;
w10016 <= w130 and not w10015;
w10017 <= w134 and not w10016;
w10018 <= w138 and not w10017;
w10019 <= w142 and not w10018;
w10020 <= w146 and not w10019;
w10021 <= w150 and not w10020;
w10022 <= w154 and not w10021;
w10023 <= w158 and not w10022;
w10024 <= w162 and not w10023;
w10025 <= w166 and not w10024;
w10026 <= w170 and not w10025;
w10027 <= w174 and not w10026;
w10028 <= w178 and not w10027;
w10029 <= w182 and not w10028;
w10030 <= w186 and not w10029;
w10031 <= w190 and not w10030;
w10032 <= w194 and not w10031;
w10033 <= w198 and not w10032;
w10034 <= w202 and not w10033;
w10035 <= w206 and not w10034;
w10036 <= w210 and not w10035;
w10037 <= w214 and not w10036;
w10038 <= w218 and not w10037;
w10039 <= w222 and not w10038;
w10040 <= w226 and not w10039;
w10041 <= w230 and not w10040;
w10042 <= w234 and not w10041;
w10043 <= w238 and not w10042;
w10044 <= w242 and not w10043;
w10045 <= w246 and not w10044;
w10046 <= w250 and not w10045;
w10047 <= w254 and not w10046;
w10048 <= w258 and not w10047;
w10049 <= w262 and not w10048;
w10050 <= w266 and not w10049;
w10051 <= w270 and not w10050;
w10052 <= w274 and not w10051;
w10053 <= w278 and not w10052;
w10054 <= req(107) and not w280;
w10055 <= not w10053 and w10054;
w10056 <= w289 and not w624;
w10057 <= w294 and not w10056;
w10058 <= w298 and not w10057;
w10059 <= w302 and not w10058;
w10060 <= w306 and not w10059;
w10061 <= w310 and not w10060;
w10062 <= w314 and not w10061;
w10063 <= w318 and not w10062;
w10064 <= w322 and not w10063;
w10065 <= w326 and not w10064;
w10066 <= w330 and not w10065;
w10067 <= w334 and not w10066;
w10068 <= w1098 and not w10067;
w10069 <= w1100 and not w10068;
w10070 <= w1364 and not w10069;
w10071 <= w345 and not w10070;
w10072 <= w349 and not w10071;
w10073 <= w353 and not w10072;
w10074 <= w357 and not w10073;
w10075 <= w361 and not w10074;
w10076 <= w365 and not w10075;
w10077 <= w369 and not w10076;
w10078 <= w373 and not w10077;
w10079 <= w377 and not w10078;
w10080 <= w381 and not w10079;
w10081 <= w385 and not w10080;
w10082 <= w389 and not w10081;
w10083 <= w393 and not w10082;
w10084 <= w397 and not w10083;
w10085 <= w401 and not w10084;
w10086 <= w405 and not w10085;
w10087 <= w409 and not w10086;
w10088 <= w413 and not w10087;
w10089 <= w417 and not w10088;
w10090 <= w421 and not w10089;
w10091 <= w425 and not w10090;
w10092 <= w429 and not w10091;
w10093 <= w433 and not w10092;
w10094 <= w437 and not w10093;
w10095 <= w441 and not w10094;
w10096 <= w445 and not w10095;
w10097 <= w449 and not w10096;
w10098 <= w453 and not w10097;
w10099 <= w457 and not w10098;
w10100 <= w461 and not w10099;
w10101 <= w465 and not w10100;
w10102 <= w469 and not w10101;
w10103 <= w473 and not w10102;
w10104 <= w477 and not w10103;
w10105 <= w481 and not w10104;
w10106 <= w485 and not w10105;
w10107 <= w489 and not w10106;
w10108 <= w493 and not w10107;
w10109 <= w497 and not w10108;
w10110 <= w501 and not w10109;
w10111 <= w505 and not w10110;
w10112 <= w509 and not w10111;
w10113 <= w513 and not w10112;
w10114 <= w517 and not w10113;
w10115 <= w521 and not w10114;
w10116 <= w525 and not w10115;
w10117 <= w529 and not w10116;
w10118 <= w533 and not w10117;
w10119 <= w537 and not w10118;
w10120 <= w541 and not w10119;
w10121 <= w545 and not w10120;
w10122 <= w549 and not w10121;
w10123 <= w553 and not w10122;
w10124 <= w557 and not w10123;
w10125 <= w561 and not w10124;
w10126 <= w565 and not w10125;
w10127 <= w569 and not w10126;
w10128 <= w573 and not w10127;
w10129 <= w577 and not w10128;
w10130 <= w581 and not w10129;
w10131 <= w585 and not w10130;
w10132 <= w589 and not w10131;
w10133 <= w593 and not w10132;
w10134 <= w597 and not w10133;
w10135 <= w601 and not w10134;
w10136 <= w605 and not w10135;
w10137 <= w609 and not w10136;
w10138 <= w613 and not w10137;
w10139 <= w617 and not w10138;
w10140 <= req(108) and not w619;
w10141 <= not w10139 and w10140;
w10142 <= w628 and not w961;
w10143 <= w633 and not w10142;
w10144 <= w637 and not w10143;
w10145 <= w641 and not w10144;
w10146 <= w645 and not w10145;
w10147 <= w649 and not w10146;
w10148 <= w653 and not w10147;
w10149 <= w657 and not w10148;
w10150 <= w661 and not w10149;
w10151 <= w665 and not w10150;
w10152 <= w669 and not w10151;
w10153 <= w673 and not w10152;
w10154 <= w1188 and not w10153;
w10155 <= w1190 and not w10154;
w10156 <= w1451 and not w10155;
w10157 <= w682 and not w10156;
w10158 <= w686 and not w10157;
w10159 <= w690 and not w10158;
w10160 <= w694 and not w10159;
w10161 <= w698 and not w10160;
w10162 <= w702 and not w10161;
w10163 <= w706 and not w10162;
w10164 <= w710 and not w10163;
w10165 <= w714 and not w10164;
w10166 <= w718 and not w10165;
w10167 <= w722 and not w10166;
w10168 <= w726 and not w10167;
w10169 <= w730 and not w10168;
w10170 <= w734 and not w10169;
w10171 <= w738 and not w10170;
w10172 <= w742 and not w10171;
w10173 <= w746 and not w10172;
w10174 <= w750 and not w10173;
w10175 <= w754 and not w10174;
w10176 <= w758 and not w10175;
w10177 <= w762 and not w10176;
w10178 <= w766 and not w10177;
w10179 <= w770 and not w10178;
w10180 <= w774 and not w10179;
w10181 <= w778 and not w10180;
w10182 <= w782 and not w10181;
w10183 <= w786 and not w10182;
w10184 <= w790 and not w10183;
w10185 <= w794 and not w10184;
w10186 <= w798 and not w10185;
w10187 <= w802 and not w10186;
w10188 <= w806 and not w10187;
w10189 <= w810 and not w10188;
w10190 <= w814 and not w10189;
w10191 <= w818 and not w10190;
w10192 <= w822 and not w10191;
w10193 <= w826 and not w10192;
w10194 <= w830 and not w10193;
w10195 <= w834 and not w10194;
w10196 <= w838 and not w10195;
w10197 <= w842 and not w10196;
w10198 <= w846 and not w10197;
w10199 <= w850 and not w10198;
w10200 <= w854 and not w10199;
w10201 <= w858 and not w10200;
w10202 <= w862 and not w10201;
w10203 <= w866 and not w10202;
w10204 <= w870 and not w10203;
w10205 <= w874 and not w10204;
w10206 <= w878 and not w10205;
w10207 <= w882 and not w10206;
w10208 <= w886 and not w10207;
w10209 <= w890 and not w10208;
w10210 <= w894 and not w10209;
w10211 <= w898 and not w10210;
w10212 <= w902 and not w10211;
w10213 <= w906 and not w10212;
w10214 <= w910 and not w10213;
w10215 <= w914 and not w10214;
w10216 <= w918 and not w10215;
w10217 <= w922 and not w10216;
w10218 <= w926 and not w10217;
w10219 <= w930 and not w10218;
w10220 <= w934 and not w10219;
w10221 <= w938 and not w10220;
w10222 <= w942 and not w10221;
w10223 <= w946 and not w10222;
w10224 <= w950 and not w10223;
w10225 <= w954 and not w10224;
w10226 <= req(109) and not w956;
w10227 <= not w10225 and w10226;
w10228 <= not w293 and w965;
w10229 <= w970 and not w10228;
w10230 <= w974 and not w10229;
w10231 <= w978 and not w10230;
w10232 <= w982 and not w10231;
w10233 <= w986 and not w10232;
w10234 <= w990 and not w10233;
w10235 <= w994 and not w10234;
w10236 <= w998 and not w10235;
w10237 <= w1002 and not w10236;
w10238 <= w1006 and not w10237;
w10239 <= w1010 and not w10238;
w10240 <= w1277 and not w10239;
w10241 <= w6 and not w10240;
w10242 <= w10 and not w10241;
w10243 <= w14 and not w10242;
w10244 <= w18 and not w10243;
w10245 <= w22 and not w10244;
w10246 <= w26 and not w10245;
w10247 <= w30 and not w10246;
w10248 <= w34 and not w10247;
w10249 <= w38 and not w10248;
w10250 <= w42 and not w10249;
w10251 <= w46 and not w10250;
w10252 <= w50 and not w10251;
w10253 <= w54 and not w10252;
w10254 <= w58 and not w10253;
w10255 <= w62 and not w10254;
w10256 <= w66 and not w10255;
w10257 <= w70 and not w10256;
w10258 <= w74 and not w10257;
w10259 <= w78 and not w10258;
w10260 <= w82 and not w10259;
w10261 <= w86 and not w10260;
w10262 <= w90 and not w10261;
w10263 <= w94 and not w10262;
w10264 <= w98 and not w10263;
w10265 <= w102 and not w10264;
w10266 <= w106 and not w10265;
w10267 <= w110 and not w10266;
w10268 <= w114 and not w10267;
w10269 <= w118 and not w10268;
w10270 <= w122 and not w10269;
w10271 <= w126 and not w10270;
w10272 <= w130 and not w10271;
w10273 <= w134 and not w10272;
w10274 <= w138 and not w10273;
w10275 <= w142 and not w10274;
w10276 <= w146 and not w10275;
w10277 <= w150 and not w10276;
w10278 <= w154 and not w10277;
w10279 <= w158 and not w10278;
w10280 <= w162 and not w10279;
w10281 <= w166 and not w10280;
w10282 <= w170 and not w10281;
w10283 <= w174 and not w10282;
w10284 <= w178 and not w10283;
w10285 <= w182 and not w10284;
w10286 <= w186 and not w10285;
w10287 <= w190 and not w10286;
w10288 <= w194 and not w10287;
w10289 <= w198 and not w10288;
w10290 <= w202 and not w10289;
w10291 <= w206 and not w10290;
w10292 <= w210 and not w10291;
w10293 <= w214 and not w10292;
w10294 <= w218 and not w10293;
w10295 <= w222 and not w10294;
w10296 <= w226 and not w10295;
w10297 <= w230 and not w10296;
w10298 <= w234 and not w10297;
w10299 <= w238 and not w10298;
w10300 <= w242 and not w10299;
w10301 <= w246 and not w10300;
w10302 <= w250 and not w10301;
w10303 <= w254 and not w10302;
w10304 <= w258 and not w10303;
w10305 <= w262 and not w10304;
w10306 <= w266 and not w10305;
w10307 <= w270 and not w10306;
w10308 <= w274 and not w10307;
w10309 <= w278 and not w10308;
w10310 <= w282 and not w10309;
w10311 <= w286 and not w10310;
w10312 <= req(110) and not w288;
w10313 <= not w10311 and w10312;
w10314 <= w297 and not w632;
w10315 <= w302 and not w10314;
w10316 <= w306 and not w10315;
w10317 <= w310 and not w10316;
w10318 <= w314 and not w10317;
w10319 <= w318 and not w10318;
w10320 <= w322 and not w10319;
w10321 <= w326 and not w10320;
w10322 <= w330 and not w10321;
w10323 <= w334 and not w10322;
w10324 <= w1098 and not w10323;
w10325 <= w1100 and not w10324;
w10326 <= w1364 and not w10325;
w10327 <= w345 and not w10326;
w10328 <= w349 and not w10327;
w10329 <= w353 and not w10328;
w10330 <= w357 and not w10329;
w10331 <= w361 and not w10330;
w10332 <= w365 and not w10331;
w10333 <= w369 and not w10332;
w10334 <= w373 and not w10333;
w10335 <= w377 and not w10334;
w10336 <= w381 and not w10335;
w10337 <= w385 and not w10336;
w10338 <= w389 and not w10337;
w10339 <= w393 and not w10338;
w10340 <= w397 and not w10339;
w10341 <= w401 and not w10340;
w10342 <= w405 and not w10341;
w10343 <= w409 and not w10342;
w10344 <= w413 and not w10343;
w10345 <= w417 and not w10344;
w10346 <= w421 and not w10345;
w10347 <= w425 and not w10346;
w10348 <= w429 and not w10347;
w10349 <= w433 and not w10348;
w10350 <= w437 and not w10349;
w10351 <= w441 and not w10350;
w10352 <= w445 and not w10351;
w10353 <= w449 and not w10352;
w10354 <= w453 and not w10353;
w10355 <= w457 and not w10354;
w10356 <= w461 and not w10355;
w10357 <= w465 and not w10356;
w10358 <= w469 and not w10357;
w10359 <= w473 and not w10358;
w10360 <= w477 and not w10359;
w10361 <= w481 and not w10360;
w10362 <= w485 and not w10361;
w10363 <= w489 and not w10362;
w10364 <= w493 and not w10363;
w10365 <= w497 and not w10364;
w10366 <= w501 and not w10365;
w10367 <= w505 and not w10366;
w10368 <= w509 and not w10367;
w10369 <= w513 and not w10368;
w10370 <= w517 and not w10369;
w10371 <= w521 and not w10370;
w10372 <= w525 and not w10371;
w10373 <= w529 and not w10372;
w10374 <= w533 and not w10373;
w10375 <= w537 and not w10374;
w10376 <= w541 and not w10375;
w10377 <= w545 and not w10376;
w10378 <= w549 and not w10377;
w10379 <= w553 and not w10378;
w10380 <= w557 and not w10379;
w10381 <= w561 and not w10380;
w10382 <= w565 and not w10381;
w10383 <= w569 and not w10382;
w10384 <= w573 and not w10383;
w10385 <= w577 and not w10384;
w10386 <= w581 and not w10385;
w10387 <= w585 and not w10386;
w10388 <= w589 and not w10387;
w10389 <= w593 and not w10388;
w10390 <= w597 and not w10389;
w10391 <= w601 and not w10390;
w10392 <= w605 and not w10391;
w10393 <= w609 and not w10392;
w10394 <= w613 and not w10393;
w10395 <= w617 and not w10394;
w10396 <= w621 and not w10395;
w10397 <= w625 and not w10396;
w10398 <= req(111) and not w627;
w10399 <= not w10397 and w10398;
w10400 <= w636 and not w969;
w10401 <= w641 and not w10400;
w10402 <= w645 and not w10401;
w10403 <= w649 and not w10402;
w10404 <= w653 and not w10403;
w10405 <= w657 and not w10404;
w10406 <= w661 and not w10405;
w10407 <= w665 and not w10406;
w10408 <= w669 and not w10407;
w10409 <= w673 and not w10408;
w10410 <= w1188 and not w10409;
w10411 <= w1190 and not w10410;
w10412 <= w1451 and not w10411;
w10413 <= w682 and not w10412;
w10414 <= w686 and not w10413;
w10415 <= w690 and not w10414;
w10416 <= w694 and not w10415;
w10417 <= w698 and not w10416;
w10418 <= w702 and not w10417;
w10419 <= w706 and not w10418;
w10420 <= w710 and not w10419;
w10421 <= w714 and not w10420;
w10422 <= w718 and not w10421;
w10423 <= w722 and not w10422;
w10424 <= w726 and not w10423;
w10425 <= w730 and not w10424;
w10426 <= w734 and not w10425;
w10427 <= w738 and not w10426;
w10428 <= w742 and not w10427;
w10429 <= w746 and not w10428;
w10430 <= w750 and not w10429;
w10431 <= w754 and not w10430;
w10432 <= w758 and not w10431;
w10433 <= w762 and not w10432;
w10434 <= w766 and not w10433;
w10435 <= w770 and not w10434;
w10436 <= w774 and not w10435;
w10437 <= w778 and not w10436;
w10438 <= w782 and not w10437;
w10439 <= w786 and not w10438;
w10440 <= w790 and not w10439;
w10441 <= w794 and not w10440;
w10442 <= w798 and not w10441;
w10443 <= w802 and not w10442;
w10444 <= w806 and not w10443;
w10445 <= w810 and not w10444;
w10446 <= w814 and not w10445;
w10447 <= w818 and not w10446;
w10448 <= w822 and not w10447;
w10449 <= w826 and not w10448;
w10450 <= w830 and not w10449;
w10451 <= w834 and not w10450;
w10452 <= w838 and not w10451;
w10453 <= w842 and not w10452;
w10454 <= w846 and not w10453;
w10455 <= w850 and not w10454;
w10456 <= w854 and not w10455;
w10457 <= w858 and not w10456;
w10458 <= w862 and not w10457;
w10459 <= w866 and not w10458;
w10460 <= w870 and not w10459;
w10461 <= w874 and not w10460;
w10462 <= w878 and not w10461;
w10463 <= w882 and not w10462;
w10464 <= w886 and not w10463;
w10465 <= w890 and not w10464;
w10466 <= w894 and not w10465;
w10467 <= w898 and not w10466;
w10468 <= w902 and not w10467;
w10469 <= w906 and not w10468;
w10470 <= w910 and not w10469;
w10471 <= w914 and not w10470;
w10472 <= w918 and not w10471;
w10473 <= w922 and not w10472;
w10474 <= w926 and not w10473;
w10475 <= w930 and not w10474;
w10476 <= w934 and not w10475;
w10477 <= w938 and not w10476;
w10478 <= w942 and not w10477;
w10479 <= w946 and not w10478;
w10480 <= w950 and not w10479;
w10481 <= w954 and not w10480;
w10482 <= w958 and not w10481;
w10483 <= w962 and not w10482;
w10484 <= req(112) and not w964;
w10485 <= not w10483 and w10484;
w10486 <= not w301 and w973;
w10487 <= w978 and not w10486;
w10488 <= w982 and not w10487;
w10489 <= w986 and not w10488;
w10490 <= w990 and not w10489;
w10491 <= w994 and not w10490;
w10492 <= w998 and not w10491;
w10493 <= w1002 and not w10492;
w10494 <= w1006 and not w10493;
w10495 <= w1010 and not w10494;
w10496 <= w1277 and not w10495;
w10497 <= w6 and not w10496;
w10498 <= w10 and not w10497;
w10499 <= w14 and not w10498;
w10500 <= w18 and not w10499;
w10501 <= w22 and not w10500;
w10502 <= w26 and not w10501;
w10503 <= w30 and not w10502;
w10504 <= w34 and not w10503;
w10505 <= w38 and not w10504;
w10506 <= w42 and not w10505;
w10507 <= w46 and not w10506;
w10508 <= w50 and not w10507;
w10509 <= w54 and not w10508;
w10510 <= w58 and not w10509;
w10511 <= w62 and not w10510;
w10512 <= w66 and not w10511;
w10513 <= w70 and not w10512;
w10514 <= w74 and not w10513;
w10515 <= w78 and not w10514;
w10516 <= w82 and not w10515;
w10517 <= w86 and not w10516;
w10518 <= w90 and not w10517;
w10519 <= w94 and not w10518;
w10520 <= w98 and not w10519;
w10521 <= w102 and not w10520;
w10522 <= w106 and not w10521;
w10523 <= w110 and not w10522;
w10524 <= w114 and not w10523;
w10525 <= w118 and not w10524;
w10526 <= w122 and not w10525;
w10527 <= w126 and not w10526;
w10528 <= w130 and not w10527;
w10529 <= w134 and not w10528;
w10530 <= w138 and not w10529;
w10531 <= w142 and not w10530;
w10532 <= w146 and not w10531;
w10533 <= w150 and not w10532;
w10534 <= w154 and not w10533;
w10535 <= w158 and not w10534;
w10536 <= w162 and not w10535;
w10537 <= w166 and not w10536;
w10538 <= w170 and not w10537;
w10539 <= w174 and not w10538;
w10540 <= w178 and not w10539;
w10541 <= w182 and not w10540;
w10542 <= w186 and not w10541;
w10543 <= w190 and not w10542;
w10544 <= w194 and not w10543;
w10545 <= w198 and not w10544;
w10546 <= w202 and not w10545;
w10547 <= w206 and not w10546;
w10548 <= w210 and not w10547;
w10549 <= w214 and not w10548;
w10550 <= w218 and not w10549;
w10551 <= w222 and not w10550;
w10552 <= w226 and not w10551;
w10553 <= w230 and not w10552;
w10554 <= w234 and not w10553;
w10555 <= w238 and not w10554;
w10556 <= w242 and not w10555;
w10557 <= w246 and not w10556;
w10558 <= w250 and not w10557;
w10559 <= w254 and not w10558;
w10560 <= w258 and not w10559;
w10561 <= w262 and not w10560;
w10562 <= w266 and not w10561;
w10563 <= w270 and not w10562;
w10564 <= w274 and not w10563;
w10565 <= w278 and not w10564;
w10566 <= w282 and not w10565;
w10567 <= w286 and not w10566;
w10568 <= w290 and not w10567;
w10569 <= w294 and not w10568;
w10570 <= req(113) and not w296;
w10571 <= not w10569 and w10570;
w10572 <= w305 and not w640;
w10573 <= w310 and not w10572;
w10574 <= w314 and not w10573;
w10575 <= w318 and not w10574;
w10576 <= w322 and not w10575;
w10577 <= w326 and not w10576;
w10578 <= w330 and not w10577;
w10579 <= w334 and not w10578;
w10580 <= w1098 and not w10579;
w10581 <= w1100 and not w10580;
w10582 <= w1364 and not w10581;
w10583 <= w345 and not w10582;
w10584 <= w349 and not w10583;
w10585 <= w353 and not w10584;
w10586 <= w357 and not w10585;
w10587 <= w361 and not w10586;
w10588 <= w365 and not w10587;
w10589 <= w369 and not w10588;
w10590 <= w373 and not w10589;
w10591 <= w377 and not w10590;
w10592 <= w381 and not w10591;
w10593 <= w385 and not w10592;
w10594 <= w389 and not w10593;
w10595 <= w393 and not w10594;
w10596 <= w397 and not w10595;
w10597 <= w401 and not w10596;
w10598 <= w405 and not w10597;
w10599 <= w409 and not w10598;
w10600 <= w413 and not w10599;
w10601 <= w417 and not w10600;
w10602 <= w421 and not w10601;
w10603 <= w425 and not w10602;
w10604 <= w429 and not w10603;
w10605 <= w433 and not w10604;
w10606 <= w437 and not w10605;
w10607 <= w441 and not w10606;
w10608 <= w445 and not w10607;
w10609 <= w449 and not w10608;
w10610 <= w453 and not w10609;
w10611 <= w457 and not w10610;
w10612 <= w461 and not w10611;
w10613 <= w465 and not w10612;
w10614 <= w469 and not w10613;
w10615 <= w473 and not w10614;
w10616 <= w477 and not w10615;
w10617 <= w481 and not w10616;
w10618 <= w485 and not w10617;
w10619 <= w489 and not w10618;
w10620 <= w493 and not w10619;
w10621 <= w497 and not w10620;
w10622 <= w501 and not w10621;
w10623 <= w505 and not w10622;
w10624 <= w509 and not w10623;
w10625 <= w513 and not w10624;
w10626 <= w517 and not w10625;
w10627 <= w521 and not w10626;
w10628 <= w525 and not w10627;
w10629 <= w529 and not w10628;
w10630 <= w533 and not w10629;
w10631 <= w537 and not w10630;
w10632 <= w541 and not w10631;
w10633 <= w545 and not w10632;
w10634 <= w549 and not w10633;
w10635 <= w553 and not w10634;
w10636 <= w557 and not w10635;
w10637 <= w561 and not w10636;
w10638 <= w565 and not w10637;
w10639 <= w569 and not w10638;
w10640 <= w573 and not w10639;
w10641 <= w577 and not w10640;
w10642 <= w581 and not w10641;
w10643 <= w585 and not w10642;
w10644 <= w589 and not w10643;
w10645 <= w593 and not w10644;
w10646 <= w597 and not w10645;
w10647 <= w601 and not w10646;
w10648 <= w605 and not w10647;
w10649 <= w609 and not w10648;
w10650 <= w613 and not w10649;
w10651 <= w617 and not w10650;
w10652 <= w621 and not w10651;
w10653 <= w625 and not w10652;
w10654 <= w629 and not w10653;
w10655 <= w633 and not w10654;
w10656 <= req(114) and not w635;
w10657 <= not w10655 and w10656;
w10658 <= w644 and not w977;
w10659 <= w649 and not w10658;
w10660 <= w653 and not w10659;
w10661 <= w657 and not w10660;
w10662 <= w661 and not w10661;
w10663 <= w665 and not w10662;
w10664 <= w669 and not w10663;
w10665 <= w673 and not w10664;
w10666 <= w1188 and not w10665;
w10667 <= w1190 and not w10666;
w10668 <= w1451 and not w10667;
w10669 <= w682 and not w10668;
w10670 <= w686 and not w10669;
w10671 <= w690 and not w10670;
w10672 <= w694 and not w10671;
w10673 <= w698 and not w10672;
w10674 <= w702 and not w10673;
w10675 <= w706 and not w10674;
w10676 <= w710 and not w10675;
w10677 <= w714 and not w10676;
w10678 <= w718 and not w10677;
w10679 <= w722 and not w10678;
w10680 <= w726 and not w10679;
w10681 <= w730 and not w10680;
w10682 <= w734 and not w10681;
w10683 <= w738 and not w10682;
w10684 <= w742 and not w10683;
w10685 <= w746 and not w10684;
w10686 <= w750 and not w10685;
w10687 <= w754 and not w10686;
w10688 <= w758 and not w10687;
w10689 <= w762 and not w10688;
w10690 <= w766 and not w10689;
w10691 <= w770 and not w10690;
w10692 <= w774 and not w10691;
w10693 <= w778 and not w10692;
w10694 <= w782 and not w10693;
w10695 <= w786 and not w10694;
w10696 <= w790 and not w10695;
w10697 <= w794 and not w10696;
w10698 <= w798 and not w10697;
w10699 <= w802 and not w10698;
w10700 <= w806 and not w10699;
w10701 <= w810 and not w10700;
w10702 <= w814 and not w10701;
w10703 <= w818 and not w10702;
w10704 <= w822 and not w10703;
w10705 <= w826 and not w10704;
w10706 <= w830 and not w10705;
w10707 <= w834 and not w10706;
w10708 <= w838 and not w10707;
w10709 <= w842 and not w10708;
w10710 <= w846 and not w10709;
w10711 <= w850 and not w10710;
w10712 <= w854 and not w10711;
w10713 <= w858 and not w10712;
w10714 <= w862 and not w10713;
w10715 <= w866 and not w10714;
w10716 <= w870 and not w10715;
w10717 <= w874 and not w10716;
w10718 <= w878 and not w10717;
w10719 <= w882 and not w10718;
w10720 <= w886 and not w10719;
w10721 <= w890 and not w10720;
w10722 <= w894 and not w10721;
w10723 <= w898 and not w10722;
w10724 <= w902 and not w10723;
w10725 <= w906 and not w10724;
w10726 <= w910 and not w10725;
w10727 <= w914 and not w10726;
w10728 <= w918 and not w10727;
w10729 <= w922 and not w10728;
w10730 <= w926 and not w10729;
w10731 <= w930 and not w10730;
w10732 <= w934 and not w10731;
w10733 <= w938 and not w10732;
w10734 <= w942 and not w10733;
w10735 <= w946 and not w10734;
w10736 <= w950 and not w10735;
w10737 <= w954 and not w10736;
w10738 <= w958 and not w10737;
w10739 <= w962 and not w10738;
w10740 <= w966 and not w10739;
w10741 <= w970 and not w10740;
w10742 <= req(115) and not w972;
w10743 <= not w10741 and w10742;
w10744 <= not w309 and w981;
w10745 <= w986 and not w10744;
w10746 <= w990 and not w10745;
w10747 <= w994 and not w10746;
w10748 <= w998 and not w10747;
w10749 <= w1002 and not w10748;
w10750 <= w1006 and not w10749;
w10751 <= w1010 and not w10750;
w10752 <= w1277 and not w10751;
w10753 <= w6 and not w10752;
w10754 <= w10 and not w10753;
w10755 <= w14 and not w10754;
w10756 <= w18 and not w10755;
w10757 <= w22 and not w10756;
w10758 <= w26 and not w10757;
w10759 <= w30 and not w10758;
w10760 <= w34 and not w10759;
w10761 <= w38 and not w10760;
w10762 <= w42 and not w10761;
w10763 <= w46 and not w10762;
w10764 <= w50 and not w10763;
w10765 <= w54 and not w10764;
w10766 <= w58 and not w10765;
w10767 <= w62 and not w10766;
w10768 <= w66 and not w10767;
w10769 <= w70 and not w10768;
w10770 <= w74 and not w10769;
w10771 <= w78 and not w10770;
w10772 <= w82 and not w10771;
w10773 <= w86 and not w10772;
w10774 <= w90 and not w10773;
w10775 <= w94 and not w10774;
w10776 <= w98 and not w10775;
w10777 <= w102 and not w10776;
w10778 <= w106 and not w10777;
w10779 <= w110 and not w10778;
w10780 <= w114 and not w10779;
w10781 <= w118 and not w10780;
w10782 <= w122 and not w10781;
w10783 <= w126 and not w10782;
w10784 <= w130 and not w10783;
w10785 <= w134 and not w10784;
w10786 <= w138 and not w10785;
w10787 <= w142 and not w10786;
w10788 <= w146 and not w10787;
w10789 <= w150 and not w10788;
w10790 <= w154 and not w10789;
w10791 <= w158 and not w10790;
w10792 <= w162 and not w10791;
w10793 <= w166 and not w10792;
w10794 <= w170 and not w10793;
w10795 <= w174 and not w10794;
w10796 <= w178 and not w10795;
w10797 <= w182 and not w10796;
w10798 <= w186 and not w10797;
w10799 <= w190 and not w10798;
w10800 <= w194 and not w10799;
w10801 <= w198 and not w10800;
w10802 <= w202 and not w10801;
w10803 <= w206 and not w10802;
w10804 <= w210 and not w10803;
w10805 <= w214 and not w10804;
w10806 <= w218 and not w10805;
w10807 <= w222 and not w10806;
w10808 <= w226 and not w10807;
w10809 <= w230 and not w10808;
w10810 <= w234 and not w10809;
w10811 <= w238 and not w10810;
w10812 <= w242 and not w10811;
w10813 <= w246 and not w10812;
w10814 <= w250 and not w10813;
w10815 <= w254 and not w10814;
w10816 <= w258 and not w10815;
w10817 <= w262 and not w10816;
w10818 <= w266 and not w10817;
w10819 <= w270 and not w10818;
w10820 <= w274 and not w10819;
w10821 <= w278 and not w10820;
w10822 <= w282 and not w10821;
w10823 <= w286 and not w10822;
w10824 <= w290 and not w10823;
w10825 <= w294 and not w10824;
w10826 <= w298 and not w10825;
w10827 <= w302 and not w10826;
w10828 <= req(116) and not w304;
w10829 <= not w10827 and w10828;
w10830 <= w313 and not w648;
w10831 <= w318 and not w10830;
w10832 <= w322 and not w10831;
w10833 <= w326 and not w10832;
w10834 <= w330 and not w10833;
w10835 <= w334 and not w10834;
w10836 <= w1098 and not w10835;
w10837 <= w1100 and not w10836;
w10838 <= w1364 and not w10837;
w10839 <= w345 and not w10838;
w10840 <= w349 and not w10839;
w10841 <= w353 and not w10840;
w10842 <= w357 and not w10841;
w10843 <= w361 and not w10842;
w10844 <= w365 and not w10843;
w10845 <= w369 and not w10844;
w10846 <= w373 and not w10845;
w10847 <= w377 and not w10846;
w10848 <= w381 and not w10847;
w10849 <= w385 and not w10848;
w10850 <= w389 and not w10849;
w10851 <= w393 and not w10850;
w10852 <= w397 and not w10851;
w10853 <= w401 and not w10852;
w10854 <= w405 and not w10853;
w10855 <= w409 and not w10854;
w10856 <= w413 and not w10855;
w10857 <= w417 and not w10856;
w10858 <= w421 and not w10857;
w10859 <= w425 and not w10858;
w10860 <= w429 and not w10859;
w10861 <= w433 and not w10860;
w10862 <= w437 and not w10861;
w10863 <= w441 and not w10862;
w10864 <= w445 and not w10863;
w10865 <= w449 and not w10864;
w10866 <= w453 and not w10865;
w10867 <= w457 and not w10866;
w10868 <= w461 and not w10867;
w10869 <= w465 and not w10868;
w10870 <= w469 and not w10869;
w10871 <= w473 and not w10870;
w10872 <= w477 and not w10871;
w10873 <= w481 and not w10872;
w10874 <= w485 and not w10873;
w10875 <= w489 and not w10874;
w10876 <= w493 and not w10875;
w10877 <= w497 and not w10876;
w10878 <= w501 and not w10877;
w10879 <= w505 and not w10878;
w10880 <= w509 and not w10879;
w10881 <= w513 and not w10880;
w10882 <= w517 and not w10881;
w10883 <= w521 and not w10882;
w10884 <= w525 and not w10883;
w10885 <= w529 and not w10884;
w10886 <= w533 and not w10885;
w10887 <= w537 and not w10886;
w10888 <= w541 and not w10887;
w10889 <= w545 and not w10888;
w10890 <= w549 and not w10889;
w10891 <= w553 and not w10890;
w10892 <= w557 and not w10891;
w10893 <= w561 and not w10892;
w10894 <= w565 and not w10893;
w10895 <= w569 and not w10894;
w10896 <= w573 and not w10895;
w10897 <= w577 and not w10896;
w10898 <= w581 and not w10897;
w10899 <= w585 and not w10898;
w10900 <= w589 and not w10899;
w10901 <= w593 and not w10900;
w10902 <= w597 and not w10901;
w10903 <= w601 and not w10902;
w10904 <= w605 and not w10903;
w10905 <= w609 and not w10904;
w10906 <= w613 and not w10905;
w10907 <= w617 and not w10906;
w10908 <= w621 and not w10907;
w10909 <= w625 and not w10908;
w10910 <= w629 and not w10909;
w10911 <= w633 and not w10910;
w10912 <= w637 and not w10911;
w10913 <= w641 and not w10912;
w10914 <= req(117) and not w643;
w10915 <= not w10913 and w10914;
w10916 <= w652 and not w985;
w10917 <= w657 and not w10916;
w10918 <= w661 and not w10917;
w10919 <= w665 and not w10918;
w10920 <= w669 and not w10919;
w10921 <= w673 and not w10920;
w10922 <= w1188 and not w10921;
w10923 <= w1190 and not w10922;
w10924 <= w1451 and not w10923;
w10925 <= w682 and not w10924;
w10926 <= w686 and not w10925;
w10927 <= w690 and not w10926;
w10928 <= w694 and not w10927;
w10929 <= w698 and not w10928;
w10930 <= w702 and not w10929;
w10931 <= w706 and not w10930;
w10932 <= w710 and not w10931;
w10933 <= w714 and not w10932;
w10934 <= w718 and not w10933;
w10935 <= w722 and not w10934;
w10936 <= w726 and not w10935;
w10937 <= w730 and not w10936;
w10938 <= w734 and not w10937;
w10939 <= w738 and not w10938;
w10940 <= w742 and not w10939;
w10941 <= w746 and not w10940;
w10942 <= w750 and not w10941;
w10943 <= w754 and not w10942;
w10944 <= w758 and not w10943;
w10945 <= w762 and not w10944;
w10946 <= w766 and not w10945;
w10947 <= w770 and not w10946;
w10948 <= w774 and not w10947;
w10949 <= w778 and not w10948;
w10950 <= w782 and not w10949;
w10951 <= w786 and not w10950;
w10952 <= w790 and not w10951;
w10953 <= w794 and not w10952;
w10954 <= w798 and not w10953;
w10955 <= w802 and not w10954;
w10956 <= w806 and not w10955;
w10957 <= w810 and not w10956;
w10958 <= w814 and not w10957;
w10959 <= w818 and not w10958;
w10960 <= w822 and not w10959;
w10961 <= w826 and not w10960;
w10962 <= w830 and not w10961;
w10963 <= w834 and not w10962;
w10964 <= w838 and not w10963;
w10965 <= w842 and not w10964;
w10966 <= w846 and not w10965;
w10967 <= w850 and not w10966;
w10968 <= w854 and not w10967;
w10969 <= w858 and not w10968;
w10970 <= w862 and not w10969;
w10971 <= w866 and not w10970;
w10972 <= w870 and not w10971;
w10973 <= w874 and not w10972;
w10974 <= w878 and not w10973;
w10975 <= w882 and not w10974;
w10976 <= w886 and not w10975;
w10977 <= w890 and not w10976;
w10978 <= w894 and not w10977;
w10979 <= w898 and not w10978;
w10980 <= w902 and not w10979;
w10981 <= w906 and not w10980;
w10982 <= w910 and not w10981;
w10983 <= w914 and not w10982;
w10984 <= w918 and not w10983;
w10985 <= w922 and not w10984;
w10986 <= w926 and not w10985;
w10987 <= w930 and not w10986;
w10988 <= w934 and not w10987;
w10989 <= w938 and not w10988;
w10990 <= w942 and not w10989;
w10991 <= w946 and not w10990;
w10992 <= w950 and not w10991;
w10993 <= w954 and not w10992;
w10994 <= w958 and not w10993;
w10995 <= w962 and not w10994;
w10996 <= w966 and not w10995;
w10997 <= w970 and not w10996;
w10998 <= w974 and not w10997;
w10999 <= w978 and not w10998;
w11000 <= req(118) and not w980;
w11001 <= not w10999 and w11000;
w11002 <= not w317 and w989;
w11003 <= w994 and not w11002;
w11004 <= w998 and not w11003;
w11005 <= w1002 and not w11004;
w11006 <= w1006 and not w11005;
w11007 <= w1010 and not w11006;
w11008 <= w1277 and not w11007;
w11009 <= w6 and not w11008;
w11010 <= w10 and not w11009;
w11011 <= w14 and not w11010;
w11012 <= w18 and not w11011;
w11013 <= w22 and not w11012;
w11014 <= w26 and not w11013;
w11015 <= w30 and not w11014;
w11016 <= w34 and not w11015;
w11017 <= w38 and not w11016;
w11018 <= w42 and not w11017;
w11019 <= w46 and not w11018;
w11020 <= w50 and not w11019;
w11021 <= w54 and not w11020;
w11022 <= w58 and not w11021;
w11023 <= w62 and not w11022;
w11024 <= w66 and not w11023;
w11025 <= w70 and not w11024;
w11026 <= w74 and not w11025;
w11027 <= w78 and not w11026;
w11028 <= w82 and not w11027;
w11029 <= w86 and not w11028;
w11030 <= w90 and not w11029;
w11031 <= w94 and not w11030;
w11032 <= w98 and not w11031;
w11033 <= w102 and not w11032;
w11034 <= w106 and not w11033;
w11035 <= w110 and not w11034;
w11036 <= w114 and not w11035;
w11037 <= w118 and not w11036;
w11038 <= w122 and not w11037;
w11039 <= w126 and not w11038;
w11040 <= w130 and not w11039;
w11041 <= w134 and not w11040;
w11042 <= w138 and not w11041;
w11043 <= w142 and not w11042;
w11044 <= w146 and not w11043;
w11045 <= w150 and not w11044;
w11046 <= w154 and not w11045;
w11047 <= w158 and not w11046;
w11048 <= w162 and not w11047;
w11049 <= w166 and not w11048;
w11050 <= w170 and not w11049;
w11051 <= w174 and not w11050;
w11052 <= w178 and not w11051;
w11053 <= w182 and not w11052;
w11054 <= w186 and not w11053;
w11055 <= w190 and not w11054;
w11056 <= w194 and not w11055;
w11057 <= w198 and not w11056;
w11058 <= w202 and not w11057;
w11059 <= w206 and not w11058;
w11060 <= w210 and not w11059;
w11061 <= w214 and not w11060;
w11062 <= w218 and not w11061;
w11063 <= w222 and not w11062;
w11064 <= w226 and not w11063;
w11065 <= w230 and not w11064;
w11066 <= w234 and not w11065;
w11067 <= w238 and not w11066;
w11068 <= w242 and not w11067;
w11069 <= w246 and not w11068;
w11070 <= w250 and not w11069;
w11071 <= w254 and not w11070;
w11072 <= w258 and not w11071;
w11073 <= w262 and not w11072;
w11074 <= w266 and not w11073;
w11075 <= w270 and not w11074;
w11076 <= w274 and not w11075;
w11077 <= w278 and not w11076;
w11078 <= w282 and not w11077;
w11079 <= w286 and not w11078;
w11080 <= w290 and not w11079;
w11081 <= w294 and not w11080;
w11082 <= w298 and not w11081;
w11083 <= w302 and not w11082;
w11084 <= w306 and not w11083;
w11085 <= w310 and not w11084;
w11086 <= req(119) and not w312;
w11087 <= not w11085 and w11086;
w11088 <= w321 and not w656;
w11089 <= w326 and not w11088;
w11090 <= w330 and not w11089;
w11091 <= w334 and not w11090;
w11092 <= w1098 and not w11091;
w11093 <= w1100 and not w11092;
w11094 <= w1364 and not w11093;
w11095 <= w345 and not w11094;
w11096 <= w349 and not w11095;
w11097 <= w353 and not w11096;
w11098 <= w357 and not w11097;
w11099 <= w361 and not w11098;
w11100 <= w365 and not w11099;
w11101 <= w369 and not w11100;
w11102 <= w373 and not w11101;
w11103 <= w377 and not w11102;
w11104 <= w381 and not w11103;
w11105 <= w385 and not w11104;
w11106 <= w389 and not w11105;
w11107 <= w393 and not w11106;
w11108 <= w397 and not w11107;
w11109 <= w401 and not w11108;
w11110 <= w405 and not w11109;
w11111 <= w409 and not w11110;
w11112 <= w413 and not w11111;
w11113 <= w417 and not w11112;
w11114 <= w421 and not w11113;
w11115 <= w425 and not w11114;
w11116 <= w429 and not w11115;
w11117 <= w433 and not w11116;
w11118 <= w437 and not w11117;
w11119 <= w441 and not w11118;
w11120 <= w445 and not w11119;
w11121 <= w449 and not w11120;
w11122 <= w453 and not w11121;
w11123 <= w457 and not w11122;
w11124 <= w461 and not w11123;
w11125 <= w465 and not w11124;
w11126 <= w469 and not w11125;
w11127 <= w473 and not w11126;
w11128 <= w477 and not w11127;
w11129 <= w481 and not w11128;
w11130 <= w485 and not w11129;
w11131 <= w489 and not w11130;
w11132 <= w493 and not w11131;
w11133 <= w497 and not w11132;
w11134 <= w501 and not w11133;
w11135 <= w505 and not w11134;
w11136 <= w509 and not w11135;
w11137 <= w513 and not w11136;
w11138 <= w517 and not w11137;
w11139 <= w521 and not w11138;
w11140 <= w525 and not w11139;
w11141 <= w529 and not w11140;
w11142 <= w533 and not w11141;
w11143 <= w537 and not w11142;
w11144 <= w541 and not w11143;
w11145 <= w545 and not w11144;
w11146 <= w549 and not w11145;
w11147 <= w553 and not w11146;
w11148 <= w557 and not w11147;
w11149 <= w561 and not w11148;
w11150 <= w565 and not w11149;
w11151 <= w569 and not w11150;
w11152 <= w573 and not w11151;
w11153 <= w577 and not w11152;
w11154 <= w581 and not w11153;
w11155 <= w585 and not w11154;
w11156 <= w589 and not w11155;
w11157 <= w593 and not w11156;
w11158 <= w597 and not w11157;
w11159 <= w601 and not w11158;
w11160 <= w605 and not w11159;
w11161 <= w609 and not w11160;
w11162 <= w613 and not w11161;
w11163 <= w617 and not w11162;
w11164 <= w621 and not w11163;
w11165 <= w625 and not w11164;
w11166 <= w629 and not w11165;
w11167 <= w633 and not w11166;
w11168 <= w637 and not w11167;
w11169 <= w641 and not w11168;
w11170 <= w645 and not w11169;
w11171 <= w649 and not w11170;
w11172 <= req(120) and not w651;
w11173 <= not w11171 and w11172;
w11174 <= w660 and not w993;
w11175 <= w665 and not w11174;
w11176 <= w669 and not w11175;
w11177 <= w673 and not w11176;
w11178 <= w1188 and not w11177;
w11179 <= w1190 and not w11178;
w11180 <= w1451 and not w11179;
w11181 <= w682 and not w11180;
w11182 <= w686 and not w11181;
w11183 <= w690 and not w11182;
w11184 <= w694 and not w11183;
w11185 <= w698 and not w11184;
w11186 <= w702 and not w11185;
w11187 <= w706 and not w11186;
w11188 <= w710 and not w11187;
w11189 <= w714 and not w11188;
w11190 <= w718 and not w11189;
w11191 <= w722 and not w11190;
w11192 <= w726 and not w11191;
w11193 <= w730 and not w11192;
w11194 <= w734 and not w11193;
w11195 <= w738 and not w11194;
w11196 <= w742 and not w11195;
w11197 <= w746 and not w11196;
w11198 <= w750 and not w11197;
w11199 <= w754 and not w11198;
w11200 <= w758 and not w11199;
w11201 <= w762 and not w11200;
w11202 <= w766 and not w11201;
w11203 <= w770 and not w11202;
w11204 <= w774 and not w11203;
w11205 <= w778 and not w11204;
w11206 <= w782 and not w11205;
w11207 <= w786 and not w11206;
w11208 <= w790 and not w11207;
w11209 <= w794 and not w11208;
w11210 <= w798 and not w11209;
w11211 <= w802 and not w11210;
w11212 <= w806 and not w11211;
w11213 <= w810 and not w11212;
w11214 <= w814 and not w11213;
w11215 <= w818 and not w11214;
w11216 <= w822 and not w11215;
w11217 <= w826 and not w11216;
w11218 <= w830 and not w11217;
w11219 <= w834 and not w11218;
w11220 <= w838 and not w11219;
w11221 <= w842 and not w11220;
w11222 <= w846 and not w11221;
w11223 <= w850 and not w11222;
w11224 <= w854 and not w11223;
w11225 <= w858 and not w11224;
w11226 <= w862 and not w11225;
w11227 <= w866 and not w11226;
w11228 <= w870 and not w11227;
w11229 <= w874 and not w11228;
w11230 <= w878 and not w11229;
w11231 <= w882 and not w11230;
w11232 <= w886 and not w11231;
w11233 <= w890 and not w11232;
w11234 <= w894 and not w11233;
w11235 <= w898 and not w11234;
w11236 <= w902 and not w11235;
w11237 <= w906 and not w11236;
w11238 <= w910 and not w11237;
w11239 <= w914 and not w11238;
w11240 <= w918 and not w11239;
w11241 <= w922 and not w11240;
w11242 <= w926 and not w11241;
w11243 <= w930 and not w11242;
w11244 <= w934 and not w11243;
w11245 <= w938 and not w11244;
w11246 <= w942 and not w11245;
w11247 <= w946 and not w11246;
w11248 <= w950 and not w11247;
w11249 <= w954 and not w11248;
w11250 <= w958 and not w11249;
w11251 <= w962 and not w11250;
w11252 <= w966 and not w11251;
w11253 <= w970 and not w11252;
w11254 <= w974 and not w11253;
w11255 <= w978 and not w11254;
w11256 <= w982 and not w11255;
w11257 <= w986 and not w11256;
w11258 <= req(121) and not w988;
w11259 <= not w11257 and w11258;
w11260 <= not w325 and w997;
w11261 <= w1002 and not w11260;
w11262 <= w1006 and not w11261;
w11263 <= w1010 and not w11262;
w11264 <= w1277 and not w11263;
w11265 <= w6 and not w11264;
w11266 <= w10 and not w11265;
w11267 <= w14 and not w11266;
w11268 <= w18 and not w11267;
w11269 <= w22 and not w11268;
w11270 <= w26 and not w11269;
w11271 <= w30 and not w11270;
w11272 <= w34 and not w11271;
w11273 <= w38 and not w11272;
w11274 <= w42 and not w11273;
w11275 <= w46 and not w11274;
w11276 <= w50 and not w11275;
w11277 <= w54 and not w11276;
w11278 <= w58 and not w11277;
w11279 <= w62 and not w11278;
w11280 <= w66 and not w11279;
w11281 <= w70 and not w11280;
w11282 <= w74 and not w11281;
w11283 <= w78 and not w11282;
w11284 <= w82 and not w11283;
w11285 <= w86 and not w11284;
w11286 <= w90 and not w11285;
w11287 <= w94 and not w11286;
w11288 <= w98 and not w11287;
w11289 <= w102 and not w11288;
w11290 <= w106 and not w11289;
w11291 <= w110 and not w11290;
w11292 <= w114 and not w11291;
w11293 <= w118 and not w11292;
w11294 <= w122 and not w11293;
w11295 <= w126 and not w11294;
w11296 <= w130 and not w11295;
w11297 <= w134 and not w11296;
w11298 <= w138 and not w11297;
w11299 <= w142 and not w11298;
w11300 <= w146 and not w11299;
w11301 <= w150 and not w11300;
w11302 <= w154 and not w11301;
w11303 <= w158 and not w11302;
w11304 <= w162 and not w11303;
w11305 <= w166 and not w11304;
w11306 <= w170 and not w11305;
w11307 <= w174 and not w11306;
w11308 <= w178 and not w11307;
w11309 <= w182 and not w11308;
w11310 <= w186 and not w11309;
w11311 <= w190 and not w11310;
w11312 <= w194 and not w11311;
w11313 <= w198 and not w11312;
w11314 <= w202 and not w11313;
w11315 <= w206 and not w11314;
w11316 <= w210 and not w11315;
w11317 <= w214 and not w11316;
w11318 <= w218 and not w11317;
w11319 <= w222 and not w11318;
w11320 <= w226 and not w11319;
w11321 <= w230 and not w11320;
w11322 <= w234 and not w11321;
w11323 <= w238 and not w11322;
w11324 <= w242 and not w11323;
w11325 <= w246 and not w11324;
w11326 <= w250 and not w11325;
w11327 <= w254 and not w11326;
w11328 <= w258 and not w11327;
w11329 <= w262 and not w11328;
w11330 <= w266 and not w11329;
w11331 <= w270 and not w11330;
w11332 <= w274 and not w11331;
w11333 <= w278 and not w11332;
w11334 <= w282 and not w11333;
w11335 <= w286 and not w11334;
w11336 <= w290 and not w11335;
w11337 <= w294 and not w11336;
w11338 <= w298 and not w11337;
w11339 <= w302 and not w11338;
w11340 <= w306 and not w11339;
w11341 <= w310 and not w11340;
w11342 <= w314 and not w11341;
w11343 <= w318 and not w11342;
w11344 <= req(122) and not w320;
w11345 <= not w11343 and w11344;
w11346 <= w329 and not w664;
w11347 <= w334 and not w11346;
w11348 <= w1098 and not w11347;
w11349 <= w1100 and not w11348;
w11350 <= w1364 and not w11349;
w11351 <= w345 and not w11350;
w11352 <= w349 and not w11351;
w11353 <= w353 and not w11352;
w11354 <= w357 and not w11353;
w11355 <= w361 and not w11354;
w11356 <= w365 and not w11355;
w11357 <= w369 and not w11356;
w11358 <= w373 and not w11357;
w11359 <= w377 and not w11358;
w11360 <= w381 and not w11359;
w11361 <= w385 and not w11360;
w11362 <= w389 and not w11361;
w11363 <= w393 and not w11362;
w11364 <= w397 and not w11363;
w11365 <= w401 and not w11364;
w11366 <= w405 and not w11365;
w11367 <= w409 and not w11366;
w11368 <= w413 and not w11367;
w11369 <= w417 and not w11368;
w11370 <= w421 and not w11369;
w11371 <= w425 and not w11370;
w11372 <= w429 and not w11371;
w11373 <= w433 and not w11372;
w11374 <= w437 and not w11373;
w11375 <= w441 and not w11374;
w11376 <= w445 and not w11375;
w11377 <= w449 and not w11376;
w11378 <= w453 and not w11377;
w11379 <= w457 and not w11378;
w11380 <= w461 and not w11379;
w11381 <= w465 and not w11380;
w11382 <= w469 and not w11381;
w11383 <= w473 and not w11382;
w11384 <= w477 and not w11383;
w11385 <= w481 and not w11384;
w11386 <= w485 and not w11385;
w11387 <= w489 and not w11386;
w11388 <= w493 and not w11387;
w11389 <= w497 and not w11388;
w11390 <= w501 and not w11389;
w11391 <= w505 and not w11390;
w11392 <= w509 and not w11391;
w11393 <= w513 and not w11392;
w11394 <= w517 and not w11393;
w11395 <= w521 and not w11394;
w11396 <= w525 and not w11395;
w11397 <= w529 and not w11396;
w11398 <= w533 and not w11397;
w11399 <= w537 and not w11398;
w11400 <= w541 and not w11399;
w11401 <= w545 and not w11400;
w11402 <= w549 and not w11401;
w11403 <= w553 and not w11402;
w11404 <= w557 and not w11403;
w11405 <= w561 and not w11404;
w11406 <= w565 and not w11405;
w11407 <= w569 and not w11406;
w11408 <= w573 and not w11407;
w11409 <= w577 and not w11408;
w11410 <= w581 and not w11409;
w11411 <= w585 and not w11410;
w11412 <= w589 and not w11411;
w11413 <= w593 and not w11412;
w11414 <= w597 and not w11413;
w11415 <= w601 and not w11414;
w11416 <= w605 and not w11415;
w11417 <= w609 and not w11416;
w11418 <= w613 and not w11417;
w11419 <= w617 and not w11418;
w11420 <= w621 and not w11419;
w11421 <= w625 and not w11420;
w11422 <= w629 and not w11421;
w11423 <= w633 and not w11422;
w11424 <= w637 and not w11423;
w11425 <= w641 and not w11424;
w11426 <= w645 and not w11425;
w11427 <= w649 and not w11426;
w11428 <= w653 and not w11427;
w11429 <= w657 and not w11428;
w11430 <= req(123) and not w659;
w11431 <= not w11429 and w11430;
w11432 <= w668 and not w1001;
w11433 <= w673 and not w11432;
w11434 <= w1188 and not w11433;
w11435 <= w1190 and not w11434;
w11436 <= w1451 and not w11435;
w11437 <= w682 and not w11436;
w11438 <= w686 and not w11437;
w11439 <= w690 and not w11438;
w11440 <= w694 and not w11439;
w11441 <= w698 and not w11440;
w11442 <= w702 and not w11441;
w11443 <= w706 and not w11442;
w11444 <= w710 and not w11443;
w11445 <= w714 and not w11444;
w11446 <= w718 and not w11445;
w11447 <= w722 and not w11446;
w11448 <= w726 and not w11447;
w11449 <= w730 and not w11448;
w11450 <= w734 and not w11449;
w11451 <= w738 and not w11450;
w11452 <= w742 and not w11451;
w11453 <= w746 and not w11452;
w11454 <= w750 and not w11453;
w11455 <= w754 and not w11454;
w11456 <= w758 and not w11455;
w11457 <= w762 and not w11456;
w11458 <= w766 and not w11457;
w11459 <= w770 and not w11458;
w11460 <= w774 and not w11459;
w11461 <= w778 and not w11460;
w11462 <= w782 and not w11461;
w11463 <= w786 and not w11462;
w11464 <= w790 and not w11463;
w11465 <= w794 and not w11464;
w11466 <= w798 and not w11465;
w11467 <= w802 and not w11466;
w11468 <= w806 and not w11467;
w11469 <= w810 and not w11468;
w11470 <= w814 and not w11469;
w11471 <= w818 and not w11470;
w11472 <= w822 and not w11471;
w11473 <= w826 and not w11472;
w11474 <= w830 and not w11473;
w11475 <= w834 and not w11474;
w11476 <= w838 and not w11475;
w11477 <= w842 and not w11476;
w11478 <= w846 and not w11477;
w11479 <= w850 and not w11478;
w11480 <= w854 and not w11479;
w11481 <= w858 and not w11480;
w11482 <= w862 and not w11481;
w11483 <= w866 and not w11482;
w11484 <= w870 and not w11483;
w11485 <= w874 and not w11484;
w11486 <= w878 and not w11485;
w11487 <= w882 and not w11486;
w11488 <= w886 and not w11487;
w11489 <= w890 and not w11488;
w11490 <= w894 and not w11489;
w11491 <= w898 and not w11490;
w11492 <= w902 and not w11491;
w11493 <= w906 and not w11492;
w11494 <= w910 and not w11493;
w11495 <= w914 and not w11494;
w11496 <= w918 and not w11495;
w11497 <= w922 and not w11496;
w11498 <= w926 and not w11497;
w11499 <= w930 and not w11498;
w11500 <= w934 and not w11499;
w11501 <= w938 and not w11500;
w11502 <= w942 and not w11501;
w11503 <= w946 and not w11502;
w11504 <= w950 and not w11503;
w11505 <= w954 and not w11504;
w11506 <= w958 and not w11505;
w11507 <= w962 and not w11506;
w11508 <= w966 and not w11507;
w11509 <= w970 and not w11508;
w11510 <= w974 and not w11509;
w11511 <= w978 and not w11510;
w11512 <= w982 and not w11511;
w11513 <= w986 and not w11512;
w11514 <= w990 and not w11513;
w11515 <= w994 and not w11514;
w11516 <= req(124) and not w996;
w11517 <= not w11515 and w11516;
w11518 <= not w333 and w1005;
w11519 <= w1010 and not w11518;
w11520 <= w1277 and not w11519;
w11521 <= w6 and not w11520;
w11522 <= w10 and not w11521;
w11523 <= w14 and not w11522;
w11524 <= w18 and not w11523;
w11525 <= w22 and not w11524;
w11526 <= w26 and not w11525;
w11527 <= w30 and not w11526;
w11528 <= w34 and not w11527;
w11529 <= w38 and not w11528;
w11530 <= w42 and not w11529;
w11531 <= w46 and not w11530;
w11532 <= w50 and not w11531;
w11533 <= w54 and not w11532;
w11534 <= w58 and not w11533;
w11535 <= w62 and not w11534;
w11536 <= w66 and not w11535;
w11537 <= w70 and not w11536;
w11538 <= w74 and not w11537;
w11539 <= w78 and not w11538;
w11540 <= w82 and not w11539;
w11541 <= w86 and not w11540;
w11542 <= w90 and not w11541;
w11543 <= w94 and not w11542;
w11544 <= w98 and not w11543;
w11545 <= w102 and not w11544;
w11546 <= w106 and not w11545;
w11547 <= w110 and not w11546;
w11548 <= w114 and not w11547;
w11549 <= w118 and not w11548;
w11550 <= w122 and not w11549;
w11551 <= w126 and not w11550;
w11552 <= w130 and not w11551;
w11553 <= w134 and not w11552;
w11554 <= w138 and not w11553;
w11555 <= w142 and not w11554;
w11556 <= w146 and not w11555;
w11557 <= w150 and not w11556;
w11558 <= w154 and not w11557;
w11559 <= w158 and not w11558;
w11560 <= w162 and not w11559;
w11561 <= w166 and not w11560;
w11562 <= w170 and not w11561;
w11563 <= w174 and not w11562;
w11564 <= w178 and not w11563;
w11565 <= w182 and not w11564;
w11566 <= w186 and not w11565;
w11567 <= w190 and not w11566;
w11568 <= w194 and not w11567;
w11569 <= w198 and not w11568;
w11570 <= w202 and not w11569;
w11571 <= w206 and not w11570;
w11572 <= w210 and not w11571;
w11573 <= w214 and not w11572;
w11574 <= w218 and not w11573;
w11575 <= w222 and not w11574;
w11576 <= w226 and not w11575;
w11577 <= w230 and not w11576;
w11578 <= w234 and not w11577;
w11579 <= w238 and not w11578;
w11580 <= w242 and not w11579;
w11581 <= w246 and not w11580;
w11582 <= w250 and not w11581;
w11583 <= w254 and not w11582;
w11584 <= w258 and not w11583;
w11585 <= w262 and not w11584;
w11586 <= w266 and not w11585;
w11587 <= w270 and not w11586;
w11588 <= w274 and not w11587;
w11589 <= w278 and not w11588;
w11590 <= w282 and not w11589;
w11591 <= w286 and not w11590;
w11592 <= w290 and not w11591;
w11593 <= w294 and not w11592;
w11594 <= w298 and not w11593;
w11595 <= w302 and not w11594;
w11596 <= w306 and not w11595;
w11597 <= w310 and not w11596;
w11598 <= w314 and not w11597;
w11599 <= w318 and not w11598;
w11600 <= w322 and not w11599;
w11601 <= w326 and not w11600;
w11602 <= req(125) and not w328;
w11603 <= not w11601 and w11602;
w11604 <= not w672 and w1097;
w11605 <= w1100 and not w11604;
w11606 <= w1364 and not w11605;
w11607 <= w345 and not w11606;
w11608 <= w349 and not w11607;
w11609 <= w353 and not w11608;
w11610 <= w357 and not w11609;
w11611 <= w361 and not w11610;
w11612 <= w365 and not w11611;
w11613 <= w369 and not w11612;
w11614 <= w373 and not w11613;
w11615 <= w377 and not w11614;
w11616 <= w381 and not w11615;
w11617 <= w385 and not w11616;
w11618 <= w389 and not w11617;
w11619 <= w393 and not w11618;
w11620 <= w397 and not w11619;
w11621 <= w401 and not w11620;
w11622 <= w405 and not w11621;
w11623 <= w409 and not w11622;
w11624 <= w413 and not w11623;
w11625 <= w417 and not w11624;
w11626 <= w421 and not w11625;
w11627 <= w425 and not w11626;
w11628 <= w429 and not w11627;
w11629 <= w433 and not w11628;
w11630 <= w437 and not w11629;
w11631 <= w441 and not w11630;
w11632 <= w445 and not w11631;
w11633 <= w449 and not w11632;
w11634 <= w453 and not w11633;
w11635 <= w457 and not w11634;
w11636 <= w461 and not w11635;
w11637 <= w465 and not w11636;
w11638 <= w469 and not w11637;
w11639 <= w473 and not w11638;
w11640 <= w477 and not w11639;
w11641 <= w481 and not w11640;
w11642 <= w485 and not w11641;
w11643 <= w489 and not w11642;
w11644 <= w493 and not w11643;
w11645 <= w497 and not w11644;
w11646 <= w501 and not w11645;
w11647 <= w505 and not w11646;
w11648 <= w509 and not w11647;
w11649 <= w513 and not w11648;
w11650 <= w517 and not w11649;
w11651 <= w521 and not w11650;
w11652 <= w525 and not w11651;
w11653 <= w529 and not w11652;
w11654 <= w533 and not w11653;
w11655 <= w537 and not w11654;
w11656 <= w541 and not w11655;
w11657 <= w545 and not w11656;
w11658 <= w549 and not w11657;
w11659 <= w553 and not w11658;
w11660 <= w557 and not w11659;
w11661 <= w561 and not w11660;
w11662 <= w565 and not w11661;
w11663 <= w569 and not w11662;
w11664 <= w573 and not w11663;
w11665 <= w577 and not w11664;
w11666 <= w581 and not w11665;
w11667 <= w585 and not w11666;
w11668 <= w589 and not w11667;
w11669 <= w593 and not w11668;
w11670 <= w597 and not w11669;
w11671 <= w601 and not w11670;
w11672 <= w605 and not w11671;
w11673 <= w609 and not w11672;
w11674 <= w613 and not w11673;
w11675 <= w617 and not w11674;
w11676 <= w621 and not w11675;
w11677 <= w625 and not w11676;
w11678 <= w629 and not w11677;
w11679 <= w633 and not w11678;
w11680 <= w637 and not w11679;
w11681 <= w641 and not w11680;
w11682 <= w645 and not w11681;
w11683 <= w649 and not w11682;
w11684 <= w653 and not w11683;
w11685 <= w657 and not w11684;
w11686 <= w661 and not w11685;
w11687 <= w665 and not w11686;
w11688 <= req(126) and not w667;
w11689 <= not w11687 and w11688;
w11690 <= not w1009 and w1187;
w11691 <= w1190 and not w11690;
w11692 <= w1451 and not w11691;
w11693 <= w682 and not w11692;
w11694 <= w686 and not w11693;
w11695 <= w690 and not w11694;
w11696 <= w694 and not w11695;
w11697 <= w698 and not w11696;
w11698 <= w702 and not w11697;
w11699 <= w706 and not w11698;
w11700 <= w710 and not w11699;
w11701 <= w714 and not w11700;
w11702 <= w718 and not w11701;
w11703 <= w722 and not w11702;
w11704 <= w726 and not w11703;
w11705 <= w730 and not w11704;
w11706 <= w734 and not w11705;
w11707 <= w738 and not w11706;
w11708 <= w742 and not w11707;
w11709 <= w746 and not w11708;
w11710 <= w750 and not w11709;
w11711 <= w754 and not w11710;
w11712 <= w758 and not w11711;
w11713 <= w762 and not w11712;
w11714 <= w766 and not w11713;
w11715 <= w770 and not w11714;
w11716 <= w774 and not w11715;
w11717 <= w778 and not w11716;
w11718 <= w782 and not w11717;
w11719 <= w786 and not w11718;
w11720 <= w790 and not w11719;
w11721 <= w794 and not w11720;
w11722 <= w798 and not w11721;
w11723 <= w802 and not w11722;
w11724 <= w806 and not w11723;
w11725 <= w810 and not w11724;
w11726 <= w814 and not w11725;
w11727 <= w818 and not w11726;
w11728 <= w822 and not w11727;
w11729 <= w826 and not w11728;
w11730 <= w830 and not w11729;
w11731 <= w834 and not w11730;
w11732 <= w838 and not w11731;
w11733 <= w842 and not w11732;
w11734 <= w846 and not w11733;
w11735 <= w850 and not w11734;
w11736 <= w854 and not w11735;
w11737 <= w858 and not w11736;
w11738 <= w862 and not w11737;
w11739 <= w866 and not w11738;
w11740 <= w870 and not w11739;
w11741 <= w874 and not w11740;
w11742 <= w878 and not w11741;
w11743 <= w882 and not w11742;
w11744 <= w886 and not w11743;
w11745 <= w890 and not w11744;
w11746 <= w894 and not w11745;
w11747 <= w898 and not w11746;
w11748 <= w902 and not w11747;
w11749 <= w906 and not w11748;
w11750 <= w910 and not w11749;
w11751 <= w914 and not w11750;
w11752 <= w918 and not w11751;
w11753 <= w922 and not w11752;
w11754 <= w926 and not w11753;
w11755 <= w930 and not w11754;
w11756 <= w934 and not w11755;
w11757 <= w938 and not w11756;
w11758 <= w942 and not w11757;
w11759 <= w946 and not w11758;
w11760 <= w950 and not w11759;
w11761 <= w954 and not w11760;
w11762 <= w958 and not w11761;
w11763 <= w962 and not w11762;
w11764 <= w966 and not w11763;
w11765 <= w970 and not w11764;
w11766 <= w974 and not w11765;
w11767 <= w978 and not w11766;
w11768 <= w982 and not w11767;
w11769 <= w986 and not w11768;
w11770 <= w990 and not w11769;
w11771 <= w994 and not w11770;
w11772 <= w998 and not w11771;
w11773 <= w1002 and not w11772;
w11774 <= req(127) and not w1004;
w11775 <= not w11773 and w11774;
w11776 <= w2 and w17;
w11777 <= w33 and w49;
w11778 <= w65 and w81;
w11779 <= w97 and w113;
w11780 <= w129 and w145;
w11781 <= w161 and w177;
w11782 <= w193 and w209;
w11783 <= w225 and w241;
w11784 <= w257 and w273;
w11785 <= w289 and w305;
w11786 <= w321 and w348;
w11787 <= w364 and w380;
w11788 <= w396 and w412;
w11789 <= w428 and w444;
w11790 <= w460 and w476;
w11791 <= w492 and w508;
w11792 <= w524 and w540;
w11793 <= w556 and w572;
w11794 <= w588 and w604;
w11795 <= w620 and w636;
w11796 <= w652 and w668;
w11797 <= w678 and w693;
w11798 <= w709 and w725;
w11799 <= w741 and w757;
w11800 <= w773 and w789;
w11801 <= w805 and w821;
w11802 <= w837 and w853;
w11803 <= w869 and w885;
w11804 <= w901 and w917;
w11805 <= w933 and w949;
w11806 <= w965 and w981;
w11807 <= w997 and w1097;
w11808 <= w11806 and w11807;
w11809 <= w11804 and w11805;
w11810 <= w11802 and w11803;
w11811 <= w11800 and w11801;
w11812 <= w11798 and w11799;
w11813 <= w11796 and w11797;
w11814 <= w11794 and w11795;
w11815 <= w11792 and w11793;
w11816 <= w11790 and w11791;
w11817 <= w11788 and w11789;
w11818 <= w11786 and w11787;
w11819 <= w11784 and w11785;
w11820 <= w11782 and w11783;
w11821 <= w11780 and w11781;
w11822 <= w11778 and w11779;
w11823 <= w11776 and w11777;
w11824 <= w11822 and w11823;
w11825 <= w11820 and w11821;
w11826 <= w11818 and w11819;
w11827 <= w11816 and w11817;
w11828 <= w11814 and w11815;
w11829 <= w11812 and w11813;
w11830 <= w11810 and w11811;
w11831 <= w11808 and w11809;
w11832 <= w11830 and w11831;
w11833 <= w11828 and w11829;
w11834 <= w11826 and w11827;
w11835 <= w11824 and w11825;
w11836 <= w11834 and w11835;
w11837 <= w11832 and w11833;
w11838 <= w11836 and w11837;
one <= '1';
grant(0) <= w338;-- level 87
grant(1) <= w677;-- level 87
grant(2) <= w1014;-- level 87
grant(3) <= w1104;-- level 87
grant(4) <= w1194;-- level 87
grant(5) <= w1281;-- level 87
grant(6) <= w1368;-- level 87
grant(7) <= w1455;-- level 87
grant(8) <= w1541;-- level 87
grant(9) <= w1627;-- level 87
grant(10) <= w1713;-- level 87
grant(11) <= w1799;-- level 87
grant(12) <= w1885;-- level 87
grant(13) <= w1971;-- level 87
grant(14) <= w2057;-- level 87
grant(15) <= w2143;-- level 87
grant(16) <= w2229;-- level 87
grant(17) <= w2315;-- level 87
grant(18) <= w2401;-- level 87
grant(19) <= w2487;-- level 87
grant(20) <= w2573;-- level 87
grant(21) <= w2659;-- level 87
grant(22) <= w2745;-- level 87
grant(23) <= w2831;-- level 87
grant(24) <= w2917;-- level 87
grant(25) <= w3003;-- level 87
grant(26) <= w3089;-- level 87
grant(27) <= w3175;-- level 87
grant(28) <= w3261;-- level 87
grant(29) <= w3347;-- level 87
grant(30) <= w3433;-- level 87
grant(31) <= w3519;-- level 87
grant(32) <= w3605;-- level 87
grant(33) <= w3691;-- level 87
grant(34) <= w3777;-- level 87
grant(35) <= w3863;-- level 87
grant(36) <= w3949;-- level 87
grant(37) <= w4035;-- level 87
grant(38) <= w4121;-- level 87
grant(39) <= w4207;-- level 87
grant(40) <= w4293;-- level 87
grant(41) <= w4379;-- level 87
grant(42) <= w4465;-- level 87
grant(43) <= w4551;-- level 87
grant(44) <= w4637;-- level 87
grant(45) <= w4723;-- level 87
grant(46) <= w4809;-- level 87
grant(47) <= w4895;-- level 87
grant(48) <= w4981;-- level 87
grant(49) <= w5067;-- level 87
grant(50) <= w5153;-- level 87
grant(51) <= w5239;-- level 87
grant(52) <= w5325;-- level 87
grant(53) <= w5411;-- level 87
grant(54) <= w5497;-- level 87
grant(55) <= w5583;-- level 87
grant(56) <= w5669;-- level 87
grant(57) <= w5755;-- level 87
grant(58) <= w5841;-- level 87
grant(59) <= w5927;-- level 87
grant(60) <= w6013;-- level 87
grant(61) <= w6099;-- level 87
grant(62) <= w6185;-- level 87
grant(63) <= w6271;-- level 87
grant(64) <= w6357;-- level 87
grant(65) <= w6443;-- level 87
grant(66) <= w6529;-- level 87
grant(67) <= w6615;-- level 87
grant(68) <= w6701;-- level 87
grant(69) <= w6787;-- level 87
grant(70) <= w6873;-- level 87
grant(71) <= w6959;-- level 87
grant(72) <= w7045;-- level 87
grant(73) <= w7131;-- level 87
grant(74) <= w7217;-- level 87
grant(75) <= w7303;-- level 87
grant(76) <= w7389;-- level 87
grant(77) <= w7475;-- level 87
grant(78) <= w7561;-- level 87
grant(79) <= w7647;-- level 87
grant(80) <= w7733;-- level 87
grant(81) <= w7819;-- level 87
grant(82) <= w7905;-- level 87
grant(83) <= w7991;-- level 87
grant(84) <= w8077;-- level 87
grant(85) <= w8163;-- level 87
grant(86) <= w8249;-- level 87
grant(87) <= w8335;-- level 87
grant(88) <= w8421;-- level 87
grant(89) <= w8507;-- level 87
grant(90) <= w8593;-- level 87
grant(91) <= w8679;-- level 87
grant(92) <= w8765;-- level 87
grant(93) <= w8851;-- level 87
grant(94) <= w8937;-- level 87
grant(95) <= w9023;-- level 87
grant(96) <= w9109;-- level 87
grant(97) <= w9195;-- level 87
grant(98) <= w9281;-- level 87
grant(99) <= w9367;-- level 87
grant(100) <= w9453;-- level 87
grant(101) <= w9539;-- level 87
grant(102) <= w9625;-- level 87
grant(103) <= w9711;-- level 87
grant(104) <= w9797;-- level 87
grant(105) <= w9883;-- level 87
grant(106) <= w9969;-- level 87
grant(107) <= w10055;-- level 87
grant(108) <= w10141;-- level 87
grant(109) <= w10227;-- level 87
grant(110) <= w10313;-- level 87
grant(111) <= w10399;-- level 87
grant(112) <= w10485;-- level 87
grant(113) <= w10571;-- level 87
grant(114) <= w10657;-- level 87
grant(115) <= w10743;-- level 87
grant(116) <= w10829;-- level 87
grant(117) <= w10915;-- level 87
grant(118) <= w11001;-- level 87
grant(119) <= w11087;-- level 87
grant(120) <= w11173;-- level 87
grant(121) <= w11259;-- level 87
grant(122) <= w11345;-- level 87
grant(123) <= w11431;-- level 87
grant(124) <= w11517;-- level 87
grant(125) <= w11603;-- level 87
grant(126) <= w11689;-- level 87
grant(127) <= w11775;-- level 87
anyGrant <= not w11838;-- level 7
end Behavioral;