
	`include "spi_if.sv";
	`include "apb_if.sv";

package proj_pkg;


endpackage
