module top;

import "DPI" function void string_sv2c(); 

initial 
begin 
    string_sv2c(); 
end 

endmodule
