`ifdef ATCPIT100_CFG_VH
`else
`define ATCPIT100_CFG_VH

//-------------------------------------------------
// Number of PIT Channels
//-------------------------------------------------
//`define ATCPIT100_NUM_CHANNEL_1
//`define ATCPIT100_NUM_CHANNEL_2
//`define ATCPIT100_NUM_CHANNEL_3
`define ATCPIT100_NUM_CHANNEL_4

`endif // ATCPIT100_CFG_VH
