library ieee;
use ieee.std_logic_1164.all;

entity top is
	port( a: in std_logic_vector(63 downto 0);
	asquared: out std_logic_vector(127 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483: std_logic;

begin

w0 <= a(0) and a(1);
w1 <= a(1) and not w0;
w2 <= a(0) and a(2);
w3 <= w0 and w2;
w4 <= not w0 and not w2;
w5 <= not w3 and not w4;
w6 <= a(1) and a(2);
w7 <= a(2) and not w6;
w8 <= a(0) and a(3);
w9 <= not w7 and not w8;
w10 <= w7 and w8;
w11 <= not w9 and not w10;
w12 <= w3 and not w11;
w13 <= not w3 and w11;
w14 <= not w12 and not w13;
w15 <= a(3) and a(4);
w16 <= w0 and w15;
w17 <= a(1) and a(3);
w18 <= a(0) and a(4);
w19 <= not w17 and not w18;
w20 <= not w16 and not w19;
w21 <= not w6 and not w20;
w22 <= w6 and w20;
w23 <= not w21 and not w22;
w24 <= a(2) and a(3);
w25 <= a(0) and w24;
w26 <= not w23 and not w25;
w27 <= w23 and w25;
w28 <= not w26 and not w27;
w29 <= a(1) and a(4);
w30 <= a(0) and a(5);
w31 <= not w29 and not w30;
w32 <= a(4) and a(5);
w33 <= w0 and w32;
w34 <= not w31 and not w33;
w35 <= w16 and w34;
w36 <= not w33 and not w35;
w37 <= not w31 and w36;
w38 <= w16 and not w35;
w39 <= not w37 and not w38;
w40 <= a(3) and not w24;
w41 <= w39 and not w40;
w42 <= not w39 and w40;
w43 <= not w41 and not w42;
w44 <= not w21 and w25;
w45 <= not w22 and not w44;
w46 <= not w43 and w45;
w47 <= w43 and not w45;
w48 <= not w46 and not w47;
w49 <= not w41 and not w45;
w50 <= not w42 and not w49;
w51 <= a(6) and w25;
w52 <= a(0) and not w51;
w53 <= a(6) and w52;
w54 <= w24 and not w51;
w55 <= not w53 and not w54;
w56 <= w6 and w32;
w57 <= a(1) and a(5);
w58 <= a(2) and a(4);
w59 <= not w57 and not w58;
w60 <= not w56 and not w59;
w61 <= w55 and not w60;
w62 <= not w55 and w60;
w63 <= not w61 and not w62;
w64 <= w36 and not w63;
w65 <= not w36 and w63;
w66 <= not w64 and not w65;
w67 <= w50 and not w66;
w68 <= not w50 and not w64;
w69 <= not w65 and w68;
w70 <= not w67 and not w69;
w71 <= w24 and w32;
w72 <= a(0) and a(7);
w73 <= w15 and w72;
w74 <= a(5) and a(7);
w75 <= w2 and w74;
w76 <= not w73 and not w75;
w77 <= not w71 and not w76;
w78 <= not w71 and not w77;
w79 <= a(2) and a(5);
w80 <= not w15 and not w79;
w81 <= w78 and not w80;
w82 <= w72 and not w77;
w83 <= not w81 and not w82;
w84 <= not w51 and not w62;
w85 <= a(1) and a(6);
w86 <= w56 and not w85;
w87 <= w56 and not w86;
w88 <= not a(4) and not w85;
w89 <= a(4) and w85;
w90 <= not w86 and not w89;
w91 <= not w88 and w90;
w92 <= not w87 and not w91;
w93 <= not w84 and not w92;
w94 <= w84 and not w91;
w95 <= not w87 and w94;
w96 <= not w93 and not w95;
w97 <= w83 and not w96;
w98 <= not w83 and w96;
w99 <= not w97 and not w98;
w100 <= not w65 and not w68;
w101 <= not w99 and w100;
w102 <= w99 and not w100;
w103 <= not w101 and not w102;
w104 <= not w86 and not w93;
w105 <= a(1) and a(7);
w106 <= a(3) and a(5);
w107 <= w105 and w106;
w108 <= w105 and not w107;
w109 <= w106 and not w107;
w110 <= not w108 and not w109;
w111 <= not w78 and not w110;
w112 <= not w78 and not w111;
w113 <= not w110 and not w111;
w114 <= not w112 and not w113;
w115 <= a(0) and a(8);
w116 <= a(2) and a(6);
w117 <= not w115 and not w116;
w118 <= a(6) and a(8);
w119 <= w2 and w118;
w120 <= not w117 and not w119;
w121 <= w89 and w120;
w122 <= not w119 and not w121;
w123 <= not w117 and w122;
w124 <= w89 and not w121;
w125 <= not w123 and not w124;
w126 <= not w114 and not w125;
w127 <= w114 and w125;
w128 <= not w126 and not w127;
w129 <= w104 and not w128;
w130 <= not w104 and w128;
w131 <= not w129 and not w130;
w132 <= not w97 and not w100;
w133 <= not w98 and not w132;
w134 <= not w131 and w133;
w135 <= w131 and not w133;
w136 <= not w134 and not w135;
w137 <= not w111 and not w126;
w138 <= a(5) and a(6);
w139 <= w15 and w138;
w140 <= w58 and w74;
w141 <= a(6) and a(7);
w142 <= w24 and w141;
w143 <= not w140 and not w142;
w144 <= not w139 and not w143;
w145 <= not w139 and not w144;
w146 <= a(3) and a(6);
w147 <= not w32 and not w146;
w148 <= w145 and not w147;
w149 <= a(2) and a(7);
w150 <= not w144 and w149;
w151 <= not w148 and not w150;
w152 <= not w122 and not w151;
w153 <= not w122 and not w152;
w154 <= not w151 and not w152;
w155 <= not w153 and not w154;
w156 <= a(0) and a(9);
w157 <= w107 and not w156;
w158 <= not w107 and w156;
w159 <= not w157 and not w158;
w160 <= a(5) and a(8);
w161 <= a(1) and w160;
w162 <= a(5) and not w161;
w163 <= a(1) and not w161;
w164 <= a(8) and w163;
w165 <= not w162 and not w164;
w166 <= not w159 and not w165;
w167 <= w159 and w165;
w168 <= not w166 and not w167;
w169 <= not w155 and w168;
w170 <= not w154 and not w168;
w171 <= not w153 and w170;
w172 <= not w169 and not w171;
w173 <= not w137 and w172;
w174 <= w137 and not w172;
w175 <= not w173 and not w174;
w176 <= not w129 and not w133;
w177 <= not w130 and not w176;
w178 <= not w175 and w177;
w179 <= w175 and not w177;
w180 <= not w178 and not w179;
w181 <= not w174 and not w177;
w182 <= not w173 and not w181;
w183 <= not w152 and not w169;
w184 <= a(8) and a(10);
w185 <= w2 and w184;
w186 <= a(7) and a(8);
w187 <= w24 and w186;
w188 <= not w185 and not w187;
w189 <= a(0) and a(10);
w190 <= a(3) and a(7);
w191 <= w189 and w190;
w192 <= not w188 and not w191;
w193 <= a(2) and not w192;
w194 <= a(8) and w193;
w195 <= not w191 and not w192;
w196 <= not w189 and not w190;
w197 <= w195 and not w196;
w198 <= not w194 and not w197;
w199 <= w107 and w156;
w200 <= not w166 and not w199;
w201 <= not w198 and w200;
w202 <= w198 and not w200;
w203 <= not w201 and not w202;
w204 <= a(9) and w89;
w205 <= a(1) and a(9);
w206 <= a(4) and a(6);
w207 <= not w205 and not w206;
w208 <= not w204 and not w207;
w209 <= w161 and w208;
w210 <= w161 and not w209;
w211 <= w208 and not w209;
w212 <= not w210 and not w211;
w213 <= not w145 and not w212;
w214 <= w145 and not w211;
w215 <= not w210 and w214;
w216 <= not w213 and not w215;
w217 <= not w203 and w216;
w218 <= w203 and not w216;
w219 <= not w217 and not w218;
w220 <= w183 and not w219;
w221 <= not w183 and w219;
w222 <= not w220 and not w221;
w223 <= w182 and not w222;
w224 <= not w182 and not w220;
w225 <= not w221 and w224;
w226 <= not w223 and not w225;
w227 <= not w198 and not w200;
w228 <= not w217 and not w227;
w229 <= a(10) and w85;
w230 <= a(6) and not w229;
w231 <= a(1) and not w229;
w232 <= a(10) and w231;
w233 <= not w230 and not w232;
w234 <= not w195 and not w233;
w235 <= not w195 and not w234;
w236 <= not w233 and not w234;
w237 <= not w235 and not w236;
w238 <= a(8) and a(9);
w239 <= w24 and w238;
w240 <= a(2) and a(9);
w241 <= a(3) and a(8);
w242 <= not w240 and not w241;
w243 <= not w239 and not w242;
w244 <= w204 and w243;
w245 <= w204 and not w244;
w246 <= not w239 and not w244;
w247 <= not w242 and w246;
w248 <= not w245 and not w247;
w249 <= not w237 and not w248;
w250 <= not w237 and not w249;
w251 <= not w248 and not w249;
w252 <= not w250 and not w251;
w253 <= not w209 and not w213;
w254 <= w32 and w141;
w255 <= a(0) and a(11);
w256 <= a(4) and a(7);
w257 <= not w138 and not w256;
w258 <= not w254 and not w257;
w259 <= w255 and w258;
w260 <= not w254 and not w259;
w261 <= not w257 and w260;
w262 <= w255 and not w259;
w263 <= not w261 and not w262;
w264 <= not w253 and not w263;
w265 <= not w253 and not w264;
w266 <= not w263 and not w264;
w267 <= not w265 and not w266;
w268 <= not w252 and not w267;
w269 <= w252 and not w266;
w270 <= not w265 and w269;
w271 <= not w268 and not w270;
w272 <= w228 and not w271;
w273 <= not w228 and w271;
w274 <= not w272 and not w273;
w275 <= not w221 and not w224;
w276 <= not w274 and w275;
w277 <= w274 and not w275;
w278 <= not w276 and not w277;
w279 <= not w272 and not w275;
w280 <= not w273 and not w279;
w281 <= not w264 and not w268;
w282 <= w246 and w260;
w283 <= not w246 and not w260;
w284 <= not w282 and not w283;
w285 <= a(3) and a(9);
w286 <= a(10) and a(12);
w287 <= w2 and w286;
w288 <= a(0) and a(12);
w289 <= w285 and w288;
w290 <= a(9) and a(10);
w291 <= w24 and w290;
w292 <= not w289 and not w291;
w293 <= not w287 and not w292;
w294 <= w285 and not w293;
w295 <= not w287 and not w293;
w296 <= a(2) and a(10);
w297 <= not w288 and not w296;
w298 <= w295 and not w297;
w299 <= not w294 and not w298;
w300 <= w284 and not w299;
w301 <= w284 and not w300;
w302 <= not w299 and not w300;
w303 <= not w301 and not w302;
w304 <= not w234 and not w249;
w305 <= a(4) and a(8);
w306 <= not w229 and not w305;
w307 <= w229 and w305;
w308 <= a(5) and a(11);
w309 <= w105 and w308;
w310 <= a(1) and a(11);
w311 <= not w74 and not w310;
w312 <= not w309 and not w311;
w313 <= not w307 and w312;
w314 <= not w306 and w313;
w315 <= not w307 and not w314;
w316 <= not w306 and w315;
w317 <= w312 and not w314;
w318 <= not w316 and not w317;
w319 <= not w304 and not w318;
w320 <= w304 and w318;
w321 <= not w319 and not w320;
w322 <= not w303 and w321;
w323 <= w303 and not w321;
w324 <= not w322 and not w323;
w325 <= w281 and not w324;
w326 <= not w281 and w324;
w327 <= not w325 and not w326;
w328 <= w280 and not w327;
w329 <= not w280 and not w325;
w330 <= not w326 and w329;
w331 <= not w328 and not w330;
w332 <= a(9) and a(13);
w333 <= w18 and w332;
w334 <= w15 and w290;
w335 <= a(3) and a(13);
w336 <= w189 and w335;
w337 <= not w334 and not w336;
w338 <= not w333 and not w337;
w339 <= a(3) and not w338;
w340 <= a(10) and w339;
w341 <= not w333 and not w338;
w342 <= a(0) and a(13);
w343 <= a(4) and a(9);
w344 <= not w342 and not w343;
w345 <= w341 and not w344;
w346 <= not w340 and not w345;
w347 <= w315 and not w346;
w348 <= not w315 and w346;
w349 <= not w347 and not w348;
w350 <= a(2) and a(11);
w351 <= not w141 and not w160;
w352 <= w138 and w186;
w353 <= w350 and not w352;
w354 <= not w351 and w353;
w355 <= w350 and not w354;
w356 <= not w352 and not w354;
w357 <= not w351 and w356;
w358 <= not w355 and not w357;
w359 <= not w349 and not w358;
w360 <= w349 and w358;
w361 <= not w359 and not w360;
w362 <= not w283 and not w300;
w363 <= not a(12) and w309;
w364 <= a(12) and w105;
w365 <= a(1) and a(12);
w366 <= not a(7) and not w365;
w367 <= not w364 and not w366;
w368 <= not w309 and not w367;
w369 <= not w363 and not w368;
w370 <= not w295 and w369;
w371 <= w295 and not w369;
w372 <= not w370 and not w371;
w373 <= w362 and not w372;
w374 <= not w362 and w372;
w375 <= not w373 and not w374;
w376 <= not w319 and not w322;
w377 <= not w375 and w376;
w378 <= w375 and not w376;
w379 <= not w377 and not w378;
w380 <= not w361 and not w379;
w381 <= w361 and w379;
w382 <= not w380 and not w381;
w383 <= not w326 and not w329;
w384 <= not w382 and w383;
w385 <= w382 and not w383;
w386 <= not w384 and not w385;
w387 <= not w380 and not w383;
w388 <= not w381 and not w387;
w389 <= not w374 and not w378;
w390 <= a(1) and a(13);
w391 <= not w118 and not w390;
w392 <= w118 and w390;
w393 <= not w356 and not w392;
w394 <= not w391 and w393;
w395 <= not w356 and not w394;
w396 <= not w392 and not w394;
w397 <= not w391 and w396;
w398 <= not w395 and not w397;
w399 <= not w341 and not w398;
w400 <= not w341 and not w399;
w401 <= not w398 and not w399;
w402 <= not w400 and not w401;
w403 <= not w315 and not w346;
w404 <= not w359 and not w403;
w405 <= w402 and w404;
w406 <= not w402 and not w404;
w407 <= not w405 and not w406;
w408 <= a(11) and a(12);
w409 <= w24 and w408;
w410 <= a(3) and a(14);
w411 <= w255 and w410;
w412 <= a(12) and a(14);
w413 <= w2 and w412;
w414 <= not w411 and not w413;
w415 <= not w409 and not w414;
w416 <= not w409 and not w415;
w417 <= a(2) and a(12);
w418 <= a(3) and a(11);
w419 <= not w417 and not w418;
w420 <= w416 and not w419;
w421 <= a(14) and not w415;
w422 <= a(0) and w421;
w423 <= not w420 and not w422;
w424 <= w32 and w290;
w425 <= a(4) and a(10);
w426 <= a(5) and a(9);
w427 <= not w425 and not w426;
w428 <= not w424 and not w427;
w429 <= w364 and w428;
w430 <= w364 and not w429;
w431 <= not w424 and not w429;
w432 <= not w427 and w431;
w433 <= not w430 and not w432;
w434 <= not w423 and not w433;
w435 <= not w423 and not w434;
w436 <= not w433 and not w434;
w437 <= not w435 and not w436;
w438 <= not w363 and not w370;
w439 <= w437 and w438;
w440 <= not w437 and not w438;
w441 <= not w439 and not w440;
w442 <= w407 and not w441;
w443 <= not w407 and w441;
w444 <= not w442 and not w443;
w445 <= not w389 and not w444;
w446 <= w389 and w444;
w447 <= not w445 and not w446;
w448 <= w388 and not w447;
w449 <= not w388 and not w446;
w450 <= not w445 and w449;
w451 <= not w448 and not w450;
w452 <= not w445 and not w449;
w453 <= w407 and w441;
w454 <= not w406 and not w453;
w455 <= a(4) and a(11);
w456 <= not w392 and not w455;
w457 <= w392 and w455;
w458 <= a(1) and a(14);
w459 <= a(8) and not w458;
w460 <= not a(8) and w458;
w461 <= not w459 and not w460;
w462 <= not w457 and not w461;
w463 <= not w456 and w462;
w464 <= not w457 and not w463;
w465 <= not w456 and w464;
w466 <= not w461 and not w463;
w467 <= not w465 and not w466;
w468 <= a(6) and a(9);
w469 <= not w186 and not w468;
w470 <= w186 and w468;
w471 <= a(2) and not w470;
w472 <= a(13) and w471;
w473 <= not w469 and w472;
w474 <= a(13) and not w473;
w475 <= a(2) and w474;
w476 <= not w470 and not w473;
w477 <= not w469 and w476;
w478 <= not w475 and not w477;
w479 <= not w467 and not w478;
w480 <= not w467 and not w479;
w481 <= not w478 and not w479;
w482 <= not w480 and not w481;
w483 <= not w394 and not w399;
w484 <= w482 and w483;
w485 <= not w482 and not w483;
w486 <= not w484 and not w485;
w487 <= w416 and w431;
w488 <= not w416 and not w431;
w489 <= not w487 and not w488;
w490 <= a(5) and a(10);
w491 <= a(10) and a(15);
w492 <= a(0) and w491;
w493 <= a(3) and w286;
w494 <= not w492 and not w493;
w495 <= a(0) and a(15);
w496 <= a(3) and a(12);
w497 <= w495 and w496;
w498 <= a(5) and not w497;
w499 <= not w494 and w498;
w500 <= w490 and not w499;
w501 <= not w497 and not w499;
w502 <= not w495 and not w496;
w503 <= w501 and not w502;
w504 <= not w500 and not w503;
w505 <= w489 and not w504;
w506 <= w489 and not w505;
w507 <= not w504 and not w505;
w508 <= not w506 and not w507;
w509 <= not w434 and not w440;
w510 <= w508 and w509;
w511 <= not w508 and not w509;
w512 <= not w510 and not w511;
w513 <= w486 and not w512;
w514 <= not w486 and w512;
w515 <= not w513 and not w514;
w516 <= not w454 and not w515;
w517 <= w454 and w515;
w518 <= not w516 and not w517;
w519 <= not w452 and not w518;
w520 <= w452 and w518;
w521 <= not w519 and not w520;
w522 <= w486 and w512;
w523 <= not w511 and not w522;
w524 <= w464 and w501;
w525 <= not w464 and not w501;
w526 <= not w524 and not w525;
w527 <= a(6) and a(16);
w528 <= w189 and w527;
w529 <= a(10) and a(11);
w530 <= w138 and w529;
w531 <= a(0) and a(16);
w532 <= w308 and w531;
w533 <= not w530 and not w532;
w534 <= not w528 and not w533;
w535 <= w308 and not w534;
w536 <= not w528 and not w534;
w537 <= a(6) and a(10);
w538 <= not w531 and not w537;
w539 <= w536 and not w538;
w540 <= not w535 and not w539;
w541 <= w526 and not w540;
w542 <= w526 and not w541;
w543 <= not w540 and not w541;
w544 <= not w542 and not w543;
w545 <= not w479 and not w485;
w546 <= w544 and w545;
w547 <= not w544 and not w545;
w548 <= not w546 and not w547;
w549 <= not w488 and not w505;
w550 <= a(4) and a(12);
w551 <= a(13) and a(14);
w552 <= w24 and w551;
w553 <= w58 and w412;
w554 <= a(12) and a(13);
w555 <= w15 and w554;
w556 <= not w553 and not w555;
w557 <= not w552 and not w556;
w558 <= w550 and not w557;
w559 <= not w552 and not w557;
w560 <= a(2) and a(14);
w561 <= not w335 and not w560;
w562 <= w559 and not w561;
w563 <= not w558 and not w562;
w564 <= not w549 and not w563;
w565 <= not w549 and not w564;
w566 <= not w563 and not w564;
w567 <= not w565 and not w566;
w568 <= a(8) and w458;
w569 <= a(7) and a(9);
w570 <= a(1) and a(15);
w571 <= w569 and w570;
w572 <= not w569 and not w570;
w573 <= not w571 and not w572;
w574 <= w568 and w573;
w575 <= w568 and not w574;
w576 <= not w568 and w573;
w577 <= not w575 and not w576;
w578 <= not w476 and not w577;
w579 <= not w476 and not w578;
w580 <= not w577 and not w578;
w581 <= not w579 and not w580;
w582 <= not w567 and not w581;
w583 <= not w567 and not w582;
w584 <= not w581 and not w582;
w585 <= not w583 and not w584;
w586 <= not w548 and w585;
w587 <= w548 and not w585;
w588 <= not w586 and not w587;
w589 <= not w523 and w588;
w590 <= w523 and not w588;
w591 <= not w589 and not w590;
w592 <= not w452 and not w517;
w593 <= not w516 and not w592;
w594 <= not w591 and w593;
w595 <= w591 and not w593;
w596 <= not w594 and not w595;
w597 <= not w547 and not w587;
w598 <= a(5) and a(12);
w599 <= a(0) and a(17);
w600 <= not w598 and not w599;
w601 <= w598 and w599;
w602 <= not w600 and not w601;
w603 <= w571 and w602;
w604 <= not w601 and not w603;
w605 <= not w600 and w604;
w606 <= w571 and not w603;
w607 <= not w605 and not w606;
w608 <= a(7) and a(10);
w609 <= not w238 and not w608;
w610 <= w186 and w290;
w611 <= w410 and not w610;
w612 <= not w609 and w611;
w613 <= w410 and not w612;
w614 <= not w610 and not w612;
w615 <= not w609 and w614;
w616 <= not w613 and not w615;
w617 <= not w607 and not w616;
w618 <= not w607 and not w617;
w619 <= not w616 and not w617;
w620 <= not w618 and not w619;
w621 <= a(6) and a(11);
w622 <= a(11) and a(15);
w623 <= a(2) and w622;
w624 <= a(11) and a(13);
w625 <= a(4) and w624;
w626 <= not w623 and not w625;
w627 <= a(13) and a(15);
w628 <= w58 and w627;
w629 <= a(6) and not w628;
w630 <= not w626 and w629;
w631 <= w621 and not w630;
w632 <= not w628 and not w630;
w633 <= a(2) and a(15);
w634 <= a(4) and a(13);
w635 <= not w633 and not w634;
w636 <= w632 and not w635;
w637 <= not w631 and not w636;
w638 <= not w620 and not w637;
w639 <= not w620 and not w638;
w640 <= not w637 and not w638;
w641 <= not w639 and not w640;
w642 <= not w564 and not w582;
w643 <= w641 and w642;
w644 <= not w641 and not w642;
w645 <= not w643 and not w644;
w646 <= not w574 and not w578;
w647 <= not w525 and not w541;
w648 <= w646 and w647;
w649 <= not w646 and not w647;
w650 <= not w648 and not w649;
w651 <= a(1) and a(16);
w652 <= not a(9) and not w651;
w653 <= a(9) and a(16);
w654 <= a(1) and w653;
w655 <= not w559 and not w654;
w656 <= not w652 and w655;
w657 <= not w559 and not w656;
w658 <= not w654 and not w656;
w659 <= not w652 and w658;
w660 <= not w657 and not w659;
w661 <= not w536 and not w660;
w662 <= not w536 and not w661;
w663 <= not w660 and not w661;
w664 <= not w662 and not w663;
w665 <= not w650 and w664;
w666 <= w650 and not w664;
w667 <= not w665 and not w666;
w668 <= w645 and w667;
w669 <= not w645 and not w667;
w670 <= not w668 and not w669;
w671 <= not w597 and w670;
w672 <= w597 and not w670;
w673 <= not w671 and not w672;
w674 <= not w590 and not w593;
w675 <= not w589 and not w674;
w676 <= not w673 and w675;
w677 <= w673 and not w675;
w678 <= not w676 and not w677;
w679 <= not w672 and not w675;
w680 <= not w671 and not w679;
w681 <= not w644 and not w668;
w682 <= a(7) and a(18);
w683 <= w255 and w682;
w684 <= w74 and w624;
w685 <= not w683 and not w684;
w686 <= a(0) and a(18);
w687 <= a(5) and a(13);
w688 <= w686 and w687;
w689 <= not w685 and not w688;
w690 <= not w688 and not w689;
w691 <= not w686 and not w687;
w692 <= w690 and not w691;
w693 <= a(11) and not w689;
w694 <= a(7) and w693;
w695 <= not w692 and not w694;
w696 <= a(4) and a(14);
w697 <= a(15) and a(16);
w698 <= w24 and w697;
w699 <= a(14) and a(16);
w700 <= w58 and w699;
w701 <= a(14) and a(15);
w702 <= w15 and w701;
w703 <= not w700 and not w702;
w704 <= not w698 and not w703;
w705 <= w696 and not w704;
w706 <= not w698 and not w704;
w707 <= a(3) and a(15);
w708 <= a(2) and a(16);
w709 <= not w707 and not w708;
w710 <= w706 and not w709;
w711 <= not w705 and not w710;
w712 <= not w695 and not w711;
w713 <= not w695 and not w712;
w714 <= not w711 and not w712;
w715 <= not w713 and not w714;
w716 <= a(1) and a(17);
w717 <= w184 and w716;
w718 <= w184 and not w717;
w719 <= not w184 and w716;
w720 <= not w718 and not w719;
w721 <= a(6) and a(12);
w722 <= not w654 and not w721;
w723 <= w654 and w721;
w724 <= not w720 and not w723;
w725 <= not w722 and w724;
w726 <= not w720 and not w725;
w727 <= not w723 and not w725;
w728 <= not w722 and w727;
w729 <= not w726 and not w728;
w730 <= not w715 and not w729;
w731 <= not w715 and not w730;
w732 <= not w729 and not w730;
w733 <= not w731 and not w732;
w734 <= not w649 and not w666;
w735 <= not w733 and not w734;
w736 <= not w733 and not w735;
w737 <= not w734 and not w735;
w738 <= not w736 and not w737;
w739 <= w614 and w632;
w740 <= not w614 and not w632;
w741 <= not w739 and not w740;
w742 <= w604 and not w741;
w743 <= not w604 and w741;
w744 <= not w742 and not w743;
w745 <= not w656 and not w661;
w746 <= not w617 and not w638;
w747 <= w745 and w746;
w748 <= not w745 and not w746;
w749 <= not w747 and not w748;
w750 <= w744 and w749;
w751 <= not w744 and not w749;
w752 <= not w750 and not w751;
w753 <= not w738 and w752;
w754 <= w738 and not w752;
w755 <= not w753 and not w754;
w756 <= not w681 and w755;
w757 <= w681 and not w755;
w758 <= not w756 and not w757;
w759 <= w680 and not w758;
w760 <= not w680 and not w757;
w761 <= not w756 and w760;
w762 <= not w759 and not w761;
w763 <= w690 and w727;
w764 <= not w690 and not w727;
w765 <= not w763 and not w764;
w766 <= a(3) and a(16);
w767 <= a(8) and a(11);
w768 <= not w290 and not w767;
w769 <= w290 and w767;
w770 <= w766 and not w769;
w771 <= not w768 and w770;
w772 <= w766 and not w771;
w773 <= not w769 and not w771;
w774 <= not w768 and w773;
w775 <= not w772 and not w774;
w776 <= w765 and not w775;
w777 <= w765 and not w776;
w778 <= not w775 and not w776;
w779 <= not w777 and not w778;
w780 <= not w712 and not w730;
w781 <= a(1) and a(18);
w782 <= w717 and not w781;
w783 <= w717 and not w782;
w784 <= not a(10) and not w781;
w785 <= a(10) and w781;
w786 <= not w782 and not w785;
w787 <= not w784 and w786;
w788 <= not w783 and not w787;
w789 <= not w706 and not w788;
w790 <= w706 and not w787;
w791 <= not w783 and w790;
w792 <= not w789 and not w791;
w793 <= not w780 and w792;
w794 <= w780 and not w792;
w795 <= not w793 and not w794;
w796 <= not w779 and w795;
w797 <= w779 and not w795;
w798 <= not w796 and not w797;
w799 <= a(15) and a(17);
w800 <= w58 and w799;
w801 <= a(15) and w18;
w802 <= a(17) and w2;
w803 <= not w801 and not w802;
w804 <= a(19) and not w800;
w805 <= not w803 and w804;
w806 <= not w800 and not w805;
w807 <= a(2) and a(17);
w808 <= a(4) and a(15);
w809 <= not w807 and not w808;
w810 <= w806 and not w809;
w811 <= a(19) and not w805;
w812 <= a(0) and w811;
w813 <= not w810 and not w812;
w814 <= w141 and w554;
w815 <= w74 and w412;
w816 <= w138 and w551;
w817 <= not w815 and not w816;
w818 <= not w814 and not w817;
w819 <= a(14) and not w818;
w820 <= a(5) and w819;
w821 <= not w814 and not w818;
w822 <= a(6) and a(13);
w823 <= a(7) and a(12);
w824 <= not w822 and not w823;
w825 <= w821 and not w824;
w826 <= not w820 and not w825;
w827 <= not w813 and not w826;
w828 <= not w813 and not w827;
w829 <= not w826 and not w827;
w830 <= not w828 and not w829;
w831 <= not w740 and not w743;
w832 <= w830 and w831;
w833 <= not w830 and not w831;
w834 <= not w832 and not w833;
w835 <= not w748 and not w750;
w836 <= w834 and not w835;
w837 <= not w834 and w835;
w838 <= not w836 and not w837;
w839 <= w798 and w838;
w840 <= not w798 and not w838;
w841 <= not w839 and not w840;
w842 <= not w735 and not w753;
w843 <= not w841 and w842;
w844 <= w841 and not w842;
w845 <= not w843 and not w844;
w846 <= not w756 and not w760;
w847 <= not w845 and w846;
w848 <= w845 and not w846;
w849 <= not w847 and not w848;
w850 <= not w843 and not w846;
w851 <= not w844 and not w850;
w852 <= not w836 and not w839;
w853 <= not w782 and not w789;
w854 <= a(16) and a(17);
w855 <= w15 and w854;
w856 <= a(16) and a(18);
w857 <= w58 and w856;
w858 <= a(17) and a(18);
w859 <= w24 and w858;
w860 <= not w857 and not w859;
w861 <= not w855 and not w860;
w862 <= a(18) and not w861;
w863 <= a(2) and w862;
w864 <= not w855 and not w861;
w865 <= a(3) and a(17);
w866 <= a(4) and a(16);
w867 <= not w865 and not w866;
w868 <= w864 and not w867;
w869 <= not w863 and not w868;
w870 <= not w853 and not w869;
w871 <= not w853 and not w870;
w872 <= not w869 and not w870;
w873 <= not w871 and not w872;
w874 <= not w764 and not w776;
w875 <= w873 and w874;
w876 <= not w873 and not w874;
w877 <= not w875 and not w876;
w878 <= not w793 and not w796;
w879 <= not w877 and w878;
w880 <= w877 and not w878;
w881 <= not w879 and not w880;
w882 <= a(9) and a(11);
w883 <= a(1) and a(19);
w884 <= not w882 and not w883;
w885 <= w882 and w883;
w886 <= not w773 and not w885;
w887 <= not w884 and w886;
w888 <= not w773 and not w887;
w889 <= not w885 and not w887;
w890 <= not w884 and w889;
w891 <= not w888 and not w890;
w892 <= not w806 and not w891;
w893 <= not w806 and not w892;
w894 <= not w891 and not w892;
w895 <= not w893 and not w894;
w896 <= not w827 and not w833;
w897 <= w895 and w896;
w898 <= not w895 and not w896;
w899 <= not w897 and not w898;
w900 <= a(0) and a(20);
w901 <= a(7) and a(13);
w902 <= not w900 and not w901;
w903 <= w900 and w901;
w904 <= not w902 and not w903;
w905 <= w785 and w904;
w906 <= not w785 and not w904;
w907 <= not w905 and not w906;
w908 <= not w821 and w907;
w909 <= w821 and not w907;
w910 <= not w908 and not w909;
w911 <= w138 and w701;
w912 <= w118 and w412;
w913 <= a(8) and a(15);
w914 <= w598 and w913;
w915 <= not w912 and not w914;
w916 <= not w911 and not w915;
w917 <= a(12) and not w916;
w918 <= a(8) and w917;
w919 <= not w911 and not w916;
w920 <= a(5) and a(15);
w921 <= a(6) and a(14);
w922 <= not w920 and not w921;
w923 <= w919 and not w922;
w924 <= not w918 and not w923;
w925 <= w910 and not w924;
w926 <= w910 and not w925;
w927 <= not w924 and not w925;
w928 <= not w926 and not w927;
w929 <= w899 and not w928;
w930 <= not w899 and w928;
w931 <= w881 and not w930;
w932 <= not w929 and w931;
w933 <= w881 and not w932;
w934 <= not w930 and not w932;
w935 <= not w929 and w934;
w936 <= not w933 and not w935;
w937 <= not w852 and not w936;
w938 <= w852 and w936;
w939 <= not w937 and not w938;
w940 <= not w851 and w939;
w941 <= w851 and not w939;
w942 <= not w940 and not w941;
w943 <= not w880 and not w932;
w944 <= w864 and w919;
w945 <= not w864 and not w919;
w946 <= not w944 and not w945;
w947 <= not w903 and not w905;
w948 <= not w946 and w947;
w949 <= w946 and not w947;
w950 <= not w948 and not w949;
w951 <= not w870 and not w876;
w952 <= not w950 and w951;
w953 <= w950 and not w951;
w954 <= not w952 and not w953;
w955 <= a(18) and a(19);
w956 <= w24 and w955;
w957 <= a(19) and w708;
w958 <= a(3) and w856;
w959 <= not w957 and not w958;
w960 <= a(5) and not w956;
w961 <= not w959 and w960;
w962 <= not w956 and not w961;
w963 <= a(2) and a(19);
w964 <= a(3) and a(18);
w965 <= not w963 and not w964;
w966 <= w962 and not w965;
w967 <= a(16) and not w961;
w968 <= a(5) and w967;
w969 <= not w966 and not w968;
w970 <= w186 and w551;
w971 <= w118 and w627;
w972 <= w141 and w701;
w973 <= not w971 and not w972;
w974 <= not w970 and not w973;
w975 <= a(15) and not w974;
w976 <= a(6) and w975;
w977 <= not w970 and not w974;
w978 <= a(7) and a(14);
w979 <= a(8) and a(13);
w980 <= not w978 and not w979;
w981 <= w977 and not w980;
w982 <= not w976 and not w981;
w983 <= not w969 and not w982;
w984 <= not w969 and not w983;
w985 <= not w982 and not w983;
w986 <= not w984 and not w985;
w987 <= a(4) and a(17);
w988 <= a(9) and a(12);
w989 <= not w529 and not w988;
w990 <= w290 and w408;
w991 <= w987 and not w990;
w992 <= not w989 and w991;
w993 <= w987 and not w992;
w994 <= not w990 and not w992;
w995 <= not w989 and w994;
w996 <= not w993 and not w995;
w997 <= not w986 and not w996;
w998 <= not w986 and not w997;
w999 <= not w996 and not w997;
w1000 <= not w998 and not w999;
w1001 <= not w954 and w1000;
w1002 <= w954 and not w1000;
w1003 <= not w1001 and not w1002;
w1004 <= not w887 and not w892;
w1005 <= a(0) and a(21);
w1006 <= w885 and not w1005;
w1007 <= not w885 and w1005;
w1008 <= not w1006 and not w1007;
w1009 <= a(1) and a(20);
w1010 <= a(11) and w1009;
w1011 <= a(11) and not w1010;
w1012 <= w1009 and not w1010;
w1013 <= not w1011 and not w1012;
w1014 <= not w1008 and not w1013;
w1015 <= w1008 and w1013;
w1016 <= not w1014 and not w1015;
w1017 <= w1004 and not w1016;
w1018 <= not w1004 and w1016;
w1019 <= not w1017 and not w1018;
w1020 <= not w908 and not w925;
w1021 <= not w1019 and w1020;
w1022 <= w1019 and not w1020;
w1023 <= not w1021 and not w1022;
w1024 <= not w898 and not w929;
w1025 <= w1023 and not w1024;
w1026 <= not w1023 and w1024;
w1027 <= not w1025 and not w1026;
w1028 <= w1003 and w1027;
w1029 <= not w1003 and not w1027;
w1030 <= not w1028 and not w1029;
w1031 <= not w943 and w1030;
w1032 <= w943 and not w1030;
w1033 <= not w1031 and not w1032;
w1034 <= not w851 and not w938;
w1035 <= not w937 and not w1034;
w1036 <= not w1033 and w1035;
w1037 <= w1033 and not w1035;
w1038 <= not w1036 and not w1037;
w1039 <= not w1032 and not w1035;
w1040 <= not w1031 and not w1039;
w1041 <= not w1025 and not w1028;
w1042 <= w962 and w977;
w1043 <= not w962 and not w977;
w1044 <= not w1042 and not w1043;
w1045 <= w885 and w1005;
w1046 <= not w1014 and not w1045;
w1047 <= not w1044 and w1046;
w1048 <= w1044 and not w1046;
w1049 <= not w1047 and not w1048;
w1050 <= not w1018 and not w1022;
w1051 <= not w1049 and w1050;
w1052 <= w1049 and not w1050;
w1053 <= not w1051 and not w1052;
w1054 <= a(7) and a(15);
w1055 <= a(8) and a(14);
w1056 <= not w1054 and not w1055;
w1057 <= w186 and w701;
w1058 <= a(0) and not w1057;
w1059 <= a(22) and w1058;
w1060 <= not w1056 and w1059;
w1061 <= not w1057 and not w1060;
w1062 <= not w1056 and w1061;
w1063 <= a(22) and not w1060;
w1064 <= a(0) and w1063;
w1065 <= not w1062 and not w1064;
w1066 <= a(2) and a(20);
w1067 <= not w527 and not w1066;
w1068 <= w527 and w1066;
w1069 <= w332 and not w1068;
w1070 <= not w1067 and w1069;
w1071 <= w332 and not w1070;
w1072 <= not w1068 and not w1070;
w1073 <= not w1067 and w1072;
w1074 <= not w1071 and not w1073;
w1075 <= not w1065 and not w1074;
w1076 <= not w1065 and not w1075;
w1077 <= not w1074 and not w1075;
w1078 <= not w1076 and not w1077;
w1079 <= a(3) and a(19);
w1080 <= w32 and w858;
w1081 <= w15 and w955;
w1082 <= a(5) and a(17);
w1083 <= w1079 and w1082;
w1084 <= not w1081 and not w1083;
w1085 <= not w1080 and not w1084;
w1086 <= w1079 and not w1085;
w1087 <= not w1080 and not w1085;
w1088 <= a(4) and a(18);
w1089 <= not w1082 and not w1088;
w1090 <= w1087 and not w1089;
w1091 <= not w1086 and not w1090;
w1092 <= not w1078 and not w1091;
w1093 <= not w1078 and not w1092;
w1094 <= not w1091 and not w1092;
w1095 <= not w1093 and not w1094;
w1096 <= not w1053 and w1095;
w1097 <= w1053 and not w1095;
w1098 <= not w1096 and not w1097;
w1099 <= not w953 and not w1002;
w1100 <= not w983 and not w997;
w1101 <= not w945 and not w949;
w1102 <= a(1) and a(21);
w1103 <= w286 and w1102;
w1104 <= not w286 and not w1102;
w1105 <= not w1103 and not w1104;
w1106 <= w1010 and w1105;
w1107 <= not w1010 and not w1105;
w1108 <= not w1106 and not w1107;
w1109 <= not w994 and w1108;
w1110 <= w994 and not w1108;
w1111 <= not w1109 and not w1110;
w1112 <= not w1101 and w1111;
w1113 <= not w1101 and not w1112;
w1114 <= w1111 and not w1112;
w1115 <= not w1113 and not w1114;
w1116 <= not w1100 and not w1115;
w1117 <= w1100 and not w1114;
w1118 <= not w1113 and w1117;
w1119 <= not w1116 and not w1118;
w1120 <= not w1099 and w1119;
w1121 <= not w1099 and not w1120;
w1122 <= w1119 and not w1120;
w1123 <= not w1121 and not w1122;
w1124 <= w1098 and not w1123;
w1125 <= not w1098 and not w1122;
w1126 <= not w1121 and w1125;
w1127 <= not w1124 and not w1126;
w1128 <= not w1041 and w1127;
w1129 <= w1041 and not w1127;
w1130 <= not w1128 and not w1129;
w1131 <= w1040 and not w1130;
w1132 <= not w1040 and not w1129;
w1133 <= not w1128 and w1132;
w1134 <= not w1131 and not w1133;
w1135 <= not w1120 and not w1124;
w1136 <= not w1112 and not w1116;
w1137 <= a(18) and a(20);
w1138 <= w106 and w1137;
w1139 <= a(17) and a(20);
w1140 <= w146 and w1139;
w1141 <= w138 and w858;
w1142 <= not w1140 and not w1141;
w1143 <= not w1138 and not w1142;
w1144 <= not w1138 and not w1143;
w1145 <= a(3) and a(20);
w1146 <= a(5) and a(18);
w1147 <= not w1145 and not w1146;
w1148 <= w1144 and not w1147;
w1149 <= a(17) and not w1143;
w1150 <= a(6) and w1149;
w1151 <= not w1148 and not w1150;
w1152 <= a(4) and a(19);
w1153 <= a(10) and a(13);
w1154 <= not w408 and not w1153;
w1155 <= w529 and w554;
w1156 <= w1152 and not w1155;
w1157 <= not w1154 and w1156;
w1158 <= w1152 and not w1157;
w1159 <= not w1155 and not w1157;
w1160 <= not w1154 and w1159;
w1161 <= not w1158 and not w1160;
w1162 <= not w1151 and not w1161;
w1163 <= not w1151 and not w1162;
w1164 <= not w1161 and not w1162;
w1165 <= not w1163 and not w1164;
w1166 <= not w1106 and not w1109;
w1167 <= w1165 and w1166;
w1168 <= not w1165 and not w1166;
w1169 <= not w1167 and not w1168;
w1170 <= a(0) and a(23);
w1171 <= a(2) and a(21);
w1172 <= not w1170 and not w1171;
w1173 <= a(21) and a(23);
w1174 <= w2 and w1173;
w1175 <= not w1172 and not w1174;
w1176 <= w1103 and w1175;
w1177 <= not w1174 and not w1176;
w1178 <= not w1172 and w1177;
w1179 <= w1103 and not w1176;
w1180 <= not w1178 and not w1179;
w1181 <= w1061 and not w1180;
w1182 <= not w1061 and w1180;
w1183 <= not w1181 and not w1182;
w1184 <= w238 and w701;
w1185 <= w569 and w699;
w1186 <= w186 and w697;
w1187 <= not w1185 and not w1186;
w1188 <= not w1184 and not w1187;
w1189 <= a(16) and not w1188;
w1190 <= a(7) and w1189;
w1191 <= a(9) and a(14);
w1192 <= not w913 and not w1191;
w1193 <= not w1184 and not w1188;
w1194 <= not w1192 and w1193;
w1195 <= not w1190 and not w1194;
w1196 <= not w1183 and not w1195;
w1197 <= w1183 and w1195;
w1198 <= not w1196 and not w1197;
w1199 <= not w1169 and not w1198;
w1200 <= w1169 and w1198;
w1201 <= not w1199 and not w1200;
w1202 <= not w1136 and w1201;
w1203 <= w1136 and not w1201;
w1204 <= not w1202 and not w1203;
w1205 <= not w1052 and not w1097;
w1206 <= not w1043 and not w1048;
w1207 <= not w1075 and not w1092;
w1208 <= w1206 and w1207;
w1209 <= not w1206 and not w1207;
w1210 <= not w1208 and not w1209;
w1211 <= a(1) and a(22);
w1212 <= a(12) and w1211;
w1213 <= not a(12) and not w1211;
w1214 <= not w1212 and not w1213;
w1215 <= w1087 and not w1214;
w1216 <= not w1087 and w1214;
w1217 <= not w1215 and not w1216;
w1218 <= not w1072 and w1217;
w1219 <= w1072 and not w1217;
w1220 <= not w1218 and not w1219;
w1221 <= w1210 and w1220;
w1222 <= not w1210 and not w1220;
w1223 <= not w1221 and not w1222;
w1224 <= not w1205 and w1223;
w1225 <= w1205 and not w1223;
w1226 <= not w1224 and not w1225;
w1227 <= w1204 and w1226;
w1228 <= not w1204 and not w1226;
w1229 <= not w1227 and not w1228;
w1230 <= w1135 and not w1229;
w1231 <= not w1135 and w1229;
w1232 <= not w1230 and not w1231;
w1233 <= not w1128 and not w1132;
w1234 <= not w1232 and w1233;
w1235 <= w1232 and not w1233;
w1236 <= not w1234 and not w1235;
w1237 <= not w1230 and not w1233;
w1238 <= not w1231 and not w1237;
w1239 <= not w1224 and not w1227;
w1240 <= not w1200 and not w1202;
w1241 <= w1144 and w1159;
w1242 <= not w1144 and not w1159;
w1243 <= not w1241 and not w1242;
w1244 <= w1193 and not w1243;
w1245 <= not w1193 and w1243;
w1246 <= not w1244 and not w1245;
w1247 <= not w1162 and not w1168;
w1248 <= not w1061 and not w1180;
w1249 <= not w1196 and not w1248;
w1250 <= w1247 and w1249;
w1251 <= not w1247 and not w1249;
w1252 <= not w1250 and not w1251;
w1253 <= w1246 and w1252;
w1254 <= not w1246 and not w1252;
w1255 <= not w1253 and not w1254;
w1256 <= not w1240 and w1255;
w1257 <= not w1240 and not w1256;
w1258 <= w1255 and not w1256;
w1259 <= not w1257 and not w1258;
w1260 <= a(0) and a(24);
w1261 <= w1212 and w1260;
w1262 <= w1212 and not w1261;
w1263 <= not w1212 and w1260;
w1264 <= not w1262 and not w1263;
w1265 <= a(1) and a(23);
w1266 <= w624 and w1265;
w1267 <= w1265 and not w1266;
w1268 <= w624 and not w1266;
w1269 <= not w1267 and not w1268;
w1270 <= not w1264 and not w1269;
w1271 <= not w1264 and not w1270;
w1272 <= not w1269 and not w1270;
w1273 <= not w1271 and not w1272;
w1274 <= a(7) and a(17);
w1275 <= a(18) and a(22);
w1276 <= w116 and w1275;
w1277 <= w141 and w858;
w1278 <= a(2) and a(22);
w1279 <= w1274 and w1278;
w1280 <= not w1277 and not w1279;
w1281 <= not w1276 and not w1280;
w1282 <= w1274 and not w1281;
w1283 <= not w1276 and not w1281;
w1284 <= a(6) and a(18);
w1285 <= not w1278 and not w1284;
w1286 <= w1283 and not w1285;
w1287 <= not w1282 and not w1286;
w1288 <= not w1273 and not w1287;
w1289 <= not w1273 and not w1288;
w1290 <= not w1287 and not w1288;
w1291 <= not w1289 and not w1290;
w1292 <= not w1216 and not w1218;
w1293 <= w1291 and w1292;
w1294 <= not w1291 and not w1292;
w1295 <= not w1293 and not w1294;
w1296 <= a(19) and a(20);
w1297 <= w32 and w1296;
w1298 <= a(19) and a(21);
w1299 <= w106 and w1298;
w1300 <= a(20) and a(21);
w1301 <= w15 and w1300;
w1302 <= not w1299 and not w1301;
w1303 <= not w1297 and not w1302;
w1304 <= a(3) and not w1303;
w1305 <= a(21) and w1304;
w1306 <= not w1297 and not w1303;
w1307 <= a(4) and a(20);
w1308 <= a(5) and a(19);
w1309 <= not w1307 and not w1308;
w1310 <= w1306 and not w1309;
w1311 <= not w1305 and not w1310;
w1312 <= w1177 and not w1311;
w1313 <= not w1177 and w1311;
w1314 <= not w1312 and not w1313;
w1315 <= a(8) and a(16);
w1316 <= w290 and w701;
w1317 <= w184 and w699;
w1318 <= w238 and w697;
w1319 <= not w1317 and not w1318;
w1320 <= not w1316 and not w1319;
w1321 <= w1315 and not w1320;
w1322 <= not w1316 and not w1320;
w1323 <= a(9) and a(15);
w1324 <= a(10) and a(14);
w1325 <= not w1323 and not w1324;
w1326 <= w1322 and not w1325;
w1327 <= not w1321 and not w1326;
w1328 <= not w1314 and not w1327;
w1329 <= w1314 and w1327;
w1330 <= not w1328 and not w1329;
w1331 <= not w1295 and not w1330;
w1332 <= w1295 and w1330;
w1333 <= not w1331 and not w1332;
w1334 <= not w1209 and not w1221;
w1335 <= w1333 and not w1334;
w1336 <= not w1333 and w1334;
w1337 <= not w1335 and not w1336;
w1338 <= not w1259 and w1337;
w1339 <= not w1258 and not w1337;
w1340 <= not w1257 and w1339;
w1341 <= not w1338 and not w1340;
w1342 <= not w1239 and w1341;
w1343 <= w1239 and not w1341;
w1344 <= not w1342 and not w1343;
w1345 <= w1238 and not w1344;
w1346 <= not w1238 and not w1343;
w1347 <= not w1342 and w1346;
w1348 <= not w1345 and not w1347;
w1349 <= not w1256 and not w1338;
w1350 <= a(0) and a(25);
w1351 <= a(2) and a(23);
w1352 <= not w1350 and not w1351;
w1353 <= a(23) and a(25);
w1354 <= w2 and w1353;
w1355 <= w491 and not w1354;
w1356 <= not w1352 and w1355;
w1357 <= not w1354 and not w1356;
w1358 <= not w1352 and w1357;
w1359 <= w491 and not w1356;
w1360 <= not w1358 and not w1359;
w1361 <= w238 and w854;
w1362 <= w569 and w856;
w1363 <= w186 and w858;
w1364 <= not w1362 and not w1363;
w1365 <= not w1361 and not w1364;
w1366 <= w682 and not w1365;
w1367 <= not w1361 and not w1365;
w1368 <= a(8) and a(17);
w1369 <= not w653 and not w1368;
w1370 <= w1367 and not w1369;
w1371 <= not w1366 and not w1370;
w1372 <= not w1360 and not w1371;
w1373 <= not w1360 and not w1372;
w1374 <= not w1371 and not w1372;
w1375 <= not w1373 and not w1374;
w1376 <= a(6) and a(19);
w1377 <= a(22) and w1079;
w1378 <= a(4) and w1298;
w1379 <= not w1377 and not w1378;
w1380 <= a(21) and a(22);
w1381 <= w15 and w1380;
w1382 <= a(6) and not w1381;
w1383 <= not w1379 and w1382;
w1384 <= w1376 and not w1383;
w1385 <= not w1381 and not w1383;
w1386 <= a(3) and a(22);
w1387 <= a(4) and a(21);
w1388 <= not w1386 and not w1387;
w1389 <= w1385 and not w1388;
w1390 <= not w1384 and not w1389;
w1391 <= not w1375 and not w1390;
w1392 <= not w1375 and not w1391;
w1393 <= not w1390 and not w1391;
w1394 <= not w1392 and not w1393;
w1395 <= not w1251 and not w1253;
w1396 <= not w1394 and not w1395;
w1397 <= not w1394 and not w1396;
w1398 <= not w1395 and not w1396;
w1399 <= not w1397 and not w1398;
w1400 <= a(1) and a(24);
w1401 <= a(13) and w1400;
w1402 <= not a(13) and not w1400;
w1403 <= not w1401 and not w1402;
w1404 <= w1266 and w1403;
w1405 <= not w1266 and not w1403;
w1406 <= not w1404 and not w1405;
w1407 <= not w1306 and w1406;
w1408 <= w1306 and not w1406;
w1409 <= not w1407 and not w1408;
w1410 <= not w1242 and not w1245;
w1411 <= a(11) and a(14);
w1412 <= not w554 and not w1411;
w1413 <= w554 and w1411;
w1414 <= a(5) and not w1413;
w1415 <= a(20) and w1414;
w1416 <= not w1412 and w1415;
w1417 <= a(5) and not w1416;
w1418 <= a(20) and w1417;
w1419 <= not w1413 and not w1416;
w1420 <= not w1412 and w1419;
w1421 <= not w1418 and not w1420;
w1422 <= not w1410 and not w1421;
w1423 <= not w1410 and not w1422;
w1424 <= not w1421 and not w1422;
w1425 <= not w1423 and not w1424;
w1426 <= w1409 and not w1425;
w1427 <= w1409 and not w1426;
w1428 <= not w1425 and not w1426;
w1429 <= not w1427 and not w1428;
w1430 <= not w1399 and not w1429;
w1431 <= not w1399 and not w1430;
w1432 <= not w1429 and not w1430;
w1433 <= not w1431 and not w1432;
w1434 <= w1283 and w1322;
w1435 <= not w1283 and not w1322;
w1436 <= not w1434 and not w1435;
w1437 <= not w1261 and not w1270;
w1438 <= not w1436 and w1437;
w1439 <= w1436 and not w1437;
w1440 <= not w1438 and not w1439;
w1441 <= not w1177 and not w1311;
w1442 <= not w1328 and not w1441;
w1443 <= not w1440 and w1442;
w1444 <= w1440 and not w1442;
w1445 <= not w1443 and not w1444;
w1446 <= not w1288 and not w1294;
w1447 <= not w1445 and w1446;
w1448 <= w1445 and not w1446;
w1449 <= not w1447 and not w1448;
w1450 <= not w1332 and not w1335;
w1451 <= w1449 and not w1450;
w1452 <= w1449 and not w1451;
w1453 <= not w1450 and not w1451;
w1454 <= not w1452 and not w1453;
w1455 <= not w1433 and not w1454;
w1456 <= w1433 and not w1453;
w1457 <= not w1452 and w1456;
w1458 <= not w1455 and not w1457;
w1459 <= w1349 and not w1458;
w1460 <= not w1349 and w1458;
w1461 <= not w1459 and not w1460;
w1462 <= not w1342 and not w1346;
w1463 <= not w1461 and w1462;
w1464 <= w1461 and not w1462;
w1465 <= not w1463 and not w1464;
w1466 <= not w1451 and not w1455;
w1467 <= a(3) and a(23);
w1468 <= a(7) and a(19);
w1469 <= not w1467 and not w1468;
w1470 <= a(19) and a(24);
w1471 <= w149 and w1470;
w1472 <= a(23) and a(24);
w1473 <= w24 and w1472;
w1474 <= not w1471 and not w1473;
w1475 <= w1467 and w1468;
w1476 <= not w1474 and not w1475;
w1477 <= not w1475 and not w1476;
w1478 <= not w1469 and w1477;
w1479 <= a(24) and not w1476;
w1480 <= a(2) and w1479;
w1481 <= not w1478 and not w1480;
w1482 <= a(9) and a(17);
w1483 <= w529 and w697;
w1484 <= w622 and w1482;
w1485 <= w290 and w854;
w1486 <= not w1484 and not w1485;
w1487 <= not w1483 and not w1486;
w1488 <= w1482 and not w1487;
w1489 <= not w1483 and not w1487;
w1490 <= a(10) and a(16);
w1491 <= not w622 and not w1490;
w1492 <= w1489 and not w1491;
w1493 <= not w1488 and not w1492;
w1494 <= not w1481 and not w1493;
w1495 <= not w1481 and not w1494;
w1496 <= not w1493 and not w1494;
w1497 <= not w1495 and not w1496;
w1498 <= w138 and w1300;
w1499 <= a(20) and a(22);
w1500 <= w206 and w1499;
w1501 <= w32 and w1380;
w1502 <= not w1500 and not w1501;
w1503 <= not w1498 and not w1502;
w1504 <= a(22) and not w1503;
w1505 <= a(4) and w1504;
w1506 <= not w1498 and not w1503;
w1507 <= a(5) and a(21);
w1508 <= a(6) and a(20);
w1509 <= not w1507 and not w1508;
w1510 <= w1506 and not w1509;
w1511 <= not w1505 and not w1510;
w1512 <= not w1497 and not w1511;
w1513 <= not w1497 and not w1512;
w1514 <= not w1511 and not w1512;
w1515 <= not w1513 and not w1514;
w1516 <= not w1444 and not w1448;
w1517 <= w1515 and w1516;
w1518 <= not w1515 and not w1516;
w1519 <= not w1517 and not w1518;
w1520 <= not w1435 and not w1439;
w1521 <= not w1404 and not w1407;
w1522 <= w1520 and w1521;
w1523 <= not w1520 and not w1521;
w1524 <= not w1522 and not w1523;
w1525 <= w1357 and w1367;
w1526 <= not w1357 and not w1367;
w1527 <= not w1525 and not w1526;
w1528 <= a(0) and a(26);
w1529 <= a(8) and a(18);
w1530 <= not w1528 and not w1529;
w1531 <= w1528 and w1529;
w1532 <= not w1530 and not w1531;
w1533 <= w1401 and w1532;
w1534 <= w1401 and not w1533;
w1535 <= not w1531 and not w1533;
w1536 <= not w1530 and w1535;
w1537 <= not w1534 and not w1536;
w1538 <= w1527 and not w1537;
w1539 <= w1527 and not w1538;
w1540 <= not w1537 and not w1538;
w1541 <= not w1539 and not w1540;
w1542 <= w1524 and not w1541;
w1543 <= not w1524 and w1541;
w1544 <= w1519 and not w1543;
w1545 <= not w1542 and w1544;
w1546 <= w1519 and not w1545;
w1547 <= not w1543 and not w1545;
w1548 <= not w1542 and w1547;
w1549 <= not w1546 and not w1548;
w1550 <= not w1396 and not w1430;
w1551 <= not w1422 and not w1426;
w1552 <= not w1372 and not w1391;
w1553 <= a(1) and a(25);
w1554 <= not w412 and not w1553;
w1555 <= w412 and w1553;
w1556 <= not w1419 and not w1555;
w1557 <= not w1554 and w1556;
w1558 <= not w1419 and not w1557;
w1559 <= not w1555 and not w1557;
w1560 <= not w1554 and w1559;
w1561 <= not w1558 and not w1560;
w1562 <= not w1385 and not w1561;
w1563 <= w1385 and not w1560;
w1564 <= not w1558 and w1563;
w1565 <= not w1562 and not w1564;
w1566 <= not w1552 and w1565;
w1567 <= w1552 and not w1565;
w1568 <= not w1566 and not w1567;
w1569 <= not w1551 and w1568;
w1570 <= w1551 and not w1568;
w1571 <= not w1569 and not w1570;
w1572 <= not w1550 and w1571;
w1573 <= w1550 and not w1571;
w1574 <= not w1572 and not w1573;
w1575 <= not w1549 and not w1574;
w1576 <= w1549 and w1574;
w1577 <= not w1575 and not w1576;
w1578 <= not w1466 and not w1577;
w1579 <= w1466 and w1577;
w1580 <= not w1578 and not w1579;
w1581 <= not w1459 and not w1462;
w1582 <= not w1460 and not w1581;
w1583 <= not w1580 and w1582;
w1584 <= w1580 and not w1582;
w1585 <= not w1583 and not w1584;
w1586 <= not w1549 and w1574;
w1587 <= not w1572 and not w1586;
w1588 <= not w1518 and not w1545;
w1589 <= a(21) and a(24);
w1590 <= w146 and w1589;
w1591 <= w15 and w1472;
w1592 <= not w1590 and not w1591;
w1593 <= a(4) and a(23);
w1594 <= a(6) and a(21);
w1595 <= w1593 and w1594;
w1596 <= not w1592 and not w1595;
w1597 <= not w1595 and not w1596;
w1598 <= not w1593 and not w1594;
w1599 <= w1597 and not w1598;
w1600 <= a(24) and not w1596;
w1601 <= a(3) and w1600;
w1602 <= not w1599 and not w1601;
w1603 <= a(12) and a(15);
w1604 <= not w551 and not w1603;
w1605 <= w554 and w701;
w1606 <= a(5) and not w1605;
w1607 <= a(22) and w1606;
w1608 <= not w1604 and w1607;
w1609 <= a(22) and not w1608;
w1610 <= a(5) and w1609;
w1611 <= not w1605 and not w1608;
w1612 <= not w1604 and w1611;
w1613 <= not w1610 and not w1612;
w1614 <= not w1602 and not w1613;
w1615 <= not w1602 and not w1614;
w1616 <= not w1613 and not w1614;
w1617 <= not w1615 and not w1616;
w1618 <= a(0) and a(27);
w1619 <= w1555 and not w1618;
w1620 <= not w1555 and w1618;
w1621 <= not w1619 and not w1620;
w1622 <= a(26) and w458;
w1623 <= a(14) and not w1622;
w1624 <= a(1) and not w1622;
w1625 <= a(26) and w1624;
w1626 <= not w1623 and not w1625;
w1627 <= not w1621 and not w1626;
w1628 <= w1621 and w1626;
w1629 <= not w1627 and not w1628;
w1630 <= w1617 and w1629;
w1631 <= not w1617 and not w1629;
w1632 <= not w1630 and not w1631;
w1633 <= w1489 and w1506;
w1634 <= not w1489 and not w1506;
w1635 <= not w1633 and not w1634;
w1636 <= w1477 and not w1635;
w1637 <= not w1477 and w1635;
w1638 <= not w1636 and not w1637;
w1639 <= not w1523 and not w1542;
w1640 <= w1638 and not w1639;
w1641 <= not w1638 and w1639;
w1642 <= not w1640 and not w1641;
w1643 <= not w1632 and w1642;
w1644 <= w1632 and not w1642;
w1645 <= not w1643 and not w1644;
w1646 <= not w1588 and w1645;
w1647 <= w1588 and not w1645;
w1648 <= not w1646 and not w1647;
w1649 <= a(11) and a(16);
w1650 <= a(20) and a(25);
w1651 <= w149 and w1650;
w1652 <= a(2) and a(25);
w1653 <= a(7) and a(20);
w1654 <= not w1652 and not w1653;
w1655 <= not w1651 and not w1654;
w1656 <= not w1649 and not w1655;
w1657 <= w1649 and w1655;
w1658 <= not w1656 and not w1657;
w1659 <= not w1535 and w1658;
w1660 <= w1535 and not w1658;
w1661 <= not w1659 and not w1660;
w1662 <= a(8) and a(19);
w1663 <= w290 and w858;
w1664 <= a(10) and a(17);
w1665 <= w1662 and w1664;
w1666 <= w238 and w955;
w1667 <= not w1665 and not w1666;
w1668 <= not w1663 and not w1667;
w1669 <= w1662 and not w1668;
w1670 <= not w1663 and not w1668;
w1671 <= a(9) and a(18);
w1672 <= not w1664 and not w1671;
w1673 <= w1670 and not w1672;
w1674 <= not w1669 and not w1673;
w1675 <= w1661 and not w1674;
w1676 <= w1661 and not w1675;
w1677 <= not w1674 and not w1675;
w1678 <= not w1676 and not w1677;
w1679 <= not w1566 and not w1569;
w1680 <= w1678 and w1679;
w1681 <= not w1678 and not w1679;
w1682 <= not w1680 and not w1681;
w1683 <= not w1557 and not w1562;
w1684 <= not w1526 and not w1538;
w1685 <= w1683 and w1684;
w1686 <= not w1683 and not w1684;
w1687 <= not w1685 and not w1686;
w1688 <= not w1494 and not w1512;
w1689 <= not w1687 and w1688;
w1690 <= w1687 and not w1688;
w1691 <= not w1689 and not w1690;
w1692 <= w1682 and w1691;
w1693 <= not w1682 and not w1691;
w1694 <= not w1692 and not w1693;
w1695 <= w1648 and w1694;
w1696 <= not w1648 and not w1694;
w1697 <= not w1695 and not w1696;
w1698 <= not w1587 and w1697;
w1699 <= w1587 and not w1697;
w1700 <= not w1698 and not w1699;
w1701 <= not w1579 and not w1582;
w1702 <= not w1578 and not w1701;
w1703 <= not w1700 and w1702;
w1704 <= w1700 and not w1702;
w1705 <= not w1703 and not w1704;
w1706 <= not w1640 and not w1643;
w1707 <= a(3) and a(25);
w1708 <= a(4) and a(24);
w1709 <= not w1707 and not w1708;
w1710 <= a(24) and a(25);
w1711 <= w15 and w1710;
w1712 <= a(8) and not w1711;
w1713 <= a(20) and w1712;
w1714 <= not w1709 and w1713;
w1715 <= a(8) and not w1714;
w1716 <= a(20) and w1715;
w1717 <= not w1711 and not w1714;
w1718 <= not w1709 and w1717;
w1719 <= not w1716 and not w1718;
w1720 <= w1555 and w1618;
w1721 <= not w1627 and not w1720;
w1722 <= not w1719 and w1721;
w1723 <= w1719 and not w1721;
w1724 <= not w1722 and not w1723;
w1725 <= a(22) and a(23);
w1726 <= w138 and w1725;
w1727 <= w74 and w1173;
w1728 <= w141 and w1380;
w1729 <= not w1727 and not w1728;
w1730 <= not w1726 and not w1729;
w1731 <= a(21) and not w1730;
w1732 <= a(7) and w1731;
w1733 <= not w1726 and not w1730;
w1734 <= a(5) and a(23);
w1735 <= a(6) and a(22);
w1736 <= not w1734 and not w1735;
w1737 <= w1733 and not w1736;
w1738 <= not w1732 and not w1737;
w1739 <= not w1724 and not w1738;
w1740 <= w1724 and w1738;
w1741 <= not w1739 and not w1740;
w1742 <= w1706 and not w1741;
w1743 <= not w1706 and w1741;
w1744 <= not w1742 and not w1743;
w1745 <= not w1617 and w1629;
w1746 <= not w1614 and not w1745;
w1747 <= not w1659 and not w1675;
w1748 <= a(1) and a(27);
w1749 <= w627 and w1748;
w1750 <= not w627 and not w1748;
w1751 <= not w1749 and not w1750;
w1752 <= w1622 and w1751;
w1753 <= w1622 and not w1752;
w1754 <= not w1622 and w1751;
w1755 <= not w1753 and not w1754;
w1756 <= not w1611 and not w1755;
w1757 <= w1611 and not w1754;
w1758 <= not w1753 and w1757;
w1759 <= not w1756 and not w1758;
w1760 <= not w1747 and w1759;
w1761 <= w1747 and not w1759;
w1762 <= not w1760 and not w1761;
w1763 <= not w1746 and w1762;
w1764 <= w1746 and not w1762;
w1765 <= not w1763 and not w1764;
w1766 <= w1744 and w1765;
w1767 <= not w1744 and not w1765;
w1768 <= not w1766 and not w1767;
w1769 <= not w1646 and not w1695;
w1770 <= not w1681 and not w1692;
w1771 <= w1597 and w1670;
w1772 <= not w1597 and not w1670;
w1773 <= not w1771 and not w1772;
w1774 <= not w1651 and not w1657;
w1775 <= not w1773 and w1774;
w1776 <= w1773 and not w1774;
w1777 <= not w1775 and not w1776;
w1778 <= not w1686 and not w1690;
w1779 <= not w1777 and w1778;
w1780 <= w1777 and not w1778;
w1781 <= not w1779 and not w1780;
w1782 <= a(11) and a(28);
w1783 <= w599 and w1782;
w1784 <= w408 and w854;
w1785 <= not w1783 and not w1784;
w1786 <= a(0) and a(28);
w1787 <= a(12) and a(16);
w1788 <= w1786 and w1787;
w1789 <= not w1785 and not w1788;
w1790 <= not w1788 and not w1789;
w1791 <= not w1786 and not w1787;
w1792 <= w1790 and not w1791;
w1793 <= a(17) and not w1789;
w1794 <= a(11) and w1793;
w1795 <= not w1792 and not w1794;
w1796 <= a(2) and a(26);
w1797 <= a(9) and a(19);
w1798 <= a(10) and a(18);
w1799 <= not w1797 and not w1798;
w1800 <= w290 and w955;
w1801 <= w1796 and not w1800;
w1802 <= not w1799 and w1801;
w1803 <= w1796 and not w1802;
w1804 <= not w1800 and not w1802;
w1805 <= not w1799 and w1804;
w1806 <= not w1803 and not w1805;
w1807 <= not w1795 and not w1806;
w1808 <= not w1795 and not w1807;
w1809 <= not w1806 and not w1807;
w1810 <= not w1808 and not w1809;
w1811 <= not w1634 and not w1637;
w1812 <= w1810 and w1811;
w1813 <= not w1810 and not w1811;
w1814 <= not w1812 and not w1813;
w1815 <= w1781 and w1814;
w1816 <= not w1781 and not w1814;
w1817 <= not w1815 and not w1816;
w1818 <= not w1770 and w1817;
w1819 <= w1770 and not w1817;
w1820 <= not w1818 and not w1819;
w1821 <= not w1769 and w1820;
w1822 <= w1769 and not w1820;
w1823 <= not w1821 and not w1822;
w1824 <= not w1768 and not w1823;
w1825 <= w1768 and w1823;
w1826 <= not w1824 and not w1825;
w1827 <= not w1699 and not w1702;
w1828 <= not w1698 and not w1827;
w1829 <= not w1826 and w1828;
w1830 <= w1826 and not w1828;
w1831 <= not w1829 and not w1830;
w1832 <= not w1818 and not w1821;
w1833 <= not w1780 and not w1815;
w1834 <= not w1760 and not w1763;
w1835 <= w1833 and w1834;
w1836 <= not w1833 and not w1834;
w1837 <= not w1835 and not w1836;
w1838 <= not w1807 and not w1813;
w1839 <= not w1719 and not w1721;
w1840 <= not w1739 and not w1839;
w1841 <= w1838 and w1840;
w1842 <= not w1838 and not w1840;
w1843 <= not w1841 and not w1842;
w1844 <= w1790 and w1804;
w1845 <= not w1790 and not w1804;
w1846 <= not w1844 and not w1845;
w1847 <= a(27) and a(29);
w1848 <= w2 and w1847;
w1849 <= a(0) and a(29);
w1850 <= a(2) and a(27);
w1851 <= not w1849 and not w1850;
w1852 <= not w1848 and not w1851;
w1853 <= w1749 and w1852;
w1854 <= w1749 and not w1853;
w1855 <= not w1848 and not w1853;
w1856 <= not w1851 and w1855;
w1857 <= not w1854 and not w1856;
w1858 <= w1846 and not w1857;
w1859 <= w1846 and not w1858;
w1860 <= not w1857 and not w1858;
w1861 <= not w1859 and not w1860;
w1862 <= w1843 and not w1861;
w1863 <= not w1843 and w1861;
w1864 <= w1837 and not w1863;
w1865 <= not w1862 and w1864;
w1866 <= w1837 and not w1865;
w1867 <= not w1863 and not w1865;
w1868 <= not w1862 and w1867;
w1869 <= not w1866 and not w1868;
w1870 <= not w1743 and not w1766;
w1871 <= not w1752 and not w1756;
w1872 <= a(6) and a(23);
w1873 <= a(13) and a(16);
w1874 <= not w701 and not w1873;
w1875 <= w701 and w1873;
w1876 <= w1872 and not w1875;
w1877 <= not w1874 and w1876;
w1878 <= w1872 and not w1877;
w1879 <= not w1875 and not w1877;
w1880 <= not w1874 and w1879;
w1881 <= not w1878 and not w1880;
w1882 <= not w1871 and not w1881;
w1883 <= not w1871 and not w1882;
w1884 <= not w1881 and not w1882;
w1885 <= not w1883 and not w1884;
w1886 <= not w1772 and not w1776;
w1887 <= w1885 and w1886;
w1888 <= not w1885 and not w1886;
w1889 <= not w1887 and not w1888;
w1890 <= a(3) and a(26);
w1891 <= a(8) and a(21);
w1892 <= not w1890 and not w1891;
w1893 <= a(21) and a(26);
w1894 <= w241 and w1893;
w1895 <= a(17) and not w1894;
w1896 <= a(12) and w1895;
w1897 <= not w1892 and w1896;
w1898 <= not w1894 and not w1897;
w1899 <= not w1892 and w1898;
w1900 <= a(17) and not w1897;
w1901 <= a(12) and w1900;
w1902 <= not w1899 and not w1901;
w1903 <= w529 and w955;
w1904 <= w882 and w1137;
w1905 <= w290 and w1296;
w1906 <= not w1904 and not w1905;
w1907 <= not w1903 and not w1906;
w1908 <= a(20) and not w1907;
w1909 <= a(9) and w1908;
w1910 <= not w1903 and not w1907;
w1911 <= a(10) and a(19);
w1912 <= a(11) and a(18);
w1913 <= not w1911 and not w1912;
w1914 <= w1910 and not w1913;
w1915 <= not w1909 and not w1914;
w1916 <= not w1902 and not w1915;
w1917 <= not w1902 and not w1916;
w1918 <= not w1915 and not w1916;
w1919 <= not w1917 and not w1918;
w1920 <= a(4) and a(25);
w1921 <= a(22) and a(24);
w1922 <= w74 and w1921;
w1923 <= w32 and w1710;
w1924 <= a(7) and a(22);
w1925 <= w1920 and w1924;
w1926 <= not w1923 and not w1925;
w1927 <= not w1922 and not w1926;
w1928 <= w1920 and not w1927;
w1929 <= not w1922 and not w1927;
w1930 <= a(5) and a(24);
w1931 <= not w1924 and not w1930;
w1932 <= w1929 and not w1931;
w1933 <= not w1928 and not w1932;
w1934 <= not w1919 and not w1933;
w1935 <= not w1919 and not w1934;
w1936 <= not w1933 and not w1934;
w1937 <= not w1935 and not w1936;
w1938 <= a(28) and w570;
w1939 <= a(1) and a(28);
w1940 <= not a(15) and not w1939;
w1941 <= not w1938 and not w1940;
w1942 <= w1733 and not w1941;
w1943 <= not w1733 and w1941;
w1944 <= not w1942 and not w1943;
w1945 <= not w1717 and w1944;
w1946 <= w1717 and not w1944;
w1947 <= not w1945 and not w1946;
w1948 <= not w1937 and w1947;
w1949 <= w1937 and not w1947;
w1950 <= not w1948 and not w1949;
w1951 <= w1889 and w1950;
w1952 <= not w1889 and not w1950;
w1953 <= not w1951 and not w1952;
w1954 <= not w1870 and w1953;
w1955 <= not w1870 and not w1954;
w1956 <= w1953 and not w1954;
w1957 <= not w1955 and not w1956;
w1958 <= not w1869 and not w1957;
w1959 <= w1869 and not w1956;
w1960 <= not w1955 and w1959;
w1961 <= not w1958 and not w1960;
w1962 <= not w1832 and w1961;
w1963 <= w1832 and not w1961;
w1964 <= not w1962 and not w1963;
w1965 <= not w1824 and not w1828;
w1966 <= not w1825 and not w1965;
w1967 <= not w1964 and w1966;
w1968 <= w1964 and not w1966;
w1969 <= not w1967 and not w1968;
w1970 <= not w1954 and not w1958;
w1971 <= a(0) and a(30);
w1972 <= w1938 and w1971;
w1973 <= w1938 and not w1972;
w1974 <= not w1938 and w1971;
w1975 <= not w1973 and not w1974;
w1976 <= a(1) and a(29);
w1977 <= w699 and w1976;
w1978 <= w1976 and not w1977;
w1979 <= w699 and not w1977;
w1980 <= not w1978 and not w1979;
w1981 <= not w1975 and not w1980;
w1982 <= not w1975 and not w1981;
w1983 <= not w1980 and not w1981;
w1984 <= not w1982 and not w1983;
w1985 <= not w1943 and not w1945;
w1986 <= w1984 and w1985;
w1987 <= not w1984 and not w1985;
w1988 <= not w1986 and not w1987;
w1989 <= not w1845 and not w1858;
w1990 <= not w1988 and w1989;
w1991 <= w1988 and not w1989;
w1992 <= not w1990 and not w1991;
w1993 <= not w1948 and not w1951;
w1994 <= not w1992 and w1993;
w1995 <= w1992 and not w1993;
w1996 <= not w1994 and not w1995;
w1997 <= w1879 and w1929;
w1998 <= not w1879 and not w1929;
w1999 <= not w1997 and not w1998;
w2000 <= a(2) and a(28);
w2001 <= a(9) and a(21);
w2002 <= not w2000 and not w2001;
w2003 <= w2000 and w2001;
w2004 <= a(17) and not w2003;
w2005 <= a(13) and w2004;
w2006 <= not w2002 and w2005;
w2007 <= a(17) and not w2006;
w2008 <= a(13) and w2007;
w2009 <= not w2003 and not w2006;
w2010 <= not w2002 and w2009;
w2011 <= not w2008 and not w2010;
w2012 <= w1999 and not w2011;
w2013 <= w1999 and not w2012;
w2014 <= not w2011 and not w2012;
w2015 <= not w2013 and not w2014;
w2016 <= not w1916 and not w1934;
w2017 <= w2015 and w2016;
w2018 <= not w2015 and not w2016;
w2019 <= not w2017 and not w2018;
w2020 <= w1898 and w1910;
w2021 <= not w1898 and not w1910;
w2022 <= not w2020 and not w2021;
w2023 <= w1855 and not w2022;
w2024 <= not w1855 and w2022;
w2025 <= not w2023 and not w2024;
w2026 <= w2019 and w2025;
w2027 <= not w2019 and not w2025;
w2028 <= not w2026 and not w2027;
w2029 <= w1996 and w2028;
w2030 <= not w1996 and not w2028;
w2031 <= not w2029 and not w2030;
w2032 <= not w1836 and not w1865;
w2033 <= a(26) and a(27);
w2034 <= w15 and w2033;
w2035 <= a(8) and a(27);
w2036 <= w1386 and w2035;
w2037 <= not w2034 and not w2036;
w2038 <= a(4) and a(26);
w2039 <= a(8) and a(22);
w2040 <= w2038 and w2039;
w2041 <= not w2037 and not w2040;
w2042 <= not w2040 and not w2041;
w2043 <= not w2038 and not w2039;
w2044 <= w2042 and not w2043;
w2045 <= a(27) and not w2041;
w2046 <= a(3) and w2045;
w2047 <= not w2044 and not w2046;
w2048 <= w141 and w1472;
w2049 <= w74 and w1353;
w2050 <= w138 and w1710;
w2051 <= not w2049 and not w2050;
w2052 <= not w2048 and not w2051;
w2053 <= a(25) and not w2052;
w2054 <= a(5) and w2053;
w2055 <= not w2048 and not w2052;
w2056 <= a(6) and a(24);
w2057 <= a(7) and a(23);
w2058 <= not w2056 and not w2057;
w2059 <= w2055 and not w2058;
w2060 <= not w2054 and not w2059;
w2061 <= not w2047 and not w2060;
w2062 <= not w2047 and not w2061;
w2063 <= not w2060 and not w2061;
w2064 <= not w2062 and not w2063;
w2065 <= w408 and w955;
w2066 <= w286 and w1137;
w2067 <= w529 and w1296;
w2068 <= not w2066 and not w2067;
w2069 <= not w2065 and not w2068;
w2070 <= a(20) and not w2069;
w2071 <= a(10) and w2070;
w2072 <= a(11) and a(19);
w2073 <= a(12) and a(18);
w2074 <= not w2072 and not w2073;
w2075 <= not w2065 and not w2069;
w2076 <= not w2074 and w2075;
w2077 <= not w2071 and not w2076;
w2078 <= not w2064 and not w2077;
w2079 <= not w2064 and not w2078;
w2080 <= not w2077 and not w2078;
w2081 <= not w2079 and not w2080;
w2082 <= not w1882 and not w1888;
w2083 <= w2081 and w2082;
w2084 <= not w2081 and not w2082;
w2085 <= not w2083 and not w2084;
w2086 <= not w1842 and not w1862;
w2087 <= w2085 and not w2086;
w2088 <= not w2085 and w2086;
w2089 <= not w2087 and not w2088;
w2090 <= not w2032 and w2089;
w2091 <= w2032 and not w2089;
w2092 <= not w2090 and not w2091;
w2093 <= w2031 and w2092;
w2094 <= not w2031 and not w2092;
w2095 <= not w2093 and not w2094;
w2096 <= not w1970 and w2095;
w2097 <= w1970 and not w2095;
w2098 <= not w2096 and not w2097;
w2099 <= not w1963 and not w1966;
w2100 <= not w1962 and not w2099;
w2101 <= not w2098 and w2100;
w2102 <= w2098 and not w2100;
w2103 <= not w2101 and not w2102;
w2104 <= not w2090 and not w2093;
w2105 <= not w1995 and not w2029;
w2106 <= not w2018 and not w2026;
w2107 <= a(24) and a(26);
w2108 <= w74 and w2107;
w2109 <= a(23) and a(26);
w2110 <= w160 and w2109;
w2111 <= w186 and w1472;
w2112 <= not w2110 and not w2111;
w2113 <= not w2108 and not w2112;
w2114 <= not w2108 and not w2113;
w2115 <= a(5) and a(26);
w2116 <= a(7) and a(24);
w2117 <= not w2115 and not w2116;
w2118 <= w2114 and not w2117;
w2119 <= a(23) and not w2113;
w2120 <= a(8) and w2119;
w2121 <= not w2118 and not w2120;
w2122 <= a(14) and a(17);
w2123 <= not w697 and not w2122;
w2124 <= w701 and w854;
w2125 <= a(6) and not w2124;
w2126 <= a(25) and w2125;
w2127 <= not w2123 and w2126;
w2128 <= a(25) and not w2127;
w2129 <= a(6) and w2128;
w2130 <= not w2124 and not w2127;
w2131 <= not w2123 and w2130;
w2132 <= not w2129 and not w2131;
w2133 <= not w2121 and not w2132;
w2134 <= not w2121 and not w2133;
w2135 <= not w2132 and not w2133;
w2136 <= not w2134 and not w2135;
w2137 <= a(27) and a(28);
w2138 <= w15 and w2137;
w2139 <= w58 and w1847;
w2140 <= a(28) and a(29);
w2141 <= w24 and w2140;
w2142 <= not w2139 and not w2141;
w2143 <= not w2138 and not w2142;
w2144 <= a(29) and not w2143;
w2145 <= a(2) and w2144;
w2146 <= a(3) and a(28);
w2147 <= a(4) and a(27);
w2148 <= not w2146 and not w2147;
w2149 <= not w2138 and not w2143;
w2150 <= not w2148 and w2149;
w2151 <= not w2145 and not w2150;
w2152 <= not w2136 and not w2151;
w2153 <= not w2136 and not w2152;
w2154 <= not w2151 and not w2152;
w2155 <= not w2153 and not w2154;
w2156 <= a(22) and a(31);
w2157 <= w156 and w2156;
w2158 <= a(10) and a(31);
w2159 <= w1005 and w2158;
w2160 <= w290 and w1380;
w2161 <= not w2159 and not w2160;
w2162 <= not w2157 and not w2161;
w2163 <= not w2157 and not w2162;
w2164 <= a(0) and a(31);
w2165 <= a(9) and a(22);
w2166 <= not w2164 and not w2165;
w2167 <= w2163 and not w2166;
w2168 <= a(21) and not w2162;
w2169 <= a(10) and w2168;
w2170 <= not w2167 and not w2169;
w2171 <= not w1972 and not w1981;
w2172 <= w554 and w955;
w2173 <= w624 and w1137;
w2174 <= w408 and w1296;
w2175 <= not w2173 and not w2174;
w2176 <= not w2172 and not w2175;
w2177 <= a(20) and not w2176;
w2178 <= a(11) and w2177;
w2179 <= not w2172 and not w2176;
w2180 <= a(12) and a(19);
w2181 <= a(13) and a(18);
w2182 <= not w2180 and not w2181;
w2183 <= w2179 and not w2182;
w2184 <= not w2178 and not w2183;
w2185 <= not w2171 and not w2184;
w2186 <= not w2171 and not w2185;
w2187 <= not w2184 and not w2185;
w2188 <= not w2186 and not w2187;
w2189 <= not w2170 and not w2188;
w2190 <= w2170 and not w2187;
w2191 <= not w2186 and w2190;
w2192 <= not w2189 and not w2191;
w2193 <= not w2155 and w2192;
w2194 <= w2155 and not w2192;
w2195 <= not w2193 and not w2194;
w2196 <= not w2106 and w2195;
w2197 <= w2106 and not w2195;
w2198 <= not w2196 and not w2197;
w2199 <= not w2105 and w2198;
w2200 <= w2105 and not w2198;
w2201 <= not w2199 and not w2200;
w2202 <= not w2084 and not w2087;
w2203 <= not w1998 and not w2012;
w2204 <= not w2021 and not w2024;
w2205 <= w2203 and w2204;
w2206 <= not w2203 and not w2204;
w2207 <= not w2205 and not w2206;
w2208 <= a(1) and a(30);
w2209 <= a(16) and w2208;
w2210 <= not a(16) and not w2208;
w2211 <= not w2209 and not w2210;
w2212 <= w1977 and w2211;
w2213 <= not w1977 and not w2211;
w2214 <= not w2212 and not w2213;
w2215 <= not w2055 and w2214;
w2216 <= w2055 and not w2214;
w2217 <= not w2215 and not w2216;
w2218 <= w2207 and w2217;
w2219 <= not w2207 and not w2217;
w2220 <= not w2218 and not w2219;
w2221 <= w2202 and not w2220;
w2222 <= not w2202 and w2220;
w2223 <= not w2221 and not w2222;
w2224 <= w2009 and w2042;
w2225 <= not w2009 and not w2042;
w2226 <= not w2224 and not w2225;
w2227 <= w2075 and not w2226;
w2228 <= not w2075 and w2226;
w2229 <= not w2227 and not w2228;
w2230 <= not w2061 and not w2078;
w2231 <= not w2229 and w2230;
w2232 <= w2229 and not w2230;
w2233 <= not w2231 and not w2232;
w2234 <= not w1987 and not w1991;
w2235 <= not w2233 and w2234;
w2236 <= w2233 and not w2234;
w2237 <= not w2235 and not w2236;
w2238 <= w2223 and w2237;
w2239 <= not w2223 and not w2237;
w2240 <= not w2238 and not w2239;
w2241 <= w2201 and w2240;
w2242 <= not w2201 and not w2240;
w2243 <= not w2241 and not w2242;
w2244 <= not w2104 and w2243;
w2245 <= w2104 and not w2243;
w2246 <= not w2244 and not w2245;
w2247 <= not w2097 and not w2100;
w2248 <= not w2096 and not w2247;
w2249 <= not w2246 and w2248;
w2250 <= w2246 and not w2248;
w2251 <= not w2249 and not w2250;
w2252 <= not w2245 and not w2248;
w2253 <= not w2244 and not w2252;
w2254 <= not w2199 and not w2241;
w2255 <= not w2222 and not w2238;
w2256 <= not w2232 and not w2236;
w2257 <= a(5) and a(27);
w2258 <= a(4) and a(28);
w2259 <= not w2257 and not w2258;
w2260 <= w32 and w2137;
w2261 <= a(23) and not w2260;
w2262 <= a(9) and w2261;
w2263 <= not w2259 and w2262;
w2264 <= not w2260 and not w2263;
w2265 <= not w2259 and w2264;
w2266 <= a(23) and not w2263;
w2267 <= a(9) and w2266;
w2268 <= not w2265 and not w2267;
w2269 <= a(25) and a(26);
w2270 <= w141 and w2269;
w2271 <= w118 and w2107;
w2272 <= w186 and w1710;
w2273 <= not w2271 and not w2272;
w2274 <= not w2270 and not w2273;
w2275 <= a(24) and not w2274;
w2276 <= a(8) and w2275;
w2277 <= not w2270 and not w2274;
w2278 <= a(6) and a(26);
w2279 <= a(7) and a(25);
w2280 <= not w2278 and not w2279;
w2281 <= w2277 and not w2280;
w2282 <= not w2276 and not w2281;
w2283 <= not w2268 and not w2282;
w2284 <= not w2268 and not w2283;
w2285 <= not w2282 and not w2283;
w2286 <= not w2284 and not w2285;
w2287 <= not w2212 and not w2215;
w2288 <= w2286 and w2287;
w2289 <= not w2286 and not w2287;
w2290 <= not w2288 and not w2289;
w2291 <= a(0) and a(32);
w2292 <= a(2) and a(30);
w2293 <= not w2291 and not w2292;
w2294 <= a(30) and a(32);
w2295 <= w2 and w2294;
w2296 <= not w2293 and not w2295;
w2297 <= w2209 and w2296;
w2298 <= not w2295 and not w2297;
w2299 <= not w2293 and w2298;
w2300 <= w2209 and not w2297;
w2301 <= not w2299 and not w2300;
w2302 <= w554 and w1296;
w2303 <= w624 and w1298;
w2304 <= w408 and w1300;
w2305 <= not w2303 and not w2304;
w2306 <= not w2302 and not w2305;
w2307 <= a(21) and not w2306;
w2308 <= a(11) and w2307;
w2309 <= not w2302 and not w2306;
w2310 <= a(12) and a(20);
w2311 <= a(13) and a(19);
w2312 <= not w2310 and not w2311;
w2313 <= w2309 and not w2312;
w2314 <= not w2308 and not w2313;
w2315 <= not w2301 and not w2314;
w2316 <= not w2301 and not w2315;
w2317 <= not w2314 and not w2315;
w2318 <= not w2316 and not w2317;
w2319 <= a(3) and a(29);
w2320 <= a(10) and a(22);
w2321 <= not w2319 and not w2320;
w2322 <= w2319 and w2320;
w2323 <= a(18) and not w2322;
w2324 <= a(14) and w2323;
w2325 <= not w2321 and w2324;
w2326 <= a(18) and not w2325;
w2327 <= a(14) and w2326;
w2328 <= not w2322 and not w2325;
w2329 <= not w2321 and w2328;
w2330 <= not w2327 and not w2329;
w2331 <= not w2318 and not w2330;
w2332 <= not w2318 and not w2331;
w2333 <= not w2330 and not w2331;
w2334 <= not w2332 and not w2333;
w2335 <= not w2290 and w2334;
w2336 <= w2290 and not w2334;
w2337 <= not w2335 and not w2336;
w2338 <= not w2256 and w2337;
w2339 <= w2256 and not w2337;
w2340 <= not w2338 and not w2339;
w2341 <= not w2255 and w2340;
w2342 <= w2255 and not w2340;
w2343 <= not w2341 and not w2342;
w2344 <= not w2206 and not w2218;
w2345 <= w2163 and w2179;
w2346 <= not w2163 and not w2179;
w2347 <= not w2345 and not w2346;
w2348 <= w2149 and not w2347;
w2349 <= not w2149 and w2347;
w2350 <= not w2348 and not w2349;
w2351 <= a(1) and a(31);
w2352 <= not w799 and not w2351;
w2353 <= w799 and w2351;
w2354 <= not w2352 and not w2353;
w2355 <= w2130 and not w2354;
w2356 <= not w2130 and w2354;
w2357 <= not w2355 and not w2356;
w2358 <= not w2114 and w2357;
w2359 <= w2114 and not w2357;
w2360 <= not w2358 and not w2359;
w2361 <= w2350 and w2360;
w2362 <= not w2350 and not w2360;
w2363 <= not w2361 and not w2362;
w2364 <= w2344 and not w2363;
w2365 <= not w2344 and w2363;
w2366 <= not w2364 and not w2365;
w2367 <= not w2185 and not w2189;
w2368 <= not w2225 and not w2228;
w2369 <= w2367 and w2368;
w2370 <= not w2367 and not w2368;
w2371 <= not w2369 and not w2370;
w2372 <= not w2133 and not w2152;
w2373 <= not w2371 and w2372;
w2374 <= w2371 and not w2372;
w2375 <= not w2373 and not w2374;
w2376 <= not w2193 and not w2196;
w2377 <= not w2375 and w2376;
w2378 <= w2375 and not w2376;
w2379 <= not w2377 and not w2378;
w2380 <= w2366 and w2379;
w2381 <= not w2366 and not w2379;
w2382 <= not w2380 and not w2381;
w2383 <= w2343 and w2382;
w2384 <= not w2343 and not w2382;
w2385 <= not w2383 and not w2384;
w2386 <= not w2254 and w2385;
w2387 <= w2254 and not w2385;
w2388 <= not w2386 and not w2387;
w2389 <= not w2253 and w2388;
w2390 <= w2253 and not w2388;
w2391 <= not w2389 and not w2390;
w2392 <= w2298 and w2309;
w2393 <= not w2298 and not w2309;
w2394 <= not w2392 and not w2393;
w2395 <= w2328 and not w2394;
w2396 <= not w2328 and w2394;
w2397 <= not w2395 and not w2396;
w2398 <= w2264 and w2277;
w2399 <= not w2264 and not w2277;
w2400 <= not w2398 and not w2399;
w2401 <= a(22) and a(33);
w2402 <= w255 and w2401;
w2403 <= w350 and w2156;
w2404 <= a(31) and a(33);
w2405 <= w2 and w2404;
w2406 <= not w2403 and not w2405;
w2407 <= not w2402 and not w2406;
w2408 <= a(31) and not w2407;
w2409 <= a(2) and w2408;
w2410 <= not w2402 and not w2407;
w2411 <= a(0) and a(33);
w2412 <= a(11) and a(22);
w2413 <= not w2411 and not w2412;
w2414 <= w2410 and not w2413;
w2415 <= not w2409 and not w2414;
w2416 <= w2400 and not w2415;
w2417 <= w2400 and not w2416;
w2418 <= not w2415 and not w2416;
w2419 <= not w2417 and not w2418;
w2420 <= not w2397 and w2419;
w2421 <= w2397 and not w2419;
w2422 <= not w2420 and not w2421;
w2423 <= a(29) and a(30);
w2424 <= w15 and w2423;
w2425 <= a(24) and a(30);
w2426 <= w285 and w2425;
w2427 <= not w2424 and not w2426;
w2428 <= a(4) and a(29);
w2429 <= a(9) and a(24);
w2430 <= w2428 and w2429;
w2431 <= not w2427 and not w2430;
w2432 <= not w2430 and not w2431;
w2433 <= not w2428 and not w2429;
w2434 <= w2432 and not w2433;
w2435 <= a(30) and not w2431;
w2436 <= a(3) and w2435;
w2437 <= not w2434 and not w2436;
w2438 <= a(5) and a(28);
w2439 <= a(25) and a(27);
w2440 <= w118 and w2439;
w2441 <= w138 and w2137;
w2442 <= a(8) and a(25);
w2443 <= w2438 and w2442;
w2444 <= not w2441 and not w2443;
w2445 <= not w2440 and not w2444;
w2446 <= w2438 and not w2445;
w2447 <= a(6) and a(27);
w2448 <= not w2442 and not w2447;
w2449 <= not w2440 and not w2445;
w2450 <= not w2448 and w2449;
w2451 <= not w2446 and not w2450;
w2452 <= not w2437 and not w2451;
w2453 <= not w2437 and not w2452;
w2454 <= not w2451 and not w2452;
w2455 <= not w2453 and not w2454;
w2456 <= a(15) and a(18);
w2457 <= not w854 and not w2456;
w2458 <= w697 and w858;
w2459 <= a(7) and not w2458;
w2460 <= a(26) and w2459;
w2461 <= not w2457 and w2460;
w2462 <= a(26) and not w2461;
w2463 <= a(7) and w2462;
w2464 <= not w2458 and not w2461;
w2465 <= not w2457 and w2464;
w2466 <= not w2463 and not w2465;
w2467 <= not w2455 and not w2466;
w2468 <= not w2455 and not w2467;
w2469 <= not w2466 and not w2467;
w2470 <= not w2468 and not w2469;
w2471 <= w2422 and w2470;
w2472 <= not w2422 and not w2470;
w2473 <= not w2471 and not w2472;
w2474 <= not w2346 and not w2349;
w2475 <= not w2315 and not w2331;
w2476 <= w2474 and w2475;
w2477 <= not w2474 and not w2475;
w2478 <= not w2476 and not w2477;
w2479 <= not w2283 and not w2289;
w2480 <= not w2478 and w2479;
w2481 <= w2478 and not w2479;
w2482 <= not w2480 and not w2481;
w2483 <= not w2336 and not w2338;
w2484 <= w2482 and not w2483;
w2485 <= not w2482 and w2483;
w2486 <= not w2484 and not w2485;
w2487 <= not w2473 and w2486;
w2488 <= w2473 and not w2486;
w2489 <= not w2487 and not w2488;
w2490 <= a(10) and a(23);
w2491 <= not w2353 and not w2490;
w2492 <= w2353 and w2490;
w2493 <= a(1) and a(32);
w2494 <= a(17) and not w2493;
w2495 <= not a(17) and w2493;
w2496 <= not w2494 and not w2495;
w2497 <= not w2492 and not w2496;
w2498 <= not w2491 and w2497;
w2499 <= not w2492 and not w2498;
w2500 <= not w2491 and w2499;
w2501 <= not w2496 and not w2498;
w2502 <= not w2500 and not w2501;
w2503 <= w551 and w1296;
w2504 <= w412 and w1298;
w2505 <= w554 and w1300;
w2506 <= not w2504 and not w2505;
w2507 <= not w2503 and not w2506;
w2508 <= a(21) and not w2507;
w2509 <= a(12) and w2508;
w2510 <= not w2503 and not w2507;
w2511 <= a(13) and a(20);
w2512 <= a(14) and a(19);
w2513 <= not w2511 and not w2512;
w2514 <= w2510 and not w2513;
w2515 <= not w2509 and not w2514;
w2516 <= not w2502 and not w2515;
w2517 <= not w2502 and not w2516;
w2518 <= not w2515 and not w2516;
w2519 <= not w2517 and not w2518;
w2520 <= not w2356 and not w2358;
w2521 <= w2519 and w2520;
w2522 <= not w2519 and not w2520;
w2523 <= not w2521 and not w2522;
w2524 <= not w2370 and not w2374;
w2525 <= not w2523 and w2524;
w2526 <= w2523 and not w2524;
w2527 <= not w2525 and not w2526;
w2528 <= not w2361 and not w2365;
w2529 <= not w2527 and w2528;
w2530 <= w2527 and not w2528;
w2531 <= not w2529 and not w2530;
w2532 <= not w2378 and not w2380;
w2533 <= w2531 and not w2532;
w2534 <= not w2531 and w2532;
w2535 <= not w2533 and not w2534;
w2536 <= w2489 and w2535;
w2537 <= not w2489 and not w2535;
w2538 <= not w2536 and not w2537;
w2539 <= not w2341 and not w2383;
w2540 <= not w2538 and w2539;
w2541 <= w2538 and not w2539;
w2542 <= not w2540 and not w2541;
w2543 <= not w2253 and not w2387;
w2544 <= not w2386 and not w2543;
w2545 <= not w2542 and w2544;
w2546 <= w2542 and not w2544;
w2547 <= not w2545 and not w2546;
w2548 <= not w2540 and not w2544;
w2549 <= not w2541 and not w2548;
w2550 <= not w2533 and not w2536;
w2551 <= w2499 and w2510;
w2552 <= not w2499 and not w2510;
w2553 <= not w2551 and not w2552;
w2554 <= a(11) and a(23);
w2555 <= a(12) and a(22);
w2556 <= not w2554 and not w2555;
w2557 <= w408 and w1725;
w2558 <= a(2) and not w2557;
w2559 <= a(32) and w2558;
w2560 <= not w2556 and w2559;
w2561 <= a(32) and not w2560;
w2562 <= a(2) and w2561;
w2563 <= not w2557 and not w2560;
w2564 <= not w2556 and w2563;
w2565 <= not w2562 and not w2564;
w2566 <= w2553 and not w2565;
w2567 <= w2553 and not w2566;
w2568 <= not w2565 and not w2566;
w2569 <= not w2567 and not w2568;
w2570 <= not w2516 and not w2522;
w2571 <= w2569 and w2570;
w2572 <= not w2569 and not w2570;
w2573 <= not w2571 and not w2572;
w2574 <= a(29) and w490;
w2575 <= a(24) and w2574;
w2576 <= w290 and w1710;
w2577 <= not w2575 and not w2576;
w2578 <= a(5) and a(29);
w2579 <= a(9) and a(25);
w2580 <= w2578 and w2579;
w2581 <= not w2577 and not w2580;
w2582 <= not w2580 and not w2581;
w2583 <= not w2578 and not w2579;
w2584 <= w2582 and not w2583;
w2585 <= a(24) and not w2581;
w2586 <= a(10) and w2585;
w2587 <= not w2584 and not w2586;
w2588 <= w701 and w1296;
w2589 <= w627 and w1298;
w2590 <= w551 and w1300;
w2591 <= not w2589 and not w2590;
w2592 <= not w2588 and not w2591;
w2593 <= a(21) and not w2592;
w2594 <= a(13) and w2593;
w2595 <= not w2588 and not w2592;
w2596 <= a(14) and a(20);
w2597 <= a(15) and a(19);
w2598 <= not w2596 and not w2597;
w2599 <= w2595 and not w2598;
w2600 <= not w2594 and not w2599;
w2601 <= not w2587 and not w2600;
w2602 <= not w2587 and not w2601;
w2603 <= not w2600 and not w2601;
w2604 <= not w2602 and not w2603;
w2605 <= w186 and w2033;
w2606 <= a(26) and a(28);
w2607 <= w118 and w2606;
w2608 <= w141 and w2137;
w2609 <= not w2607 and not w2608;
w2610 <= not w2605 and not w2609;
w2611 <= a(28) and not w2610;
w2612 <= a(6) and w2611;
w2613 <= not w2605 and not w2610;
w2614 <= a(7) and a(27);
w2615 <= a(8) and a(26);
w2616 <= not w2614 and not w2615;
w2617 <= w2613 and not w2616;
w2618 <= not w2612 and not w2617;
w2619 <= not w2604 and not w2618;
w2620 <= not w2604 and not w2619;
w2621 <= not w2618 and not w2619;
w2622 <= not w2620 and not w2621;
w2623 <= w2573 and not w2622;
w2624 <= not w2573 and w2622;
w2625 <= w2410 and w2432;
w2626 <= not w2410 and not w2432;
w2627 <= not w2625 and not w2626;
w2628 <= w2449 and not w2627;
w2629 <= not w2449 and w2627;
w2630 <= not w2628 and not w2629;
w2631 <= not w2452 and not w2467;
w2632 <= a(17) and w2493;
w2633 <= a(1) and a(33);
w2634 <= w856 and w2633;
w2635 <= not w856 and not w2633;
w2636 <= not w2634 and not w2635;
w2637 <= w2632 and w2636;
w2638 <= not w2632 and not w2636;
w2639 <= not w2637 and not w2638;
w2640 <= not w2464 and w2639;
w2641 <= w2464 and not w2639;
w2642 <= not w2640 and not w2641;
w2643 <= not w2631 and w2642;
w2644 <= w2631 and not w2642;
w2645 <= not w2643 and not w2644;
w2646 <= w2630 and w2645;
w2647 <= not w2630 and not w2645;
w2648 <= not w2646 and not w2647;
w2649 <= not w2624 and w2648;
w2650 <= not w2623 and w2649;
w2651 <= w2648 and not w2650;
w2652 <= not w2624 and not w2650;
w2653 <= not w2623 and w2652;
w2654 <= not w2651 and not w2653;
w2655 <= not w2526 and not w2530;
w2656 <= w2654 and w2655;
w2657 <= not w2654 and not w2655;
w2658 <= not w2656 and not w2657;
w2659 <= not w2484 and not w2487;
w2660 <= w2422 and not w2470;
w2661 <= not w2421 and not w2660;
w2662 <= not w2477 and not w2481;
w2663 <= w2661 and w2662;
w2664 <= not w2661 and not w2662;
w2665 <= not w2663 and not w2664;
w2666 <= not w2399 and not w2416;
w2667 <= not w2393 and not w2396;
w2668 <= a(31) and w8;
w2669 <= a(30) and w18;
w2670 <= not w2668 and not w2669;
w2671 <= a(30) and a(31);
w2672 <= w15 and w2671;
w2673 <= a(34) and not w2672;
w2674 <= not w2670 and w2673;
w2675 <= a(3) and a(31);
w2676 <= a(4) and a(30);
w2677 <= not w2675 and not w2676;
w2678 <= not w2672 and not w2677;
w2679 <= a(0) and a(34);
w2680 <= not w2678 and not w2679;
w2681 <= not w2674 and not w2680;
w2682 <= not w2667 and w2681;
w2683 <= w2667 and not w2681;
w2684 <= not w2682 and not w2683;
w2685 <= not w2666 and w2684;
w2686 <= w2666 and not w2684;
w2687 <= not w2685 and not w2686;
w2688 <= w2665 and w2687;
w2689 <= not w2665 and not w2687;
w2690 <= not w2688 and not w2689;
w2691 <= w2659 and not w2690;
w2692 <= not w2659 and w2690;
w2693 <= not w2691 and not w2692;
w2694 <= w2658 and w2693;
w2695 <= not w2658 and not w2693;
w2696 <= not w2694 and not w2695;
w2697 <= not w2550 and w2696;
w2698 <= w2550 and not w2696;
w2699 <= not w2697 and not w2698;
w2700 <= w2549 and not w2699;
w2701 <= not w2549 and not w2698;
w2702 <= not w2697 and w2701;
w2703 <= not w2700 and not w2702;
w2704 <= not w2697 and not w2701;
w2705 <= not w2692 and not w2694;
w2706 <= not w2650 and not w2657;
w2707 <= not w2626 and not w2629;
w2708 <= not w2637 and not w2640;
w2709 <= w2707 and w2708;
w2710 <= not w2707 and not w2708;
w2711 <= not w2709 and not w2710;
w2712 <= not w2552 and not w2566;
w2713 <= not w2711 and w2712;
w2714 <= w2711 and not w2712;
w2715 <= not w2713 and not w2714;
w2716 <= not w2643 and not w2646;
w2717 <= not w2715 and w2716;
w2718 <= w2715 and not w2716;
w2719 <= not w2717 and not w2718;
w2720 <= not w2572 and not w2623;
w2721 <= w2719 and not w2720;
w2722 <= not w2719 and w2720;
w2723 <= not w2721 and not w2722;
w2724 <= w2706 and not w2723;
w2725 <= not w2706 and w2723;
w2726 <= not w2724 and not w2725;
w2727 <= w118 and w1847;
w2728 <= a(27) and a(30);
w2729 <= w160 and w2728;
w2730 <= w138 and w2423;
w2731 <= not w2729 and not w2730;
w2732 <= not w2727 and not w2731;
w2733 <= not w2727 and not w2732;
w2734 <= a(6) and a(29);
w2735 <= not w2035 and not w2734;
w2736 <= w2733 and not w2735;
w2737 <= a(30) and not w2732;
w2738 <= a(5) and w2737;
w2739 <= not w2736 and not w2738;
w2740 <= a(16) and a(19);
w2741 <= not w858 and not w2740;
w2742 <= w858 and w2740;
w2743 <= a(7) and not w2742;
w2744 <= a(28) and w2743;
w2745 <= not w2741 and w2744;
w2746 <= a(28) and not w2745;
w2747 <= a(7) and w2746;
w2748 <= not w2742 and not w2745;
w2749 <= not w2741 and w2748;
w2750 <= not w2747 and not w2749;
w2751 <= not w2739 and not w2750;
w2752 <= not w2739 and not w2751;
w2753 <= not w2750 and not w2751;
w2754 <= not w2752 and not w2753;
w2755 <= a(9) and a(26);
w2756 <= a(10) and a(25);
w2757 <= not w2755 and not w2756;
w2758 <= w290 and w2269;
w2759 <= a(4) and not w2758;
w2760 <= a(31) and w2759;
w2761 <= not w2757 and w2760;
w2762 <= a(31) and not w2761;
w2763 <= a(4) and w2762;
w2764 <= not w2758 and not w2761;
w2765 <= not w2757 and w2764;
w2766 <= not w2763 and not w2765;
w2767 <= not w2754 and not w2766;
w2768 <= not w2754 and not w2767;
w2769 <= not w2766 and not w2767;
w2770 <= not w2768 and not w2769;
w2771 <= not w2682 and not w2685;
w2772 <= w2770 and w2771;
w2773 <= not w2770 and not w2771;
w2774 <= not w2772 and not w2773;
w2775 <= a(0) and a(35);
w2776 <= a(2) and a(33);
w2777 <= not w2775 and not w2776;
w2778 <= a(33) and a(35);
w2779 <= w2 and w2778;
w2780 <= not w2777 and not w2779;
w2781 <= w2634 and w2780;
w2782 <= not w2779 and not w2781;
w2783 <= not w2777 and w2782;
w2784 <= w2634 and not w2781;
w2785 <= not w2783 and not w2784;
w2786 <= a(3) and a(32);
w2787 <= a(11) and a(24);
w2788 <= a(12) and a(23);
w2789 <= not w2787 and not w2788;
w2790 <= w408 and w1472;
w2791 <= w2786 and not w2790;
w2792 <= not w2789 and w2791;
w2793 <= w2786 and not w2792;
w2794 <= not w2790 and not w2792;
w2795 <= not w2789 and w2794;
w2796 <= not w2793 and not w2795;
w2797 <= not w2785 and not w2796;
w2798 <= not w2785 and not w2797;
w2799 <= not w2796 and not w2797;
w2800 <= not w2798 and not w2799;
w2801 <= w701 and w1300;
w2802 <= w627 and w1499;
w2803 <= w551 and w1380;
w2804 <= not w2802 and not w2803;
w2805 <= not w2801 and not w2804;
w2806 <= a(22) and not w2805;
w2807 <= a(13) and w2806;
w2808 <= not w2801 and not w2805;
w2809 <= a(14) and a(21);
w2810 <= a(15) and a(20);
w2811 <= not w2809 and not w2810;
w2812 <= w2808 and not w2811;
w2813 <= not w2807 and not w2812;
w2814 <= not w2800 and not w2813;
w2815 <= not w2800 and not w2814;
w2816 <= not w2813 and not w2814;
w2817 <= not w2815 and not w2816;
w2818 <= w2774 and not w2817;
w2819 <= not w2774 and w2817;
w2820 <= not w2664 and not w2688;
w2821 <= w2563 and w2595;
w2822 <= not w2563 and not w2595;
w2823 <= not w2821 and not w2822;
w2824 <= not w2672 and not w2674;
w2825 <= not w2823 and w2824;
w2826 <= w2823 and not w2824;
w2827 <= not w2825 and not w2826;
w2828 <= not w2601 and not w2619;
w2829 <= a(34) and w781;
w2830 <= a(1) and a(34);
w2831 <= not a(18) and not w2830;
w2832 <= not w2829 and not w2831;
w2833 <= w2613 and not w2832;
w2834 <= not w2613 and w2832;
w2835 <= not w2833 and not w2834;
w2836 <= not w2582 and w2835;
w2837 <= w2582 and not w2835;
w2838 <= not w2836 and not w2837;
w2839 <= not w2828 and w2838;
w2840 <= w2828 and not w2838;
w2841 <= not w2839 and not w2840;
w2842 <= w2827 and w2841;
w2843 <= not w2827 and not w2841;
w2844 <= not w2842 and not w2843;
w2845 <= not w2820 and w2844;
w2846 <= w2820 and not w2844;
w2847 <= not w2845 and not w2846;
w2848 <= not w2819 and w2847;
w2849 <= not w2818 and w2848;
w2850 <= w2847 and not w2849;
w2851 <= not w2819 and not w2849;
w2852 <= not w2818 and w2851;
w2853 <= not w2850 and not w2852;
w2854 <= not w2726 and w2853;
w2855 <= w2726 and not w2853;
w2856 <= not w2854 and not w2855;
w2857 <= w2705 and not w2856;
w2858 <= not w2705 and w2856;
w2859 <= not w2857 and not w2858;
w2860 <= not w2704 and not w2859;
w2861 <= w2704 and w2859;
w2862 <= not w2860 and not w2861;
w2863 <= not w2725 and not w2855;
w2864 <= not w2845 and not w2849;
w2865 <= not w2822 and not w2826;
w2866 <= not w2834 and not w2836;
w2867 <= w2865 and w2866;
w2868 <= not w2865 and not w2866;
w2869 <= not w2867 and not w2868;
w2870 <= not w2797 and not w2814;
w2871 <= not w2869 and w2870;
w2872 <= w2869 and not w2870;
w2873 <= not w2871 and not w2872;
w2874 <= not w2839 and not w2842;
w2875 <= not w2873 and w2874;
w2876 <= w2873 and not w2874;
w2877 <= not w2875 and not w2876;
w2878 <= not w2773 and not w2818;
w2879 <= w2877 and not w2878;
w2880 <= not w2877 and w2878;
w2881 <= not w2879 and not w2880;
w2882 <= not w2864 and w2881;
w2883 <= w2864 and not w2881;
w2884 <= not w2882 and not w2883;
w2885 <= a(12) and a(24);
w2886 <= a(13) and a(23);
w2887 <= not w2885 and not w2886;
w2888 <= w554 and w1472;
w2889 <= a(2) and not w2888;
w2890 <= a(34) and w2889;
w2891 <= not w2887 and w2890;
w2892 <= not w2888 and not w2891;
w2893 <= not w2887 and w2892;
w2894 <= a(34) and not w2891;
w2895 <= a(2) and w2894;
w2896 <= not w2893 and not w2895;
w2897 <= a(9) and a(31);
w2898 <= w2257 and w2897;
w2899 <= w290 and w2033;
w2900 <= w2115 and w2158;
w2901 <= not w2899 and not w2900;
w2902 <= not w2898 and not w2901;
w2903 <= a(26) and not w2902;
w2904 <= a(10) and w2903;
w2905 <= not w2898 and not w2902;
w2906 <= a(5) and a(31);
w2907 <= a(9) and a(27);
w2908 <= not w2906 and not w2907;
w2909 <= w2905 and not w2908;
w2910 <= not w2904 and not w2909;
w2911 <= not w2896 and not w2910;
w2912 <= not w2896 and not w2911;
w2913 <= not w2910 and not w2911;
w2914 <= not w2912 and not w2913;
w2915 <= w186 and w2140;
w2916 <= a(28) and a(30);
w2917 <= w118 and w2916;
w2918 <= w141 and w2423;
w2919 <= not w2917 and not w2918;
w2920 <= not w2915 and not w2919;
w2921 <= a(30) and not w2920;
w2922 <= a(6) and w2921;
w2923 <= not w2915 and not w2920;
w2924 <= a(7) and a(29);
w2925 <= a(8) and a(28);
w2926 <= not w2924 and not w2925;
w2927 <= w2923 and not w2926;
w2928 <= not w2922 and not w2927;
w2929 <= not w2914 and not w2928;
w2930 <= not w2914 and not w2929;
w2931 <= not w2928 and not w2929;
w2932 <= not w2930 and not w2931;
w2933 <= not w2710 and not w2714;
w2934 <= a(0) and a(36);
w2935 <= w2829 and w2934;
w2936 <= w2829 and not w2935;
w2937 <= not w2829 and w2934;
w2938 <= not w2936 and not w2937;
w2939 <= a(1) and a(35);
w2940 <= a(17) and a(19);
w2941 <= w2939 and w2940;
w2942 <= w2939 and not w2941;
w2943 <= w2940 and not w2941;
w2944 <= not w2942 and not w2943;
w2945 <= not w2938 and not w2944;
w2946 <= not w2938 and not w2945;
w2947 <= not w2944 and not w2945;
w2948 <= not w2946 and not w2947;
w2949 <= a(32) and a(33);
w2950 <= w15 and w2949;
w2951 <= a(11) and a(25);
w2952 <= a(3) and a(33);
w2953 <= w2951 and w2952;
w2954 <= not w2950 and not w2953;
w2955 <= a(4) and a(32);
w2956 <= w2951 and w2955;
w2957 <= not w2954 and not w2956;
w2958 <= not w2956 and not w2957;
w2959 <= not w2951 and not w2955;
w2960 <= w2958 and not w2959;
w2961 <= w2952 and not w2957;
w2962 <= not w2960 and not w2961;
w2963 <= w697 and w1300;
w2964 <= w699 and w1499;
w2965 <= w701 and w1380;
w2966 <= not w2964 and not w2965;
w2967 <= not w2963 and not w2966;
w2968 <= a(22) and not w2967;
w2969 <= a(14) and w2968;
w2970 <= not w2963 and not w2967;
w2971 <= a(15) and a(21);
w2972 <= a(16) and a(20);
w2973 <= not w2971 and not w2972;
w2974 <= w2970 and not w2973;
w2975 <= not w2969 and not w2974;
w2976 <= not w2962 and not w2975;
w2977 <= not w2962 and not w2976;
w2978 <= not w2975 and not w2976;
w2979 <= not w2977 and not w2978;
w2980 <= not w2948 and w2979;
w2981 <= w2948 and not w2979;
w2982 <= not w2980 and not w2981;
w2983 <= not w2933 and not w2982;
w2984 <= not w2933 and not w2983;
w2985 <= not w2982 and not w2983;
w2986 <= not w2984 and not w2985;
w2987 <= not w2932 and not w2986;
w2988 <= not w2932 and not w2987;
w2989 <= not w2986 and not w2987;
w2990 <= not w2988 and not w2989;
w2991 <= not w2718 and not w2721;
w2992 <= w2733 and w2764;
w2993 <= not w2733 and not w2764;
w2994 <= not w2992 and not w2993;
w2995 <= w2748 and not w2994;
w2996 <= not w2748 and w2994;
w2997 <= not w2995 and not w2996;
w2998 <= w2794 and w2808;
w2999 <= not w2794 and not w2808;
w3000 <= not w2998 and not w2999;
w3001 <= w2782 and not w3000;
w3002 <= not w2782 and w3000;
w3003 <= not w3001 and not w3002;
w3004 <= not w2751 and not w2767;
w3005 <= not w3003 and w3004;
w3006 <= w3003 and not w3004;
w3007 <= not w3005 and not w3006;
w3008 <= w2997 and w3007;
w3009 <= not w2997 and not w3007;
w3010 <= not w3008 and not w3009;
w3011 <= not w2991 and w3010;
w3012 <= not w2991 and not w3011;
w3013 <= w3010 and not w3011;
w3014 <= not w3012 and not w3013;
w3015 <= not w2990 and not w3014;
w3016 <= w2990 and not w3013;
w3017 <= not w3012 and w3016;
w3018 <= not w3015 and not w3017;
w3019 <= w2884 and w3018;
w3020 <= not w2884 and not w3018;
w3021 <= not w3019 and not w3020;
w3022 <= w2863 and not w3021;
w3023 <= not w2863 and w3021;
w3024 <= not w3022 and not w3023;
w3025 <= not w2704 and not w2857;
w3026 <= not w2858 and not w3025;
w3027 <= not w3024 and w3026;
w3028 <= w3024 and not w3026;
w3029 <= not w3027 and not w3028;
w3030 <= not w2882 and not w3019;
w3031 <= not w2876 and not w2879;
w3032 <= not w2935 and not w2945;
w3033 <= w2905 and w3032;
w3034 <= not w2905 and not w3032;
w3035 <= not w3033 and not w3034;
w3036 <= w701 and w1725;
w3037 <= w627 and w1921;
w3038 <= w551 and w1472;
w3039 <= not w3037 and not w3038;
w3040 <= not w3036 and not w3039;
w3041 <= a(24) and not w3040;
w3042 <= a(13) and w3041;
w3043 <= a(14) and a(23);
w3044 <= a(15) and a(22);
w3045 <= not w3043 and not w3044;
w3046 <= not w3036 and not w3040;
w3047 <= not w3045 and w3046;
w3048 <= not w3042 and not w3047;
w3049 <= w3035 and not w3048;
w3050 <= w3035 and not w3049;
w3051 <= not w3048 and not w3049;
w3052 <= not w3050 and not w3051;
w3053 <= w2958 and w2970;
w3054 <= not w2958 and not w2970;
w3055 <= not w3053 and not w3054;
w3056 <= w2892 and not w3055;
w3057 <= not w2892 and w3055;
w3058 <= not w3056 and not w3057;
w3059 <= not w2948 and not w2979;
w3060 <= not w2976 and not w3059;
w3061 <= w3058 and not w3060;
w3062 <= not w3058 and w3060;
w3063 <= not w3061 and not w3062;
w3064 <= w3052 and w3063;
w3065 <= not w3052 and not w3063;
w3066 <= not w3064 and not w3065;
w3067 <= not w3031 and not w3066;
w3068 <= w3031 and w3066;
w3069 <= not w3067 and not w3068;
w3070 <= a(10) and a(32);
w3071 <= w2257 and w3070;
w3072 <= a(26) and a(32);
w3073 <= w308 and w3072;
w3074 <= w529 and w2033;
w3075 <= not w3073 and not w3074;
w3076 <= not w3071 and not w3075;
w3077 <= not w3071 and not w3076;
w3078 <= a(5) and a(32);
w3079 <= a(10) and a(27);
w3080 <= not w3078 and not w3079;
w3081 <= w3077 and not w3080;
w3082 <= a(26) and not w3076;
w3083 <= a(11) and w3082;
w3084 <= not w3081 and not w3083;
w3085 <= not w955 and not w1139;
w3086 <= w858 and w1296;
w3087 <= a(8) and not w3086;
w3088 <= a(29) and w3087;
w3089 <= not w3085 and w3088;
w3090 <= a(29) and not w3089;
w3091 <= a(8) and w3090;
w3092 <= not w3086 and not w3089;
w3093 <= not w3085 and w3092;
w3094 <= not w3091 and not w3093;
w3095 <= not w3084 and not w3094;
w3096 <= not w3084 and not w3095;
w3097 <= not w3094 and not w3095;
w3098 <= not w3096 and not w3097;
w3099 <= not w2999 and not w3002;
w3100 <= w3098 and w3099;
w3101 <= not w3098 and not w3099;
w3102 <= not w3100 and not w3101;
w3103 <= not w2868 and not w2872;
w3104 <= not w3102 and w3103;
w3105 <= w3102 and not w3103;
w3106 <= not w3104 and not w3105;
w3107 <= a(25) and a(33);
w3108 <= w550 and w3107;
w3109 <= a(25) and w288;
w3110 <= a(33) and w18;
w3111 <= not w3109 and not w3110;
w3112 <= a(37) and not w3108;
w3113 <= not w3111 and w3112;
w3114 <= not w3108 and not w3113;
w3115 <= a(4) and a(33);
w3116 <= a(12) and a(25);
w3117 <= not w3115 and not w3116;
w3118 <= w3114 and not w3117;
w3119 <= a(37) and not w3113;
w3120 <= a(0) and w3119;
w3121 <= not w3118 and not w3120;
w3122 <= a(2) and a(35);
w3123 <= a(3) and a(34);
w3124 <= not w3122 and not w3123;
w3125 <= a(34) and a(35);
w3126 <= w24 and w3125;
w3127 <= a(21) and not w3126;
w3128 <= a(16) and w3127;
w3129 <= not w3124 and w3128;
w3130 <= a(21) and not w3129;
w3131 <= a(16) and w3130;
w3132 <= not w3126 and not w3129;
w3133 <= not w3124 and w3132;
w3134 <= not w3131 and not w3133;
w3135 <= not w3121 and not w3134;
w3136 <= not w3121 and not w3135;
w3137 <= not w3134 and not w3135;
w3138 <= not w3136 and not w3137;
w3139 <= a(9) and a(28);
w3140 <= w141 and w2671;
w3141 <= w569 and w2916;
w3142 <= a(6) and a(31);
w3143 <= w3139 and w3142;
w3144 <= not w3141 and not w3143;
w3145 <= not w3140 and not w3144;
w3146 <= w3139 and not w3145;
w3147 <= not w3140 and not w3145;
w3148 <= a(7) and a(30);
w3149 <= not w3142 and not w3148;
w3150 <= w3147 and not w3149;
w3151 <= not w3146 and not w3150;
w3152 <= not w3138 and not w3151;
w3153 <= not w3138 and not w3152;
w3154 <= not w3151 and not w3152;
w3155 <= not w3153 and not w3154;
w3156 <= not w3106 and w3155;
w3157 <= w3106 and not w3155;
w3158 <= not w3156 and not w3157;
w3159 <= w3069 and w3158;
w3160 <= not w3069 and not w3158;
w3161 <= not w3159 and not w3160;
w3162 <= not w3011 and not w3015;
w3163 <= not w2983 and not w2987;
w3164 <= not w3006 and not w3008;
w3165 <= not w2911 and not w2929;
w3166 <= not w2993 and not w2996;
w3167 <= a(36) and w883;
w3168 <= a(1) and a(36);
w3169 <= not a(19) and not w3168;
w3170 <= not w3167 and not w3169;
w3171 <= w2941 and w3170;
w3172 <= w2941 and not w3171;
w3173 <= w3170 and not w3171;
w3174 <= not w3172 and not w3173;
w3175 <= not w2923 and not w3174;
w3176 <= w2923 and not w3173;
w3177 <= not w3172 and w3176;
w3178 <= not w3175 and not w3177;
w3179 <= not w3166 and w3178;
w3180 <= w3166 and not w3178;
w3181 <= not w3179 and not w3180;
w3182 <= not w3165 and w3181;
w3183 <= w3165 and not w3181;
w3184 <= not w3182 and not w3183;
w3185 <= not w3164 and w3184;
w3186 <= w3164 and not w3184;
w3187 <= not w3185 and not w3186;
w3188 <= not w3163 and w3187;
w3189 <= w3163 and not w3187;
w3190 <= not w3188 and not w3189;
w3191 <= not w3162 and w3190;
w3192 <= not w3162 and not w3191;
w3193 <= w3190 and not w3191;
w3194 <= not w3192 and not w3193;
w3195 <= w3161 and not w3194;
w3196 <= not w3161 and not w3193;
w3197 <= not w3192 and w3196;
w3198 <= not w3195 and not w3197;
w3199 <= not w3030 and w3198;
w3200 <= w3030 and not w3198;
w3201 <= not w3199 and not w3200;
w3202 <= not w3022 and not w3026;
w3203 <= not w3023 and not w3202;
w3204 <= not w3201 and w3203;
w3205 <= w3201 and not w3203;
w3206 <= not w3204 and not w3205;
w3207 <= not w3191 and not w3195;
w3208 <= not w3105 and not w3157;
w3209 <= not w3052 and w3063;
w3210 <= not w3061 and not w3209;
w3211 <= not w3208 and not w3210;
w3212 <= not w3208 and not w3211;
w3213 <= not w3210 and not w3211;
w3214 <= not w3212 and not w3213;
w3215 <= w3114 and w3132;
w3216 <= not w3114 and not w3132;
w3217 <= not w3215 and not w3216;
w3218 <= w3046 and not w3217;
w3219 <= not w3046 and w3217;
w3220 <= not w3218 and not w3219;
w3221 <= not w3095 and not w3101;
w3222 <= not w3220 and w3221;
w3223 <= w3220 and not w3221;
w3224 <= not w3222 and not w3223;
w3225 <= a(6) and a(32);
w3226 <= a(10) and a(28);
w3227 <= not w3225 and not w3226;
w3228 <= w138 and w2949;
w3229 <= a(5) and a(33);
w3230 <= w3226 and w3229;
w3231 <= not w3228 and not w3230;
w3232 <= w3225 and w3226;
w3233 <= not w3231 and not w3232;
w3234 <= not w3232 and not w3233;
w3235 <= not w3227 and w3234;
w3236 <= w3229 and not w3233;
w3237 <= not w3235 and not w3236;
w3238 <= w854 and w1380;
w3239 <= w697 and w1725;
w3240 <= a(17) and a(23);
w3241 <= w2971 and w3240;
w3242 <= not w3239 and not w3241;
w3243 <= not w3238 and not w3242;
w3244 <= a(23) and not w3243;
w3245 <= a(15) and w3244;
w3246 <= a(16) and a(22);
w3247 <= a(17) and a(21);
w3248 <= not w3246 and not w3247;
w3249 <= not w3238 and not w3243;
w3250 <= not w3248 and w3249;
w3251 <= not w3245 and not w3250;
w3252 <= not w3237 and not w3251;
w3253 <= not w3237 and not w3252;
w3254 <= not w3251 and not w3252;
w3255 <= not w3253 and not w3254;
w3256 <= a(9) and a(29);
w3257 <= w186 and w2671;
w3258 <= a(29) and a(31);
w3259 <= w569 and w3258;
w3260 <= w238 and w2423;
w3261 <= not w3259 and not w3260;
w3262 <= not w3257 and not w3261;
w3263 <= w3256 and not w3262;
w3264 <= not w3257 and not w3262;
w3265 <= a(7) and a(31);
w3266 <= a(8) and a(30);
w3267 <= not w3265 and not w3266;
w3268 <= w3264 and not w3267;
w3269 <= not w3263 and not w3268;
w3270 <= not w3255 and not w3269;
w3271 <= not w3255 and not w3270;
w3272 <= not w3269 and not w3270;
w3273 <= not w3271 and not w3272;
w3274 <= w3224 and not w3273;
w3275 <= not w3224 and w3273;
w3276 <= not w3214 and not w3275;
w3277 <= not w3274 and w3276;
w3278 <= not w3214 and not w3277;
w3279 <= not w3275 and not w3277;
w3280 <= not w3274 and w3279;
w3281 <= not w3278 and not w3280;
w3282 <= not w3067 and not w3159;
w3283 <= w3281 and w3282;
w3284 <= not w3281 and not w3282;
w3285 <= not w3283 and not w3284;
w3286 <= not w3185 and not w3188;
w3287 <= not w3034 and not w3049;
w3288 <= not w3135 and not w3152;
w3289 <= w3287 and w3288;
w3290 <= not w3287 and not w3288;
w3291 <= not w3289 and not w3290;
w3292 <= a(1) and a(37);
w3293 <= w1137 and w3292;
w3294 <= not w1137 and not w3292;
w3295 <= not w3293 and not w3294;
w3296 <= w3092 and not w3295;
w3297 <= not w3092 and w3295;
w3298 <= not w3296 and not w3297;
w3299 <= not w3147 and w3298;
w3300 <= w3147 and not w3298;
w3301 <= not w3299 and not w3300;
w3302 <= w3291 and w3301;
w3303 <= not w3291 and not w3301;
w3304 <= not w3302 and not w3303;
w3305 <= w3286 and not w3304;
w3306 <= not w3286 and w3304;
w3307 <= not w3305 and not w3306;
w3308 <= not w3171 and not w3175;
w3309 <= a(27) and a(34);
w3310 <= w455 and w3309;
w3311 <= w408 and w2033;
w3312 <= a(12) and a(34);
w3313 <= w2038 and w3312;
w3314 <= not w3311 and not w3313;
w3315 <= not w3310 and not w3314;
w3316 <= a(26) and not w3315;
w3317 <= a(12) and w3316;
w3318 <= not w3310 and not w3315;
w3319 <= a(4) and a(34);
w3320 <= a(11) and a(27);
w3321 <= not w3319 and not w3320;
w3322 <= w3318 and not w3321;
w3323 <= not w3317 and not w3322;
w3324 <= not w3308 and not w3323;
w3325 <= not w3308 and not w3324;
w3326 <= not w3323 and not w3324;
w3327 <= not w3325 and not w3326;
w3328 <= not w3054 and not w3057;
w3329 <= w3327 and w3328;
w3330 <= not w3327 and not w3328;
w3331 <= not w3329 and not w3330;
w3332 <= not w3179 and not w3182;
w3333 <= a(0) and a(38);
w3334 <= a(2) and a(36);
w3335 <= not w3333 and not w3334;
w3336 <= a(36) and a(38);
w3337 <= w2 and w3336;
w3338 <= not w3335 and not w3337;
w3339 <= w3167 and w3338;
w3340 <= not w3337 and not w3339;
w3341 <= not w3335 and w3340;
w3342 <= w3167 and not w3339;
w3343 <= not w3341 and not w3342;
w3344 <= w3077 and not w3343;
w3345 <= not w3077 and w3343;
w3346 <= not w3344 and not w3345;
w3347 <= a(13) and a(25);
w3348 <= a(14) and a(24);
w3349 <= not w3347 and not w3348;
w3350 <= w551 and w1710;
w3351 <= a(3) and not w3350;
w3352 <= a(35) and w3351;
w3353 <= not w3349 and w3352;
w3354 <= a(35) and not w3353;
w3355 <= a(3) and w3354;
w3356 <= not w3350 and not w3353;
w3357 <= not w3349 and w3356;
w3358 <= not w3355 and not w3357;
w3359 <= not w3346 and not w3358;
w3360 <= w3346 and w3358;
w3361 <= not w3359 and not w3360;
w3362 <= w3332 and not w3361;
w3363 <= not w3332 and w3361;
w3364 <= not w3362 and not w3363;
w3365 <= w3331 and w3364;
w3366 <= not w3331 and not w3364;
w3367 <= not w3365 and not w3366;
w3368 <= w3307 and w3367;
w3369 <= not w3307 and not w3367;
w3370 <= not w3368 and not w3369;
w3371 <= not w3285 and not w3370;
w3372 <= w3285 and w3370;
w3373 <= not w3371 and not w3372;
w3374 <= not w3207 and w3373;
w3375 <= w3207 and not w3373;
w3376 <= not w3374 and not w3375;
w3377 <= not w3200 and not w3203;
w3378 <= not w3199 and not w3377;
w3379 <= not w3376 and w3378;
w3380 <= w3376 and not w3378;
w3381 <= not w3379 and not w3380;
w3382 <= not w3284 and not w3372;
w3383 <= not w3306 and not w3368;
w3384 <= not w3363 and not w3365;
w3385 <= a(0) and a(39);
w3386 <= w3293 and w3385;
w3387 <= w3293 and not w3386;
w3388 <= not w3293 and w3385;
w3389 <= not w3387 and not w3388;
w3390 <= a(38) and w1009;
w3391 <= a(20) and not w3390;
w3392 <= a(1) and not w3390;
w3393 <= a(38) and w3392;
w3394 <= not w3391 and not w3393;
w3395 <= not w3389 and not w3394;
w3396 <= not w3389 and not w3395;
w3397 <= not w3394 and not w3395;
w3398 <= not w3396 and not w3397;
w3399 <= not w3297 and not w3299;
w3400 <= w3398 and w3399;
w3401 <= not w3398 and not w3399;
w3402 <= not w3400 and not w3401;
w3403 <= not w3216 and not w3219;
w3404 <= not w3402 and w3403;
w3405 <= w3402 and not w3403;
w3406 <= not w3404 and not w3405;
w3407 <= w3340 and w3356;
w3408 <= not w3340 and not w3356;
w3409 <= not w3407 and not w3408;
w3410 <= w3249 and not w3409;
w3411 <= not w3249 and w3409;
w3412 <= not w3410 and not w3411;
w3413 <= not w3252 and not w3270;
w3414 <= not w3077 and not w3343;
w3415 <= not w3359 and not w3414;
w3416 <= w3413 and w3415;
w3417 <= not w3413 and not w3415;
w3418 <= not w3416 and not w3417;
w3419 <= w3412 and w3418;
w3420 <= not w3412 and not w3418;
w3421 <= not w3419 and not w3420;
w3422 <= w3406 and w3421;
w3423 <= not w3406 and not w3421;
w3424 <= not w3422 and not w3423;
w3425 <= not w3384 and w3424;
w3426 <= w3384 and not w3424;
w3427 <= not w3425 and not w3426;
w3428 <= w3383 and not w3427;
w3429 <= not w3383 and w3427;
w3430 <= not w3428 and not w3429;
w3431 <= not w3211 and not w3277;
w3432 <= w3264 and w3318;
w3433 <= not w3264 and not w3318;
w3434 <= not w3432 and not w3433;
w3435 <= w3234 and not w3434;
w3436 <= not w3234 and w3434;
w3437 <= not w3435 and not w3436;
w3438 <= not w3324 and not w3330;
w3439 <= not w3437 and w3438;
w3440 <= w3437 and not w3438;
w3441 <= not w3439 and not w3440;
w3442 <= a(4) and a(35);
w3443 <= a(12) and a(27);
w3444 <= not w3442 and not w3443;
w3445 <= w3442 and w3443;
w3446 <= a(22) and not w3445;
w3447 <= a(17) and w3446;
w3448 <= not w3444 and w3447;
w3449 <= not w3445 and not w3448;
w3450 <= not w3444 and w3449;
w3451 <= a(22) and not w3448;
w3452 <= a(17) and w3451;
w3453 <= not w3450 and not w3452;
w3454 <= a(18) and a(21);
w3455 <= not w1296 and not w3454;
w3456 <= w955 and w1300;
w3457 <= a(8) and not w3456;
w3458 <= a(31) and w3457;
w3459 <= not w3455 and w3458;
w3460 <= a(31) and not w3459;
w3461 <= a(8) and w3460;
w3462 <= not w3456 and not w3459;
w3463 <= not w3455 and w3462;
w3464 <= not w3461 and not w3463;
w3465 <= not w3453 and not w3464;
w3466 <= not w3453 and not w3465;
w3467 <= not w3464 and not w3465;
w3468 <= not w3466 and not w3467;
w3469 <= a(34) and w2574;
w3470 <= a(5) and a(34);
w3471 <= w1782 and w3470;
w3472 <= w529 and w2140;
w3473 <= not w3471 and not w3472;
w3474 <= not w3469 and not w3473;
w3475 <= w1782 and not w3474;
w3476 <= not w3469 and not w3474;
w3477 <= a(10) and a(29);
w3478 <= not w3470 and not w3477;
w3479 <= w3476 and not w3478;
w3480 <= not w3475 and not w3479;
w3481 <= not w3468 and not w3480;
w3482 <= not w3468 and not w3481;
w3483 <= not w3480 and not w3481;
w3484 <= not w3482 and not w3483;
w3485 <= w3441 and not w3484;
w3486 <= not w3441 and w3484;
w3487 <= not w3431 and not w3486;
w3488 <= not w3485 and w3487;
w3489 <= not w3431 and not w3488;
w3490 <= not w3486 and not w3488;
w3491 <= not w3485 and w3490;
w3492 <= not w3489 and not w3491;
w3493 <= a(36) and a(37);
w3494 <= w24 and w3493;
w3495 <= a(13) and a(37);
w3496 <= w1796 and w3495;
w3497 <= not w3494 and not w3496;
w3498 <= a(3) and a(36);
w3499 <= a(13) and a(26);
w3500 <= w3498 and w3499;
w3501 <= not w3497 and not w3500;
w3502 <= not w3500 and not w3501;
w3503 <= not w3498 and not w3499;
w3504 <= w3502 and not w3503;
w3505 <= a(37) and not w3501;
w3506 <= a(2) and w3505;
w3507 <= not w3504 and not w3506;
w3508 <= w697 and w1472;
w3509 <= w699 and w1353;
w3510 <= w701 and w1710;
w3511 <= not w3509 and not w3510;
w3512 <= not w3508 and not w3511;
w3513 <= a(25) and not w3512;
w3514 <= a(14) and w3513;
w3515 <= not w3508 and not w3512;
w3516 <= a(15) and a(24);
w3517 <= a(16) and a(23);
w3518 <= not w3516 and not w3517;
w3519 <= w3515 and not w3518;
w3520 <= not w3514 and not w3519;
w3521 <= not w3507 and not w3520;
w3522 <= not w3507 and not w3521;
w3523 <= not w3520 and not w3521;
w3524 <= not w3522 and not w3523;
w3525 <= a(6) and a(33);
w3526 <= w569 and w2294;
w3527 <= w141 and w2949;
w3528 <= a(9) and a(30);
w3529 <= w3525 and w3528;
w3530 <= not w3527 and not w3529;
w3531 <= not w3526 and not w3530;
w3532 <= w3525 and not w3531;
w3533 <= not w3526 and not w3531;
w3534 <= a(7) and a(32);
w3535 <= not w3528 and not w3534;
w3536 <= w3533 and not w3535;
w3537 <= not w3532 and not w3536;
w3538 <= not w3524 and not w3537;
w3539 <= not w3524 and not w3538;
w3540 <= not w3537 and not w3538;
w3541 <= not w3539 and not w3540;
w3542 <= not w3290 and not w3302;
w3543 <= w3541 and w3542;
w3544 <= not w3541 and not w3542;
w3545 <= not w3543 and not w3544;
w3546 <= not w3223 and not w3274;
w3547 <= w3545 and not w3546;
w3548 <= not w3545 and w3546;
w3549 <= not w3547 and not w3548;
w3550 <= w3492 and w3549;
w3551 <= not w3492 and not w3549;
w3552 <= not w3550 and not w3551;
w3553 <= w3430 and not w3552;
w3554 <= not w3430 and w3552;
w3555 <= not w3553 and not w3554;
w3556 <= not w3382 and w3555;
w3557 <= w3382 and not w3555;
w3558 <= not w3556 and not w3557;
w3559 <= not w3375 and not w3378;
w3560 <= not w3374 and not w3559;
w3561 <= not w3558 and w3560;
w3562 <= w3558 and not w3560;
w3563 <= not w3561 and not w3562;
w3564 <= not w3557 and not w3560;
w3565 <= not w3556 and not w3564;
w3566 <= not w3429 and not w3553;
w3567 <= not w3492 and w3549;
w3568 <= not w3488 and not w3567;
w3569 <= not w3544 and not w3547;
w3570 <= not w3440 and not w3485;
w3571 <= w3476 and w3502;
w3572 <= not w3476 and not w3502;
w3573 <= not w3571 and not w3572;
w3574 <= w3449 and not w3573;
w3575 <= not w3449 and w3573;
w3576 <= not w3574 and not w3575;
w3577 <= not w3465 and not w3481;
w3578 <= not w3521 and not w3538;
w3579 <= w3577 and w3578;
w3580 <= not w3577 and not w3578;
w3581 <= not w3579 and not w3580;
w3582 <= w3576 and w3581;
w3583 <= not w3576 and not w3581;
w3584 <= not w3582 and not w3583;
w3585 <= not w3570 and w3584;
w3586 <= w3570 and not w3584;
w3587 <= not w3585 and not w3586;
w3588 <= not w3569 and w3587;
w3589 <= w3569 and not w3587;
w3590 <= not w3588 and not w3589;
w3591 <= not w3568 and w3590;
w3592 <= w3590 and not w3591;
w3593 <= not w3568 and not w3591;
w3594 <= not w3592 and not w3593;
w3595 <= w3515 and w3533;
w3596 <= not w3515 and not w3533;
w3597 <= not w3595 and not w3596;
w3598 <= not w3386 and not w3395;
w3599 <= not w3597 and w3598;
w3600 <= w3597 and not w3598;
w3601 <= not w3599 and not w3600;
w3602 <= not w3401 and not w3405;
w3603 <= not w3601 and w3602;
w3604 <= w3601 and not w3602;
w3605 <= not w3603 and not w3604;
w3606 <= a(0) and a(40);
w3607 <= a(2) and a(38);
w3608 <= not w3606 and not w3607;
w3609 <= a(38) and a(40);
w3610 <= w2 and w3609;
w3611 <= not w3608 and not w3610;
w3612 <= w1275 and w3611;
w3613 <= not w3610 and not w3612;
w3614 <= not w3608 and w3613;
w3615 <= w1275 and not w3612;
w3616 <= not w3614 and not w3615;
w3617 <= a(7) and a(33);
w3618 <= a(31) and a(32);
w3619 <= w238 and w3618;
w3620 <= w569 and w2404;
w3621 <= w186 and w2949;
w3622 <= not w3620 and not w3621;
w3623 <= not w3619 and not w3622;
w3624 <= w3617 and not w3623;
w3625 <= not w3619 and not w3623;
w3626 <= a(8) and a(32);
w3627 <= not w2897 and not w3626;
w3628 <= w3625 and not w3627;
w3629 <= not w3624 and not w3628;
w3630 <= not w3616 and not w3629;
w3631 <= not w3616 and not w3630;
w3632 <= not w3629 and not w3630;
w3633 <= not w3631 and not w3632;
w3634 <= a(35) and a(36);
w3635 <= w32 and w3634;
w3636 <= a(12) and a(36);
w3637 <= w2258 and w3636;
w3638 <= not w3635 and not w3637;
w3639 <= a(5) and a(35);
w3640 <= a(12) and a(28);
w3641 <= w3639 and w3640;
w3642 <= not w3638 and not w3641;
w3643 <= a(36) and not w3642;
w3644 <= a(4) and w3643;
w3645 <= not w3641 and not w3642;
w3646 <= not w3639 and not w3640;
w3647 <= w3645 and not w3646;
w3648 <= not w3644 and not w3647;
w3649 <= not w3633 and not w3648;
w3650 <= not w3633 and not w3649;
w3651 <= not w3648 and not w3649;
w3652 <= not w3650 and not w3651;
w3653 <= not w3605 and w3652;
w3654 <= w3605 and not w3652;
w3655 <= not w3653 and not w3654;
w3656 <= not w3422 and not w3425;
w3657 <= w3655 and not w3656;
w3658 <= not w3655 and w3656;
w3659 <= not w3657 and not w3658;
w3660 <= a(13) and a(27);
w3661 <= a(14) and a(26);
w3662 <= not w3660 and not w3661;
w3663 <= w551 and w2033;
w3664 <= a(3) and not w3663;
w3665 <= a(37) and w3664;
w3666 <= not w3662 and w3665;
w3667 <= not w3663 and not w3666;
w3668 <= not w3662 and w3667;
w3669 <= a(37) and not w3666;
w3670 <= a(3) and w3669;
w3671 <= not w3668 and not w3670;
w3672 <= w854 and w1472;
w3673 <= w799 and w1353;
w3674 <= w697 and w1710;
w3675 <= not w3673 and not w3674;
w3676 <= not w3672 and not w3675;
w3677 <= a(25) and not w3676;
w3678 <= a(15) and w3677;
w3679 <= not w3672 and not w3676;
w3680 <= a(16) and a(24);
w3681 <= not w3240 and not w3680;
w3682 <= w3679 and not w3681;
w3683 <= not w3678 and not w3682;
w3684 <= not w3671 and not w3683;
w3685 <= not w3671 and not w3684;
w3686 <= not w3683 and not w3684;
w3687 <= not w3685 and not w3686;
w3688 <= a(6) and a(34);
w3689 <= a(10) and a(30);
w3690 <= w3688 and w3689;
w3691 <= w529 and w2423;
w3692 <= a(11) and a(34);
w3693 <= w2734 and w3692;
w3694 <= not w3691 and not w3693;
w3695 <= not w3690 and not w3694;
w3696 <= a(29) and not w3695;
w3697 <= a(11) and w3696;
w3698 <= not w3690 and not w3695;
w3699 <= not w3688 and not w3689;
w3700 <= w3698 and not w3699;
w3701 <= not w3697 and not w3700;
w3702 <= not w3687 and not w3701;
w3703 <= not w3687 and not w3702;
w3704 <= not w3701 and not w3702;
w3705 <= not w3703 and not w3704;
w3706 <= not w3417 and not w3419;
w3707 <= not w3705 and not w3706;
w3708 <= w3705 and w3706;
w3709 <= not w3707 and not w3708;
w3710 <= not w3433 and not w3436;
w3711 <= not w3408 and not w3411;
w3712 <= w3710 and w3711;
w3713 <= not w3710 and not w3711;
w3714 <= not w3712 and not w3713;
w3715 <= a(1) and a(39);
w3716 <= w1298 and w3715;
w3717 <= not w1298 and not w3715;
w3718 <= not w3716 and not w3717;
w3719 <= w3390 and w3718;
w3720 <= not w3390 and not w3718;
w3721 <= not w3719 and not w3720;
w3722 <= not w3462 and w3721;
w3723 <= w3462 and not w3721;
w3724 <= not w3722 and not w3723;
w3725 <= w3714 and w3724;
w3726 <= not w3714 and not w3724;
w3727 <= not w3725 and not w3726;
w3728 <= w3709 and w3727;
w3729 <= not w3709 and not w3727;
w3730 <= not w3728 and not w3729;
w3731 <= w3659 and w3730;
w3732 <= not w3659 and not w3730;
w3733 <= not w3731 and not w3732;
w3734 <= not w3594 and w3733;
w3735 <= not w3593 and not w3733;
w3736 <= not w3592 and w3735;
w3737 <= not w3734 and not w3736;
w3738 <= not w3566 and w3737;
w3739 <= w3566 and not w3737;
w3740 <= not w3738 and not w3739;
w3741 <= w3565 and not w3740;
w3742 <= not w3565 and not w3739;
w3743 <= not w3738 and w3742;
w3744 <= not w3741 and not w3743;
w3745 <= not w3591 and not w3734;
w3746 <= not w3707 and not w3728;
w3747 <= not w3604 and not w3654;
w3748 <= w3613 and w3679;
w3749 <= not w3613 and not w3679;
w3750 <= not w3748 and not w3749;
w3751 <= w3667 and not w3750;
w3752 <= not w3667 and w3750;
w3753 <= not w3751 and not w3752;
w3754 <= not w3630 and not w3649;
w3755 <= not w3753 and w3754;
w3756 <= w3753 and not w3754;
w3757 <= not w3755 and not w3756;
w3758 <= a(40) and w1102;
w3759 <= a(1) and a(40);
w3760 <= not a(21) and not w3759;
w3761 <= not w3758 and not w3760;
w3762 <= w3625 and not w3761;
w3763 <= not w3625 and w3761;
w3764 <= not w3762 and not w3763;
w3765 <= not w3698 and w3764;
w3766 <= w3698 and not w3764;
w3767 <= not w3765 and not w3766;
w3768 <= w3757 and w3767;
w3769 <= not w3757 and not w3767;
w3770 <= not w3768 and not w3769;
w3771 <= not w3747 and w3770;
w3772 <= w3747 and not w3770;
w3773 <= not w3771 and not w3772;
w3774 <= w3746 and not w3773;
w3775 <= not w3746 and w3773;
w3776 <= not w3774 and not w3775;
w3777 <= not w3657 and not w3731;
w3778 <= not w3776 and w3777;
w3779 <= w3776 and not w3777;
w3780 <= not w3778 and not w3779;
w3781 <= not w3596 and not w3600;
w3782 <= not w3572 and not w3575;
w3783 <= w3781 and w3782;
w3784 <= not w3781 and not w3782;
w3785 <= not w3783 and not w3784;
w3786 <= not w3684 and not w3702;
w3787 <= not w3785 and w3786;
w3788 <= w3785 and not w3786;
w3789 <= not w3787 and not w3788;
w3790 <= a(39) and a(41);
w3791 <= w2 and w3790;
w3792 <= a(0) and a(41);
w3793 <= a(2) and a(39);
w3794 <= not w3792 and not w3793;
w3795 <= not w3791 and not w3794;
w3796 <= w3716 and w3795;
w3797 <= not w3716 and not w3795;
w3798 <= not w3796 and not w3797;
w3799 <= not w3645 and w3798;
w3800 <= w3645 and not w3798;
w3801 <= not w3799 and not w3800;
w3802 <= a(13) and a(28);
w3803 <= a(15) and a(26);
w3804 <= not w3802 and not w3803;
w3805 <= w627 and w2606;
w3806 <= a(3) and not w3805;
w3807 <= a(38) and w3806;
w3808 <= not w3804 and w3807;
w3809 <= a(38) and not w3808;
w3810 <= a(3) and w3809;
w3811 <= not w3805 and not w3808;
w3812 <= not w3804 and w3811;
w3813 <= not w3810 and not w3812;
w3814 <= w3801 and not w3813;
w3815 <= w3801 and not w3814;
w3816 <= not w3813 and not w3814;
w3817 <= not w3815 and not w3816;
w3818 <= not w3580 and not w3582;
w3819 <= not w3817 and not w3818;
w3820 <= not w3817 and not w3819;
w3821 <= not w3818 and not w3819;
w3822 <= not w3820 and not w3821;
w3823 <= not w3789 and w3822;
w3824 <= w3789 and not w3822;
w3825 <= not w3823 and not w3824;
w3826 <= not w3585 and not w3588;
w3827 <= a(6) and a(35);
w3828 <= a(11) and a(30);
w3829 <= not w3827 and not w3828;
w3830 <= a(30) and a(35);
w3831 <= w621 and w3830;
w3832 <= w138 and w3634;
w3833 <= a(30) and a(36);
w3834 <= w308 and w3833;
w3835 <= not w3832 and not w3834;
w3836 <= not w3831 and not w3835;
w3837 <= not w3831 and not w3836;
w3838 <= not w3829 and w3837;
w3839 <= a(36) and not w3836;
w3840 <= a(5) and w3839;
w3841 <= not w3838 and not w3840;
w3842 <= a(19) and a(22);
w3843 <= not w1300 and not w3842;
w3844 <= w1300 and w3842;
w3845 <= a(8) and not w3844;
w3846 <= a(33) and w3845;
w3847 <= not w3843 and w3846;
w3848 <= a(33) and not w3847;
w3849 <= a(8) and w3848;
w3850 <= not w3844 and not w3847;
w3851 <= not w3843 and w3850;
w3852 <= not w3849 and not w3851;
w3853 <= not w3841 and not w3852;
w3854 <= not w3841 and not w3853;
w3855 <= not w3852 and not w3853;
w3856 <= not w3854 and not w3855;
w3857 <= not w3719 and not w3722;
w3858 <= w3856 and w3857;
w3859 <= not w3856 and not w3857;
w3860 <= not w3858 and not w3859;
w3861 <= not w3713 and not w3725;
w3862 <= not w3860 and w3861;
w3863 <= w3860 and not w3861;
w3864 <= not w3862 and not w3863;
w3865 <= a(27) and a(37);
w3866 <= w696 and w3865;
w3867 <= w412 and w1847;
w3868 <= not w3866 and not w3867;
w3869 <= a(4) and a(37);
w3870 <= a(12) and a(29);
w3871 <= w3869 and w3870;
w3872 <= not w3868 and not w3871;
w3873 <= not w3871 and not w3872;
w3874 <= not w3869 and not w3870;
w3875 <= w3873 and not w3874;
w3876 <= a(27) and not w3872;
w3877 <= a(14) and w3876;
w3878 <= not w3875 and not w3877;
w3879 <= w858 and w1472;
w3880 <= w856 and w1353;
w3881 <= w854 and w1710;
w3882 <= not w3880 and not w3881;
w3883 <= not w3879 and not w3882;
w3884 <= a(25) and not w3883;
w3885 <= a(16) and w3884;
w3886 <= not w3879 and not w3883;
w3887 <= a(17) and a(24);
w3888 <= a(18) and a(23);
w3889 <= not w3887 and not w3888;
w3890 <= w3886 and not w3889;
w3891 <= not w3885 and not w3890;
w3892 <= not w3878 and not w3891;
w3893 <= not w3878 and not w3892;
w3894 <= not w3891 and not w3892;
w3895 <= not w3893 and not w3894;
w3896 <= a(32) and a(34);
w3897 <= w569 and w3896;
w3898 <= w290 and w3618;
w3899 <= a(7) and a(34);
w3900 <= w2158 and w3899;
w3901 <= not w3898 and not w3900;
w3902 <= not w3897 and not w3901;
w3903 <= w2158 and not w3902;
w3904 <= not w3897 and not w3902;
w3905 <= a(9) and a(32);
w3906 <= not w3899 and not w3905;
w3907 <= w3904 and not w3906;
w3908 <= not w3903 and not w3907;
w3909 <= not w3895 and not w3908;
w3910 <= not w3895 and not w3909;
w3911 <= not w3908 and not w3909;
w3912 <= not w3910 and not w3911;
w3913 <= not w3864 and w3912;
w3914 <= w3864 and not w3912;
w3915 <= not w3913 and not w3914;
w3916 <= not w3826 and w3915;
w3917 <= not w3826 and not w3916;
w3918 <= w3915 and not w3916;
w3919 <= not w3917 and not w3918;
w3920 <= w3825 and not w3919;
w3921 <= not w3825 and not w3918;
w3922 <= not w3917 and w3921;
w3923 <= not w3920 and not w3922;
w3924 <= w3780 and w3923;
w3925 <= not w3780 and not w3923;
w3926 <= not w3924 and not w3925;
w3927 <= w3745 and not w3926;
w3928 <= not w3745 and w3926;
w3929 <= not w3927 and not w3928;
w3930 <= not w3738 and not w3742;
w3931 <= not w3929 and w3930;
w3932 <= w3929 and not w3930;
w3933 <= not w3931 and not w3932;
w3934 <= not w3927 and not w3930;
w3935 <= not w3928 and not w3934;
w3936 <= not w3779 and not w3924;
w3937 <= not w3771 and not w3775;
w3938 <= not w3784 and not w3788;
w3939 <= a(7) and a(35);
w3940 <= a(11) and a(31);
w3941 <= w3939 and w3940;
w3942 <= a(31) and a(36);
w3943 <= w621 and w3942;
w3944 <= w141 and w3634;
w3945 <= not w3943 and not w3944;
w3946 <= not w3941 and not w3945;
w3947 <= a(6) and not w3946;
w3948 <= a(36) and w3947;
w3949 <= not w3941 and not w3946;
w3950 <= not w3939 and not w3940;
w3951 <= w3949 and not w3950;
w3952 <= not w3948 and not w3951;
w3953 <= w3904 and not w3952;
w3954 <= not w3904 and w3952;
w3955 <= not w3953 and not w3954;
w3956 <= a(33) and a(34);
w3957 <= w238 and w3956;
w3958 <= w184 and w3896;
w3959 <= w290 and w2949;
w3960 <= not w3958 and not w3959;
w3961 <= not w3957 and not w3960;
w3962 <= w3070 and not w3961;
w3963 <= not w3957 and not w3961;
w3964 <= a(8) and a(34);
w3965 <= a(9) and a(33);
w3966 <= not w3964 and not w3965;
w3967 <= w3963 and not w3966;
w3968 <= not w3962 and not w3967;
w3969 <= not w3955 and not w3968;
w3970 <= w3955 and w3968;
w3971 <= not w3969 and not w3970;
w3972 <= w3938 and not w3971;
w3973 <= not w3938 and w3971;
w3974 <= not w3972 and not w3973;
w3975 <= a(16) and a(40);
w3976 <= w1796 and w3975;
w3977 <= a(39) and a(40);
w3978 <= w24 and w3977;
w3979 <= not w3976 and not w3978;
w3980 <= a(3) and a(39);
w3981 <= a(16) and a(26);
w3982 <= w3980 and w3981;
w3983 <= not w3979 and not w3982;
w3984 <= not w3982 and not w3983;
w3985 <= not w3980 and not w3981;
w3986 <= w3984 and not w3985;
w3987 <= a(40) and not w3983;
w3988 <= a(2) and w3987;
w3989 <= not w3986 and not w3988;
w3990 <= w955 and w1472;
w3991 <= w1353 and w2940;
w3992 <= w858 and w1710;
w3993 <= not w3991 and not w3992;
w3994 <= not w3990 and not w3993;
w3995 <= a(25) and not w3994;
w3996 <= a(17) and w3995;
w3997 <= a(18) and a(24);
w3998 <= a(19) and a(23);
w3999 <= not w3997 and not w3998;
w4000 <= not w3990 and not w3994;
w4001 <= not w3999 and w4000;
w4002 <= not w3996 and not w4001;
w4003 <= not w3989 and not w4002;
w4004 <= not w3989 and not w4003;
w4005 <= not w4002 and not w4003;
w4006 <= not w4004 and not w4005;
w4007 <= a(14) and a(38);
w4008 <= w2258 and w4007;
w4009 <= w701 and w2137;
w4010 <= a(15) and a(38);
w4011 <= w2147 and w4010;
w4012 <= not w4009 and not w4011;
w4013 <= not w4008 and not w4012;
w4014 <= a(27) and not w4013;
w4015 <= a(15) and w4014;
w4016 <= not w4008 and not w4013;
w4017 <= a(4) and a(38);
w4018 <= a(14) and a(28);
w4019 <= not w4017 and not w4018;
w4020 <= w4016 and not w4019;
w4021 <= not w4015 and not w4020;
w4022 <= not w4006 and not w4021;
w4023 <= not w4006 and not w4022;
w4024 <= not w4021 and not w4022;
w4025 <= not w4023 and not w4024;
w4026 <= w3974 and not w4025;
w4027 <= not w3974 and w4025;
w4028 <= not w3937 and not w4027;
w4029 <= not w4026 and w4028;
w4030 <= not w3937 and not w4029;
w4031 <= not w4027 and not w4029;
w4032 <= not w4026 and w4031;
w4033 <= not w4030 and not w4032;
w4034 <= a(0) and a(42);
w4035 <= w3758 and w4034;
w4036 <= w3758 and not w4035;
w4037 <= not w3758 and w4034;
w4038 <= not w4036 and not w4037;
w4039 <= a(1) and a(41);
w4040 <= w1499 and w4039;
w4041 <= w4039 and not w4040;
w4042 <= w1499 and not w4040;
w4043 <= not w4041 and not w4042;
w4044 <= not w4038 and not w4043;
w4045 <= not w4038 and not w4044;
w4046 <= not w4043 and not w4044;
w4047 <= not w4045 and not w4046;
w4048 <= a(5) and a(37);
w4049 <= a(12) and a(30);
w4050 <= w4048 and w4049;
w4051 <= w554 and w2423;
w4052 <= w2578 and w3495;
w4053 <= not w4051 and not w4052;
w4054 <= not w4050 and not w4053;
w4055 <= a(29) and not w4054;
w4056 <= a(13) and w4055;
w4057 <= not w4050 and not w4054;
w4058 <= not w4048 and not w4049;
w4059 <= w4057 and not w4058;
w4060 <= not w4056 and not w4059;
w4061 <= not w4047 and not w4060;
w4062 <= not w4047 and not w4061;
w4063 <= not w4060 and not w4061;
w4064 <= not w4062 and not w4063;
w4065 <= not w3763 and not w3765;
w4066 <= w4064 and w4065;
w4067 <= not w4064 and not w4065;
w4068 <= not w4066 and not w4067;
w4069 <= not w3756 and not w3768;
w4070 <= not w4068 and w4069;
w4071 <= w4068 and not w4069;
w4072 <= not w4070 and not w4071;
w4073 <= w3850 and w3873;
w4074 <= not w3850 and not w3873;
w4075 <= not w4073 and not w4074;
w4076 <= w3837 and not w4075;
w4077 <= not w3837 and w4075;
w4078 <= not w4076 and not w4077;
w4079 <= not w3853 and not w3859;
w4080 <= not w4078 and w4079;
w4081 <= w4078 and not w4079;
w4082 <= not w4080 and not w4081;
w4083 <= w3811 and w3886;
w4084 <= not w3811 and not w3886;
w4085 <= not w4083 and not w4084;
w4086 <= not w3791 and not w3796;
w4087 <= not w4085 and w4086;
w4088 <= w4085 and not w4086;
w4089 <= not w4087 and not w4088;
w4090 <= w4082 and w4089;
w4091 <= not w4082 and not w4089;
w4092 <= not w4090 and not w4091;
w4093 <= w4072 and w4092;
w4094 <= not w4072 and not w4092;
w4095 <= not w4093 and not w4094;
w4096 <= w4033 and w4095;
w4097 <= not w4033 and not w4095;
w4098 <= not w4096 and not w4097;
w4099 <= not w3916 and not w3920;
w4100 <= not w3819 and not w3824;
w4101 <= not w3749 and not w3752;
w4102 <= not w3799 and not w3814;
w4103 <= w4101 and w4102;
w4104 <= not w4101 and not w4102;
w4105 <= not w4103 and not w4104;
w4106 <= not w3892 and not w3909;
w4107 <= not w4105 and w4106;
w4108 <= w4105 and not w4106;
w4109 <= not w4107 and not w4108;
w4110 <= not w3863 and not w3914;
w4111 <= w4109 and not w4110;
w4112 <= not w4109 and w4110;
w4113 <= not w4111 and not w4112;
w4114 <= not w4100 and w4113;
w4115 <= w4100 and not w4113;
w4116 <= not w4114 and not w4115;
w4117 <= not w4099 and w4116;
w4118 <= w4099 and not w4116;
w4119 <= not w4117 and not w4118;
w4120 <= not w4098 and w4119;
w4121 <= w4119 and not w4120;
w4122 <= not w4098 and not w4120;
w4123 <= not w4121 and not w4122;
w4124 <= not w3936 and not w4123;
w4125 <= w3936 and w4123;
w4126 <= not w4124 and not w4125;
w4127 <= not w3935 and w4126;
w4128 <= w3935 and not w4126;
w4129 <= not w4127 and not w4128;
w4130 <= not w4117 and not w4120;
w4131 <= not w4033 and w4095;
w4132 <= not w4029 and not w4131;
w4133 <= not w4071 and not w4093;
w4134 <= not w3973 and not w4026;
w4135 <= not w4003 and not w4022;
w4136 <= not w3904 and not w3952;
w4137 <= not w3969 and not w4136;
w4138 <= a(42) and w1211;
w4139 <= a(1) and a(42);
w4140 <= not a(22) and not w4139;
w4141 <= not w4138 and not w4140;
w4142 <= w4040 and w4141;
w4143 <= not w4040 and not w4141;
w4144 <= not w4142 and not w4143;
w4145 <= not w3963 and w4144;
w4146 <= w3963 and not w4144;
w4147 <= not w4145 and not w4146;
w4148 <= not w4137 and w4147;
w4149 <= not w4137 and not w4148;
w4150 <= w4147 and not w4148;
w4151 <= not w4149 and not w4150;
w4152 <= not w4135 and not w4151;
w4153 <= w4135 and not w4150;
w4154 <= not w4149 and w4153;
w4155 <= not w4152 and not w4154;
w4156 <= not w4134 and w4155;
w4157 <= w4134 and not w4155;
w4158 <= not w4156 and not w4157;
w4159 <= not w4133 and w4158;
w4160 <= w4133 and not w4158;
w4161 <= not w4159 and not w4160;
w4162 <= not w4132 and w4161;
w4163 <= not w4132 and not w4162;
w4164 <= w4161 and not w4162;
w4165 <= not w4163 and not w4164;
w4166 <= not w4111 and not w4114;
w4167 <= not w4104 and not w4108;
w4168 <= w15 and w3977;
w4169 <= a(4) and a(43);
w4170 <= w3385 and w4169;
w4171 <= not w4168 and not w4170;
w4172 <= a(0) and a(43);
w4173 <= a(3) and a(40);
w4174 <= w4172 and w4173;
w4175 <= not w4171 and not w4174;
w4176 <= not w4174 and not w4175;
w4177 <= not w4172 and not w4173;
w4178 <= w4176 and not w4177;
w4179 <= a(39) and not w4175;
w4180 <= a(4) and w4179;
w4181 <= not w4178 and not w4180;
w4182 <= w697 and w2137;
w4183 <= w699 and w1847;
w4184 <= w701 and w2140;
w4185 <= not w4183 and not w4184;
w4186 <= not w4182 and not w4185;
w4187 <= a(29) and not w4186;
w4188 <= a(14) and w4187;
w4189 <= not w4182 and not w4186;
w4190 <= a(15) and a(28);
w4191 <= a(16) and a(27);
w4192 <= not w4190 and not w4191;
w4193 <= w4189 and not w4192;
w4194 <= not w4188 and not w4193;
w4195 <= not w4181 and not w4194;
w4196 <= not w4181 and not w4195;
w4197 <= not w4194 and not w4195;
w4198 <= not w4196 and not w4197;
w4199 <= w955 and w1710;
w4200 <= w2107 and w2940;
w4201 <= w858 and w2269;
w4202 <= not w4200 and not w4201;
w4203 <= not w4199 and not w4202;
w4204 <= a(26) and not w4203;
w4205 <= a(17) and w4204;
w4206 <= a(18) and a(25);
w4207 <= not w1470 and not w4206;
w4208 <= not w4199 and not w4203;
w4209 <= not w4207 and w4208;
w4210 <= not w4205 and not w4209;
w4211 <= not w4198 and not w4210;
w4212 <= not w4198 and not w4211;
w4213 <= not w4210 and not w4211;
w4214 <= not w4212 and not w4213;
w4215 <= w184 and w2778;
w4216 <= w186 and w3634;
w4217 <= a(10) and a(36);
w4218 <= w3617 and w4217;
w4219 <= not w4216 and not w4218;
w4220 <= not w4215 and not w4219;
w4221 <= not w4215 and not w4220;
w4222 <= a(8) and a(35);
w4223 <= a(10) and a(33);
w4224 <= not w4222 and not w4223;
w4225 <= w4221 and not w4224;
w4226 <= a(36) and not w4220;
w4227 <= a(7) and w4226;
w4228 <= not w4225 and not w4227;
w4229 <= a(20) and a(23);
w4230 <= not w1380 and not w4229;
w4231 <= w1300 and w1725;
w4232 <= a(34) and not w4231;
w4233 <= a(9) and w4232;
w4234 <= not w4230 and w4233;
w4235 <= a(34) and not w4234;
w4236 <= a(9) and w4235;
w4237 <= not w4231 and not w4234;
w4238 <= not w4230 and w4237;
w4239 <= not w4236 and not w4238;
w4240 <= not w4228 and not w4239;
w4241 <= not w4228 and not w4240;
w4242 <= not w4239 and not w4240;
w4243 <= not w4241 and not w4242;
w4244 <= a(5) and a(38);
w4245 <= a(13) and a(30);
w4246 <= not w4244 and not w4245;
w4247 <= w4244 and w4245;
w4248 <= a(2) and not w4247;
w4249 <= a(41) and w4248;
w4250 <= not w4246 and w4249;
w4251 <= a(41) and not w4250;
w4252 <= a(2) and w4251;
w4253 <= not w4247 and not w4250;
w4254 <= not w4246 and w4253;
w4255 <= not w4252 and not w4254;
w4256 <= not w4243 and not w4255;
w4257 <= not w4243 and not w4256;
w4258 <= not w4255 and not w4256;
w4259 <= not w4257 and not w4258;
w4260 <= not w4214 and w4259;
w4261 <= w4214 and not w4259;
w4262 <= not w4260 and not w4261;
w4263 <= not w4167 and not w4262;
w4264 <= w4167 and w4262;
w4265 <= not w4263 and not w4264;
w4266 <= not w4166 and w4265;
w4267 <= w4166 and not w4265;
w4268 <= not w4266 and not w4267;
w4269 <= not w4061 and not w4067;
w4270 <= w3949 and w4016;
w4271 <= not w3949 and not w4016;
w4272 <= not w4270 and not w4271;
w4273 <= w4000 and not w4272;
w4274 <= not w4000 and w4272;
w4275 <= not w4273 and not w4274;
w4276 <= w3984 and w4057;
w4277 <= not w3984 and not w4057;
w4278 <= not w4276 and not w4277;
w4279 <= not w4035 and not w4044;
w4280 <= not w4278 and w4279;
w4281 <= w4278 and not w4279;
w4282 <= not w4280 and not w4281;
w4283 <= not w4275 and not w4282;
w4284 <= w4275 and w4282;
w4285 <= not w4283 and not w4284;
w4286 <= not w4269 and w4285;
w4287 <= w4269 and not w4285;
w4288 <= not w4286 and not w4287;
w4289 <= not w4074 and not w4077;
w4290 <= w408 and w3618;
w4291 <= a(12) and a(37);
w4292 <= w3142 and w4291;
w4293 <= not w4290 and not w4292;
w4294 <= a(6) and a(37);
w4295 <= a(11) and a(32);
w4296 <= w4294 and w4295;
w4297 <= not w4293 and not w4296;
w4298 <= a(31) and not w4297;
w4299 <= a(12) and w4298;
w4300 <= not w4296 and not w4297;
w4301 <= not w4294 and not w4295;
w4302 <= w4300 and not w4301;
w4303 <= not w4299 and not w4302;
w4304 <= not w4289 and not w4303;
w4305 <= not w4289 and not w4304;
w4306 <= not w4303 and not w4304;
w4307 <= not w4305 and not w4306;
w4308 <= not w4084 and not w4088;
w4309 <= w4307 and w4308;
w4310 <= not w4307 and not w4308;
w4311 <= not w4309 and not w4310;
w4312 <= not w4081 and not w4090;
w4313 <= w4311 and not w4312;
w4314 <= not w4311 and w4312;
w4315 <= not w4313 and not w4314;
w4316 <= w4288 and w4315;
w4317 <= not w4288 and not w4315;
w4318 <= not w4316 and not w4317;
w4319 <= w4268 and w4318;
w4320 <= not w4268 and not w4318;
w4321 <= not w4319 and not w4320;
w4322 <= not w4165 and w4321;
w4323 <= not w4164 and not w4321;
w4324 <= not w4163 and w4323;
w4325 <= not w4322 and not w4324;
w4326 <= not w4130 and w4325;
w4327 <= w4130 and not w4325;
w4328 <= not w4326 and not w4327;
w4329 <= not w3935 and not w4125;
w4330 <= not w4124 and not w4329;
w4331 <= not w4328 and w4330;
w4332 <= w4328 and not w4330;
w4333 <= not w4331 and not w4332;
w4334 <= not w4162 and not w4322;
w4335 <= not w4156 and not w4159;
w4336 <= not w4148 and not w4152;
w4337 <= a(15) and a(29);
w4338 <= a(17) and a(27);
w4339 <= not w4337 and not w4338;
w4340 <= w799 and w1847;
w4341 <= a(3) and not w4340;
w4342 <= a(41) and w4341;
w4343 <= not w4339 and w4342;
w4344 <= not w4340 and not w4343;
w4345 <= not w4339 and w4344;
w4346 <= a(41) and not w4343;
w4347 <= a(3) and w4346;
w4348 <= not w4345 and not w4347;
w4349 <= a(18) and a(26);
w4350 <= w1296 and w1710;
w4351 <= w1137 and w2107;
w4352 <= w955 and w2269;
w4353 <= not w4351 and not w4352;
w4354 <= not w4350 and not w4353;
w4355 <= w4349 and not w4354;
w4356 <= a(19) and a(25);
w4357 <= a(20) and a(24);
w4358 <= not w4356 and not w4357;
w4359 <= not w4350 and not w4354;
w4360 <= not w4358 and w4359;
w4361 <= not w4355 and not w4360;
w4362 <= not w4348 and not w4361;
w4363 <= not w4348 and not w4362;
w4364 <= not w4361 and not w4362;
w4365 <= not w4363 and not w4364;
w4366 <= a(6) and a(38);
w4367 <= a(11) and a(37);
w4368 <= w3617 and w4367;
w4369 <= a(33) and a(38);
w4370 <= w621 and w4369;
w4371 <= a(37) and a(38);
w4372 <= w141 and w4371;
w4373 <= not w4370 and not w4372;
w4374 <= not w4368 and not w4373;
w4375 <= w4366 and not w4374;
w4376 <= not w4368 and not w4374;
w4377 <= a(7) and a(37);
w4378 <= a(11) and a(33);
w4379 <= not w4377 and not w4378;
w4380 <= w4376 and not w4379;
w4381 <= not w4375 and not w4380;
w4382 <= not w4365 and not w4381;
w4383 <= not w4365 and not w4382;
w4384 <= not w4381 and not w4382;
w4385 <= not w4383 and not w4384;
w4386 <= w2258 and w3975;
w4387 <= w699 and w2916;
w4388 <= not w4386 and not w4387;
w4389 <= a(4) and a(40);
w4390 <= a(14) and a(30);
w4391 <= w4389 and w4390;
w4392 <= not w4388 and not w4391;
w4393 <= not w4391 and not w4392;
w4394 <= not w4389 and not w4390;
w4395 <= w4393 and not w4394;
w4396 <= a(28) and not w4392;
w4397 <= a(16) and w4396;
w4398 <= not w4395 and not w4397;
w4399 <= a(8) and a(36);
w4400 <= w290 and w3125;
w4401 <= a(34) and a(36);
w4402 <= w184 and w4401;
w4403 <= w238 and w3634;
w4404 <= not w4402 and not w4403;
w4405 <= not w4400 and not w4404;
w4406 <= w4399 and not w4405;
w4407 <= not w4400 and not w4405;
w4408 <= a(9) and a(35);
w4409 <= a(10) and a(34);
w4410 <= not w4408 and not w4409;
w4411 <= w4407 and not w4410;
w4412 <= not w4406 and not w4411;
w4413 <= not w4398 and not w4412;
w4414 <= not w4398 and not w4413;
w4415 <= not w4412 and not w4413;
w4416 <= not w4414 and not w4415;
w4417 <= a(12) and a(32);
w4418 <= a(13) and a(31);
w4419 <= not w4417 and not w4418;
w4420 <= w554 and w3618;
w4421 <= a(5) and not w4420;
w4422 <= a(39) and w4421;
w4423 <= not w4419 and w4422;
w4424 <= a(39) and not w4423;
w4425 <= a(5) and w4424;
w4426 <= not w4420 and not w4423;
w4427 <= not w4419 and w4426;
w4428 <= not w4425 and not w4427;
w4429 <= not w4416 and not w4428;
w4430 <= not w4416 and not w4429;
w4431 <= not w4428 and not w4429;
w4432 <= not w4430 and not w4431;
w4433 <= w4385 and w4432;
w4434 <= not w4385 and not w4432;
w4435 <= not w4433 and not w4434;
w4436 <= not w4336 and w4435;
w4437 <= w4336 and not w4435;
w4438 <= not w4436 and not w4437;
w4439 <= w4335 and not w4438;
w4440 <= not w4335 and w4438;
w4441 <= not w4439 and not w4440;
w4442 <= w4189 and w4300;
w4443 <= not w4189 and not w4300;
w4444 <= not w4442 and not w4443;
w4445 <= a(42) and a(44);
w4446 <= w2 and w4445;
w4447 <= a(0) and a(44);
w4448 <= a(2) and a(42);
w4449 <= not w4447 and not w4448;
w4450 <= not w4446 and not w4449;
w4451 <= w4138 and w4450;
w4452 <= w4138 and not w4451;
w4453 <= not w4446 and not w4451;
w4454 <= not w4449 and w4453;
w4455 <= not w4452 and not w4454;
w4456 <= w4444 and not w4455;
w4457 <= w4444 and not w4456;
w4458 <= not w4455 and not w4456;
w4459 <= not w4457 and not w4458;
w4460 <= a(1) and a(43);
w4461 <= not w1173 and not w4460;
w4462 <= w1173 and w4460;
w4463 <= not w4461 and not w4462;
w4464 <= w4237 and not w4463;
w4465 <= not w4237 and w4463;
w4466 <= not w4464 and not w4465;
w4467 <= not w4221 and w4466;
w4468 <= w4221 and not w4466;
w4469 <= not w4467 and not w4468;
w4470 <= not w4459 and w4469;
w4471 <= not w4459 and not w4470;
w4472 <= w4469 and not w4470;
w4473 <= not w4471 and not w4472;
w4474 <= not w4304 and not w4310;
w4475 <= w4473 and w4474;
w4476 <= not w4473 and not w4474;
w4477 <= not w4475 and not w4476;
w4478 <= not w4284 and not w4286;
w4479 <= not w4277 and not w4281;
w4480 <= not w4142 and not w4145;
w4481 <= w4479 and w4480;
w4482 <= not w4479 and not w4480;
w4483 <= not w4481 and not w4482;
w4484 <= not w4271 and not w4274;
w4485 <= not w4483 and w4484;
w4486 <= w4483 and not w4484;
w4487 <= not w4485 and not w4486;
w4488 <= not w4478 and w4487;
w4489 <= w4478 and not w4487;
w4490 <= not w4488 and not w4489;
w4491 <= not w4477 and not w4490;
w4492 <= w4477 and w4490;
w4493 <= w4441 and not w4492;
w4494 <= not w4491 and w4493;
w4495 <= w4441 and not w4494;
w4496 <= not w4492 and not w4494;
w4497 <= not w4491 and w4496;
w4498 <= not w4495 and not w4497;
w4499 <= not w4266 and not w4319;
w4500 <= not w4313 and not w4316;
w4501 <= not w4214 and not w4259;
w4502 <= not w4263 and not w4501;
w4503 <= w4176 and w4253;
w4504 <= not w4176 and not w4253;
w4505 <= not w4503 and not w4504;
w4506 <= w4208 and not w4505;
w4507 <= not w4208 and w4505;
w4508 <= not w4506 and not w4507;
w4509 <= not w4240 and not w4256;
w4510 <= not w4195 and not w4211;
w4511 <= w4509 and w4510;
w4512 <= not w4509 and not w4510;
w4513 <= not w4511 and not w4512;
w4514 <= w4508 and w4513;
w4515 <= not w4508 and not w4513;
w4516 <= not w4514 and not w4515;
w4517 <= not w4502 and w4516;
w4518 <= w4502 and not w4516;
w4519 <= not w4517 and not w4518;
w4520 <= not w4500 and w4519;
w4521 <= w4500 and not w4519;
w4522 <= not w4520 and not w4521;
w4523 <= not w4499 and w4522;
w4524 <= w4499 and not w4522;
w4525 <= not w4523 and not w4524;
w4526 <= not w4498 and not w4525;
w4527 <= w4498 and w4525;
w4528 <= not w4526 and not w4527;
w4529 <= not w4334 and not w4528;
w4530 <= w4334 and w4528;
w4531 <= not w4529 and not w4530;
w4532 <= not w4327 and not w4330;
w4533 <= not w4326 and not w4532;
w4534 <= not w4531 and w4533;
w4535 <= w4531 and not w4533;
w4536 <= not w4534 and not w4535;
w4537 <= not w4434 and not w4436;
w4538 <= not w4488 and not w4492;
w4539 <= not w4537 and w4538;
w4540 <= w4537 and not w4538;
w4541 <= not w4539 and not w4540;
w4542 <= w4344 and w4453;
w4543 <= not w4344 and not w4453;
w4544 <= not w4542 and not w4543;
w4545 <= w4359 and not w4544;
w4546 <= not w4359 and w4544;
w4547 <= not w4545 and not w4546;
w4548 <= not w4482 and not w4486;
w4549 <= not w4547 and w4548;
w4550 <= w4547 and not w4548;
w4551 <= not w4549 and not w4550;
w4552 <= a(6) and a(39);
w4553 <= not w3692 and not w4552;
w4554 <= a(34) and a(39);
w4555 <= w621 and w4554;
w4556 <= a(12) and a(39);
w4557 <= w3525 and w4556;
w4558 <= w408 and w3956;
w4559 <= not w4557 and not w4558;
w4560 <= not w4555 and not w4559;
w4561 <= not w4555 and not w4560;
w4562 <= not w4553 and w4561;
w4563 <= a(33) and not w4560;
w4564 <= a(12) and w4563;
w4565 <= not w4562 and not w4564;
w4566 <= w854 and w2140;
w4567 <= w799 and w2916;
w4568 <= w697 and w2423;
w4569 <= not w4567 and not w4568;
w4570 <= not w4566 and not w4569;
w4571 <= a(30) and not w4570;
w4572 <= a(15) and w4571;
w4573 <= not w4566 and not w4570;
w4574 <= a(16) and a(29);
w4575 <= a(17) and a(28);
w4576 <= not w4574 and not w4575;
w4577 <= w4573 and not w4576;
w4578 <= not w4572 and not w4577;
w4579 <= not w4565 and not w4578;
w4580 <= not w4565 and not w4579;
w4581 <= not w4578 and not w4579;
w4582 <= not w4580 and not w4581;
w4583 <= a(44) and w1265;
w4584 <= a(1) and not w4583;
w4585 <= a(44) and w4584;
w4586 <= a(23) and not w4583;
w4587 <= not w4585 and not w4586;
w4588 <= a(3) and a(42);
w4589 <= not w4462 and not w4588;
w4590 <= w4462 and w4588;
w4591 <= not w4587 and not w4590;
w4592 <= not w4589 and w4591;
w4593 <= not w4587 and not w4592;
w4594 <= not w4590 and not w4592;
w4595 <= not w4589 and w4594;
w4596 <= not w4593 and not w4595;
w4597 <= not w4582 and not w4596;
w4598 <= not w4582 and not w4597;
w4599 <= not w4596 and not w4597;
w4600 <= not w4598 and not w4599;
w4601 <= w4551 and not w4600;
w4602 <= not w4551 and w4600;
w4603 <= not w4541 and not w4602;
w4604 <= not w4601 and w4603;
w4605 <= not w4541 and not w4604;
w4606 <= not w4602 and not w4604;
w4607 <= not w4601 and w4606;
w4608 <= not w4605 and not w4607;
w4609 <= not w4440 and not w4494;
w4610 <= w4608 and w4609;
w4611 <= not w4608 and not w4609;
w4612 <= not w4610 and not w4611;
w4613 <= a(41) and a(43);
w4614 <= w58 and w4613;
w4615 <= a(41) and a(45);
w4616 <= w18 and w4615;
w4617 <= a(43) and a(45);
w4618 <= w2 and w4617;
w4619 <= not w4616 and not w4618;
w4620 <= not w4614 and not w4619;
w4621 <= not w4614 and not w4620;
w4622 <= a(2) and a(43);
w4623 <= a(4) and a(41);
w4624 <= not w4622 and not w4623;
w4625 <= w4621 and not w4624;
w4626 <= a(45) and not w4620;
w4627 <= a(0) and w4626;
w4628 <= not w4625 and not w4627;
w4629 <= a(7) and a(38);
w4630 <= w238 and w3493;
w4631 <= w569 and w3336;
w4632 <= w186 and w4371;
w4633 <= not w4631 and not w4632;
w4634 <= not w4630 and not w4633;
w4635 <= w4629 and not w4634;
w4636 <= a(8) and a(37);
w4637 <= a(9) and a(36);
w4638 <= not w4636 and not w4637;
w4639 <= not w4630 and not w4634;
w4640 <= not w4638 and w4639;
w4641 <= not w4635 and not w4640;
w4642 <= not w4628 and not w4641;
w4643 <= not w4628 and not w4642;
w4644 <= not w4641 and not w4642;
w4645 <= not w4643 and not w4644;
w4646 <= not w1589 and not w1725;
w4647 <= w1380 and w1472;
w4648 <= a(35) and not w4647;
w4649 <= a(10) and w4648;
w4650 <= not w4646 and w4649;
w4651 <= a(35) and not w4650;
w4652 <= a(10) and w4651;
w4653 <= not w4647 and not w4650;
w4654 <= not w4646 and w4653;
w4655 <= not w4652 and not w4654;
w4656 <= not w4645 and not w4655;
w4657 <= not w4645 and not w4656;
w4658 <= not w4655 and not w4656;
w4659 <= not w4657 and not w4658;
w4660 <= w551 and w3618;
w4661 <= a(14) and a(40);
w4662 <= w2906 and w4661;
w4663 <= not w4660 and not w4662;
w4664 <= a(5) and a(40);
w4665 <= a(13) and a(32);
w4666 <= w4664 and w4665;
w4667 <= not w4663 and not w4666;
w4668 <= not w4666 and not w4667;
w4669 <= not w4664 and not w4665;
w4670 <= w4668 and not w4669;
w4671 <= a(31) and not w4667;
w4672 <= a(14) and w4671;
w4673 <= not w4670 and not w4672;
w4674 <= w1296 and w2269;
w4675 <= w1137 and w2439;
w4676 <= w955 and w2033;
w4677 <= not w4675 and not w4676;
w4678 <= not w4674 and not w4677;
w4679 <= a(27) and not w4678;
w4680 <= a(18) and w4679;
w4681 <= not w4674 and not w4678;
w4682 <= a(19) and a(26);
w4683 <= not w1650 and not w4682;
w4684 <= w4681 and not w4683;
w4685 <= not w4680 and not w4684;
w4686 <= not w4407 and not w4685;
w4687 <= not w4407 and not w4686;
w4688 <= not w4685 and not w4686;
w4689 <= not w4687 and not w4688;
w4690 <= not w4673 and not w4689;
w4691 <= not w4673 and not w4690;
w4692 <= not w4689 and not w4690;
w4693 <= not w4691 and not w4692;
w4694 <= not w4659 and not w4693;
w4695 <= not w4659 and not w4694;
w4696 <= not w4693 and not w4694;
w4697 <= not w4695 and not w4696;
w4698 <= not w4512 and not w4514;
w4699 <= not w4697 and not w4698;
w4700 <= not w4697 and not w4699;
w4701 <= not w4698 and not w4699;
w4702 <= not w4700 and not w4701;
w4703 <= not w4517 and not w4520;
w4704 <= w4702 and w4703;
w4705 <= not w4702 and not w4703;
w4706 <= not w4704 and not w4705;
w4707 <= not w4443 and not w4456;
w4708 <= not w4504 and not w4507;
w4709 <= w4707 and w4708;
w4710 <= not w4707 and not w4708;
w4711 <= not w4709 and not w4710;
w4712 <= not w4465 and not w4467;
w4713 <= not w4711 and w4712;
w4714 <= w4711 and not w4712;
w4715 <= not w4713 and not w4714;
w4716 <= not w4470 and not w4476;
w4717 <= not w4715 and w4716;
w4718 <= w4715 and not w4716;
w4719 <= not w4717 and not w4718;
w4720 <= w4376 and w4393;
w4721 <= not w4376 and not w4393;
w4722 <= not w4720 and not w4721;
w4723 <= w4426 and not w4722;
w4724 <= not w4426 and w4722;
w4725 <= not w4723 and not w4724;
w4726 <= not w4413 and not w4429;
w4727 <= not w4362 and not w4382;
w4728 <= w4726 and w4727;
w4729 <= not w4726 and not w4727;
w4730 <= not w4728 and not w4729;
w4731 <= w4725 and w4730;
w4732 <= not w4725 and not w4730;
w4733 <= not w4731 and not w4732;
w4734 <= w4719 and w4733;
w4735 <= not w4719 and not w4733;
w4736 <= not w4734 and not w4735;
w4737 <= w4706 and w4736;
w4738 <= not w4706 and not w4736;
w4739 <= w4612 and not w4738;
w4740 <= not w4737 and w4739;
w4741 <= w4612 and not w4740;
w4742 <= not w4738 and not w4740;
w4743 <= not w4737 and w4742;
w4744 <= not w4741 and not w4743;
w4745 <= not w4498 and w4525;
w4746 <= not w4523 and not w4745;
w4747 <= not w4744 and not w4746;
w4748 <= w4744 and w4746;
w4749 <= not w4747 and not w4748;
w4750 <= not w4530 and not w4533;
w4751 <= not w4529 and not w4750;
w4752 <= not w4749 and w4751;
w4753 <= w4749 and not w4751;
w4754 <= not w4752 and not w4753;
w4755 <= not w4611 and not w4740;
w4756 <= not w4705 and not w4737;
w4757 <= not w4718 and not w4734;
w4758 <= not w4694 and not w4699;
w4759 <= w4757 and w4758;
w4760 <= not w4757 and not w4758;
w4761 <= not w4759 and not w4760;
w4762 <= a(5) and a(41);
w4763 <= a(15) and a(31);
w4764 <= not w4762 and not w4763;
w4765 <= a(31) and a(41);
w4766 <= w920 and w4765;
w4767 <= a(2) and not w4766;
w4768 <= a(44) and w4767;
w4769 <= not w4764 and w4768;
w4770 <= not w4766 and not w4769;
w4771 <= not w4764 and w4770;
w4772 <= a(44) and not w4769;
w4773 <= a(2) and w4772;
w4774 <= not w4771 and not w4773;
w4775 <= w551 and w2949;
w4776 <= w3225 and w4661;
w4777 <= not w4775 and not w4776;
w4778 <= a(6) and a(40);
w4779 <= a(13) and a(33);
w4780 <= w4778 and w4779;
w4781 <= not w4777 and not w4780;
w4782 <= a(32) and not w4781;
w4783 <= a(14) and w4782;
w4784 <= not w4780 and not w4781;
w4785 <= not w4778 and not w4779;
w4786 <= w4784 and not w4785;
w4787 <= not w4783 and not w4786;
w4788 <= not w4774 and not w4787;
w4789 <= not w4774 and not w4788;
w4790 <= not w4787 and not w4788;
w4791 <= not w4789 and not w4790;
w4792 <= not w4721 and not w4724;
w4793 <= w4791 and w4792;
w4794 <= not w4791 and not w4792;
w4795 <= not w4793 and not w4794;
w4796 <= w4573 and w4681;
w4797 <= not w4573 and not w4681;
w4798 <= not w4796 and not w4797;
w4799 <= w4561 and not w4798;
w4800 <= not w4561 and w4798;
w4801 <= not w4799 and not w4800;
w4802 <= not w4710 and not w4714;
w4803 <= not w4801 and w4802;
w4804 <= w4801 and not w4802;
w4805 <= not w4803 and not w4804;
w4806 <= w4795 and w4805;
w4807 <= not w4795 and not w4805;
w4808 <= not w4806 and not w4807;
w4809 <= w4761 and w4808;
w4810 <= not w4761 and not w4808;
w4811 <= not w4809 and not w4810;
w4812 <= not w4756 and w4811;
w4813 <= w4756 and not w4811;
w4814 <= not w4812 and not w4813;
w4815 <= w4755 and not w4814;
w4816 <= not w4755 and w4814;
w4817 <= not w4815 and not w4816;
w4818 <= not w4537 and not w4538;
w4819 <= not w4604 and not w4818;
w4820 <= not w4729 and not w4731;
w4821 <= a(0) and a(46);
w4822 <= a(4) and a(42);
w4823 <= not w4821 and not w4822;
w4824 <= a(42) and a(43);
w4825 <= w15 and w4824;
w4826 <= a(3) and a(46);
w4827 <= w4172 and w4826;
w4828 <= not w4825 and not w4827;
w4829 <= w4821 and w4822;
w4830 <= not w4828 and not w4829;
w4831 <= not w4829 and not w4830;
w4832 <= not w4823 and w4831;
w4833 <= a(43) and not w4830;
w4834 <= a(3) and w4833;
w4835 <= not w4832 and not w4834;
w4836 <= w529 and w3634;
w4837 <= a(35) and a(37);
w4838 <= w882 and w4837;
w4839 <= w290 and w3493;
w4840 <= not w4838 and not w4839;
w4841 <= not w4836 and not w4840;
w4842 <= a(37) and not w4841;
w4843 <= a(9) and w4842;
w4844 <= not w4836 and not w4841;
w4845 <= a(11) and a(35);
w4846 <= not w4217 and not w4845;
w4847 <= w4844 and not w4846;
w4848 <= not w4843 and not w4847;
w4849 <= not w4835 and not w4848;
w4850 <= not w4835 and not w4849;
w4851 <= not w4848 and not w4849;
w4852 <= not w4850 and not w4851;
w4853 <= w1300 and w2269;
w4854 <= w1298 and w2439;
w4855 <= w1296 and w2033;
w4856 <= not w4854 and not w4855;
w4857 <= not w4853 and not w4856;
w4858 <= a(27) and not w4857;
w4859 <= a(19) and w4858;
w4860 <= not w4853 and not w4857;
w4861 <= a(20) and a(26);
w4862 <= a(21) and a(25);
w4863 <= not w4861 and not w4862;
w4864 <= w4860 and not w4863;
w4865 <= not w4859 and not w4864;
w4866 <= not w4852 and not w4865;
w4867 <= not w4852 and not w4866;
w4868 <= not w4865 and not w4866;
w4869 <= not w4867 and not w4868;
w4870 <= w858 and w2140;
w4871 <= w856 and w2916;
w4872 <= w854 and w2423;
w4873 <= not w4871 and not w4872;
w4874 <= not w4870 and not w4873;
w4875 <= a(30) and not w4874;
w4876 <= a(16) and w4875;
w4877 <= not w4870 and not w4874;
w4878 <= a(17) and a(29);
w4879 <= a(18) and a(28);
w4880 <= not w4878 and not w4879;
w4881 <= w4877 and not w4880;
w4882 <= not w4876 and not w4881;
w4883 <= w4594 and not w4882;
w4884 <= not w4594 and w4882;
w4885 <= not w4883 and not w4884;
w4886 <= a(7) and a(39);
w4887 <= a(8) and a(38);
w4888 <= not w4886 and not w4887;
w4889 <= a(38) and a(39);
w4890 <= w186 and w4889;
w4891 <= w3312 and not w4890;
w4892 <= not w4888 and w4891;
w4893 <= w3312 and not w4892;
w4894 <= not w4890 and not w4892;
w4895 <= not w4888 and w4894;
w4896 <= not w4893 and not w4895;
w4897 <= not w4885 and not w4896;
w4898 <= w4885 and w4896;
w4899 <= not w4897 and not w4898;
w4900 <= not w4869 and not w4899;
w4901 <= w4869 and w4899;
w4902 <= not w4900 and not w4901;
w4903 <= not w4820 and not w4902;
w4904 <= w4820 and w4902;
w4905 <= not w4903 and not w4904;
w4906 <= not w4819 and w4905;
w4907 <= w4819 and not w4905;
w4908 <= not w4906 and not w4907;
w4909 <= not w4686 and not w4690;
w4910 <= not w4642 and not w4656;
w4911 <= w4909 and w4910;
w4912 <= not w4909 and not w4910;
w4913 <= not w4911 and not w4912;
w4914 <= not w4579 and not w4597;
w4915 <= not w4913 and w4914;
w4916 <= w4913 and not w4914;
w4917 <= not w4915 and not w4916;
w4918 <= not w4550 and not w4601;
w4919 <= w4621 and w4668;
w4920 <= not w4621 and not w4668;
w4921 <= not w4919 and not w4920;
w4922 <= w4639 and not w4921;
w4923 <= not w4639 and w4921;
w4924 <= not w4922 and not w4923;
w4925 <= not w4543 and not w4546;
w4926 <= a(1) and a(45);
w4927 <= w1921 and w4926;
w4928 <= not w1921 and not w4926;
w4929 <= not w4927 and not w4928;
w4930 <= w4583 and w4929;
w4931 <= w4583 and not w4930;
w4932 <= not w4583 and w4929;
w4933 <= not w4931 and not w4932;
w4934 <= not w4653 and not w4933;
w4935 <= w4653 and not w4932;
w4936 <= not w4931 and w4935;
w4937 <= not w4934 and not w4936;
w4938 <= not w4925 and w4937;
w4939 <= w4925 and not w4937;
w4940 <= not w4938 and not w4939;
w4941 <= w4924 and w4940;
w4942 <= not w4924 and not w4940;
w4943 <= not w4941 and not w4942;
w4944 <= not w4918 and w4943;
w4945 <= w4918 and not w4943;
w4946 <= not w4944 and not w4945;
w4947 <= w4917 and w4946;
w4948 <= not w4917 and not w4946;
w4949 <= not w4947 and not w4948;
w4950 <= w4908 and w4949;
w4951 <= not w4908 and not w4949;
w4952 <= not w4950 and not w4951;
w4953 <= not w4817 and not w4952;
w4954 <= w4817 and w4952;
w4955 <= not w4953 and not w4954;
w4956 <= not w4748 and not w4751;
w4957 <= not w4747 and not w4956;
w4958 <= not w4955 and w4957;
w4959 <= w4955 and not w4957;
w4960 <= not w4958 and not w4959;
w4961 <= not w4812 and not w4816;
w4962 <= not w4760 and not w4809;
w4963 <= not w4944 and not w4947;
w4964 <= w4962 and w4963;
w4965 <= not w4962 and not w4963;
w4966 <= not w4964 and not w4965;
w4967 <= w4770 and w4860;
w4968 <= not w4770 and not w4860;
w4969 <= not w4967 and not w4968;
w4970 <= w4831 and not w4969;
w4971 <= not w4831 and w4969;
w4972 <= not w4970 and not w4971;
w4973 <= not w4849 and not w4866;
w4974 <= not w4972 and w4973;
w4975 <= w4972 and not w4973;
w4976 <= not w4974 and not w4975;
w4977 <= not w4788 and not w4794;
w4978 <= not w4976 and w4977;
w4979 <= w4976 and not w4977;
w4980 <= not w4978 and not w4979;
w4981 <= not w4869 and w4899;
w4982 <= not w4903 and not w4981;
w4983 <= not w4804 and not w4806;
w4984 <= not w4982 and not w4983;
w4985 <= not w4982 and not w4984;
w4986 <= not w4983 and not w4984;
w4987 <= not w4985 and not w4986;
w4988 <= w4980 and not w4987;
w4989 <= not w4980 and w4987;
w4990 <= w4966 and not w4989;
w4991 <= not w4988 and w4990;
w4992 <= w4966 and not w4991;
w4993 <= not w4989 and not w4991;
w4994 <= not w4988 and w4993;
w4995 <= not w4992 and not w4994;
w4996 <= not w4906 and not w4950;
w4997 <= not w4930 and not w4934;
w4998 <= a(12) and a(40);
w4999 <= w3939 and w4998;
w5000 <= w554 and w3125;
w5001 <= a(34) and a(40);
w5002 <= w901 and w5001;
w5003 <= not w5000 and not w5002;
w5004 <= not w4999 and not w5003;
w5005 <= a(34) and not w5004;
w5006 <= a(13) and w5005;
w5007 <= not w4999 and not w5004;
w5008 <= a(7) and a(40);
w5009 <= a(12) and a(35);
w5010 <= not w5008 and not w5009;
w5011 <= w5007 and not w5010;
w5012 <= not w5006 and not w5011;
w5013 <= not w4997 and not w5012;
w5014 <= not w4997 and not w5013;
w5015 <= not w5012 and not w5013;
w5016 <= not w5014 and not w5015;
w5017 <= not w4797 and not w4800;
w5018 <= w5016 and w5017;
w5019 <= not w5016 and not w5017;
w5020 <= not w5018 and not w5019;
w5021 <= not w4938 and not w4941;
w5022 <= not w5020 and w5021;
w5023 <= w5020 and not w5021;
w5024 <= not w5022 and not w5023;
w5025 <= not w4912 and not w4916;
w5026 <= not w5024 and w5025;
w5027 <= w5024 and not w5025;
w5028 <= not w5026 and not w5027;
w5029 <= not w4594 and not w4882;
w5030 <= not w4897 and not w5029;
w5031 <= not w4920 and not w4923;
w5032 <= w5030 and w5031;
w5033 <= not w5030 and not w5031;
w5034 <= not w5032 and not w5033;
w5035 <= a(1) and a(46);
w5036 <= not a(24) and not w5035;
w5037 <= a(24) and a(46);
w5038 <= a(1) and w5037;
w5039 <= not w4844 and not w5038;
w5040 <= not w5036 and w5039;
w5041 <= not w4844 and not w5040;
w5042 <= not w5038 and not w5040;
w5043 <= not w5036 and w5042;
w5044 <= not w5041 and not w5043;
w5045 <= not w4894 and not w5044;
w5046 <= not w4894 and not w5045;
w5047 <= not w5044 and not w5045;
w5048 <= not w5046 and not w5047;
w5049 <= w5034 and not w5048;
w5050 <= w5034 and not w5049;
w5051 <= not w5048 and not w5049;
w5052 <= not w5050 and not w5051;
w5053 <= a(0) and a(47);
w5054 <= a(2) and a(45);
w5055 <= not w5053 and not w5054;
w5056 <= a(45) and a(47);
w5057 <= w2 and w5056;
w5058 <= not w5055 and not w5057;
w5059 <= w4927 and w5058;
w5060 <= not w5057 and not w5059;
w5061 <= not w5055 and w5060;
w5062 <= w4927 and not w5059;
w5063 <= not w5061 and not w5062;
w5064 <= w858 and w2423;
w5065 <= w856 and w3258;
w5066 <= w854 and w2671;
w5067 <= not w5065 and not w5066;
w5068 <= not w5064 and not w5067;
w5069 <= a(31) and not w5068;
w5070 <= a(16) and w5069;
w5071 <= not w5064 and not w5068;
w5072 <= a(17) and a(30);
w5073 <= a(18) and a(29);
w5074 <= not w5072 and not w5073;
w5075 <= w5071 and not w5074;
w5076 <= not w5070 and not w5075;
w5077 <= not w5063 and not w5076;
w5078 <= not w5063 and not w5077;
w5079 <= not w5076 and not w5077;
w5080 <= not w5078 and not w5079;
w5081 <= w1300 and w2033;
w5082 <= w1298 and w2606;
w5083 <= w1296 and w2137;
w5084 <= not w5082 and not w5083;
w5085 <= not w5081 and not w5084;
w5086 <= a(28) and not w5085;
w5087 <= a(19) and w5086;
w5088 <= not w5081 and not w5085;
w5089 <= a(20) and a(27);
w5090 <= not w1893 and not w5089;
w5091 <= w5088 and not w5090;
w5092 <= not w5087 and not w5091;
w5093 <= not w5080 and not w5092;
w5094 <= not w5080 and not w5093;
w5095 <= not w5092 and not w5093;
w5096 <= not w5094 and not w5095;
w5097 <= w4784 and w4877;
w5098 <= not w4784 and not w4877;
w5099 <= not w5097 and not w5098;
w5100 <= a(32) and a(43);
w5101 <= w808 and w5100;
w5102 <= a(43) and a(44);
w5103 <= w15 and w5102;
w5104 <= a(15) and a(44);
w5105 <= w2786 and w5104;
w5106 <= not w5103 and not w5105;
w5107 <= not w5101 and not w5106;
w5108 <= a(44) and not w5107;
w5109 <= a(3) and w5108;
w5110 <= not w5101 and not w5107;
w5111 <= a(15) and a(32);
w5112 <= not w4169 and not w5111;
w5113 <= w5110 and not w5112;
w5114 <= not w5109 and not w5113;
w5115 <= w5099 and not w5114;
w5116 <= w5099 and not w5115;
w5117 <= not w5114 and not w5115;
w5118 <= not w5116 and not w5117;
w5119 <= w882 and w3336;
w5120 <= w238 and w4889;
w5121 <= a(11) and a(39);
w5122 <= w4399 and w5121;
w5123 <= not w5120 and not w5122;
w5124 <= not w5119 and not w5123;
w5125 <= not w5119 and not w5124;
w5126 <= a(9) and a(38);
w5127 <= a(11) and a(36);
w5128 <= not w5126 and not w5127;
w5129 <= w5125 and not w5128;
w5130 <= a(39) and not w5124;
w5131 <= a(8) and w5130;
w5132 <= not w5129 and not w5131;
w5133 <= a(22) and a(25);
w5134 <= not w1472 and not w5133;
w5135 <= w1710 and w1725;
w5136 <= a(37) and not w5135;
w5137 <= a(10) and w5136;
w5138 <= not w5134 and w5137;
w5139 <= a(37) and not w5138;
w5140 <= a(10) and w5139;
w5141 <= not w5135 and not w5138;
w5142 <= not w5134 and w5141;
w5143 <= not w5140 and not w5142;
w5144 <= not w5132 and not w5143;
w5145 <= not w5132 and not w5144;
w5146 <= not w5143 and not w5144;
w5147 <= not w5145 and not w5146;
w5148 <= a(33) and a(41);
w5149 <= w921 and w5148;
w5150 <= a(41) and a(42);
w5151 <= w138 and w5150;
w5152 <= a(14) and a(42);
w5153 <= w3229 and w5152;
w5154 <= not w5151 and not w5153;
w5155 <= not w5149 and not w5154;
w5156 <= a(42) and not w5155;
w5157 <= a(5) and w5156;
w5158 <= a(6) and a(41);
w5159 <= a(14) and a(33);
w5160 <= not w5158 and not w5159;
w5161 <= not w5149 and not w5155;
w5162 <= not w5160 and w5161;
w5163 <= not w5157 and not w5162;
w5164 <= not w5147 and not w5163;
w5165 <= not w5147 and not w5164;
w5166 <= not w5163 and not w5164;
w5167 <= not w5165 and not w5166;
w5168 <= not w5118 and w5167;
w5169 <= w5118 and not w5167;
w5170 <= not w5168 and not w5169;
w5171 <= not w5096 and not w5170;
w5172 <= w5096 and w5170;
w5173 <= not w5171 and not w5172;
w5174 <= not w5052 and w5173;
w5175 <= not w5052 and not w5174;
w5176 <= w5173 and not w5174;
w5177 <= not w5175 and not w5176;
w5178 <= w5028 and not w5177;
w5179 <= not w5028 and not w5176;
w5180 <= not w5175 and w5179;
w5181 <= not w5178 and not w5180;
w5182 <= not w4996 and w5181;
w5183 <= not w4996 and not w5182;
w5184 <= w5181 and not w5182;
w5185 <= not w5183 and not w5184;
w5186 <= not w4995 and not w5185;
w5187 <= w4995 and not w5184;
w5188 <= not w5183 and w5187;
w5189 <= not w5186 and not w5188;
w5190 <= not w4961 and w5189;
w5191 <= w4961 and not w5189;
w5192 <= not w5190 and not w5191;
w5193 <= not w4953 and not w4957;
w5194 <= not w4954 and not w5193;
w5195 <= not w5192 and w5194;
w5196 <= w5192 and not w5194;
w5197 <= not w5195 and not w5196;
w5198 <= not w5191 and not w5194;
w5199 <= not w5190 and not w5198;
w5200 <= not w5182 and not w5186;
w5201 <= not w4965 and not w4991;
w5202 <= not w4984 and not w4988;
w5203 <= not w5023 and not w5027;
w5204 <= w551 and w3125;
w5205 <= w3688 and w5152;
w5206 <= not w5204 and not w5205;
w5207 <= a(6) and a(42);
w5208 <= a(13) and a(35);
w5209 <= w5207 and w5208;
w5210 <= not w5206 and not w5209;
w5211 <= not w5209 and not w5210;
w5212 <= not w5207 and not w5208;
w5213 <= w5211 and not w5212;
w5214 <= a(34) and not w5210;
w5215 <= a(14) and w5214;
w5216 <= not w5213 and not w5215;
w5217 <= a(7) and a(41);
w5218 <= w4399 and w4998;
w5219 <= a(40) and a(41);
w5220 <= w186 and w5219;
w5221 <= w3636 and w5217;
w5222 <= not w5220 and not w5221;
w5223 <= not w5218 and not w5222;
w5224 <= w5217 and not w5223;
w5225 <= a(8) and a(40);
w5226 <= not w3636 and not w5225;
w5227 <= not w5218 and not w5223;
w5228 <= not w5226 and w5227;
w5229 <= not w5224 and not w5228;
w5230 <= not w5216 and not w5229;
w5231 <= not w5216 and not w5230;
w5232 <= not w5229 and not w5230;
w5233 <= not w5231 and not w5232;
w5234 <= a(9) and a(39);
w5235 <= w529 and w4371;
w5236 <= a(37) and a(39);
w5237 <= w882 and w5236;
w5238 <= w290 and w4889;
w5239 <= not w5237 and not w5238;
w5240 <= not w5235 and not w5239;
w5241 <= w5234 and not w5240;
w5242 <= not w5235 and not w5240;
w5243 <= a(10) and a(38);
w5244 <= not w4367 and not w5243;
w5245 <= w5242 and not w5244;
w5246 <= not w5241 and not w5245;
w5247 <= not w5233 and not w5246;
w5248 <= not w5233 and not w5247;
w5249 <= not w5246 and not w5247;
w5250 <= not w5248 and not w5249;
w5251 <= not w5013 and not w5019;
w5252 <= w5250 and w5251;
w5253 <= not w5250 and not w5251;
w5254 <= not w5252 and not w5253;
w5255 <= a(33) and a(43);
w5256 <= w920 and w5255;
w5257 <= a(33) and a(44);
w5258 <= w808 and w5257;
w5259 <= w32 and w5102;
w5260 <= not w5258 and not w5259;
w5261 <= not w5256 and not w5260;
w5262 <= not w5256 and not w5261;
w5263 <= a(5) and a(43);
w5264 <= a(15) and a(33);
w5265 <= not w5263 and not w5264;
w5266 <= w5262 and not w5265;
w5267 <= a(44) and not w5261;
w5268 <= a(4) and w5267;
w5269 <= not w5266 and not w5268;
w5270 <= w1380 and w2033;
w5271 <= w1499 and w2606;
w5272 <= w1300 and w2137;
w5273 <= not w5271 and not w5272;
w5274 <= not w5270 and not w5273;
w5275 <= a(28) and not w5274;
w5276 <= a(20) and w5275;
w5277 <= a(21) and a(27);
w5278 <= a(22) and a(26);
w5279 <= not w5277 and not w5278;
w5280 <= not w5270 and not w5274;
w5281 <= not w5279 and w5280;
w5282 <= not w5276 and not w5281;
w5283 <= not w5269 and not w5282;
w5284 <= not w5269 and not w5283;
w5285 <= not w5282 and not w5283;
w5286 <= not w5284 and not w5285;
w5287 <= w955 and w2423;
w5288 <= w2940 and w3258;
w5289 <= w858 and w2671;
w5290 <= not w5288 and not w5289;
w5291 <= not w5287 and not w5290;
w5292 <= a(31) and not w5291;
w5293 <= a(17) and w5292;
w5294 <= not w5287 and not w5291;
w5295 <= a(18) and a(30);
w5296 <= a(19) and a(29);
w5297 <= not w5295 and not w5296;
w5298 <= w5294 and not w5297;
w5299 <= not w5293 and not w5298;
w5300 <= not w5286 and not w5299;
w5301 <= not w5286 and not w5300;
w5302 <= not w5299 and not w5300;
w5303 <= not w5301 and not w5302;
w5304 <= not w5254 and w5303;
w5305 <= w5254 and not w5303;
w5306 <= not w5304 and not w5305;
w5307 <= not w5203 and w5306;
w5308 <= w5203 and not w5306;
w5309 <= not w5307 and not w5308;
w5310 <= not w5202 and w5309;
w5311 <= w5202 and not w5309;
w5312 <= not w5310 and not w5311;
w5313 <= w5201 and not w5312;
w5314 <= not w5201 and w5312;
w5315 <= not w5313 and not w5314;
w5316 <= not w5174 and not w5178;
w5317 <= not w4975 and not w4979;
w5318 <= not w5033 and not w5049;
w5319 <= w5317 and w5318;
w5320 <= not w5317 and not w5318;
w5321 <= not w5319 and not w5320;
w5322 <= a(0) and a(48);
w5323 <= w5038 and w5322;
w5324 <= w5038 and not w5323;
w5325 <= not w5038 and w5322;
w5326 <= not w5324 and not w5325;
w5327 <= a(1) and a(47);
w5328 <= w1353 and w5327;
w5329 <= w5327 and not w5328;
w5330 <= w1353 and not w5328;
w5331 <= not w5329 and not w5330;
w5332 <= not w5326 and not w5331;
w5333 <= not w5326 and not w5332;
w5334 <= not w5331 and not w5332;
w5335 <= not w5333 and not w5334;
w5336 <= not w4968 and not w4971;
w5337 <= w5335 and w5336;
w5338 <= not w5335 and not w5336;
w5339 <= not w5337 and not w5338;
w5340 <= not w5098 and not w5115;
w5341 <= not w5339 and w5340;
w5342 <= w5339 and not w5340;
w5343 <= not w5341 and not w5342;
w5344 <= w5321 and w5343;
w5345 <= not w5321 and not w5343;
w5346 <= not w5344 and not w5345;
w5347 <= not w5316 and w5346;
w5348 <= not w5316 and not w5347;
w5349 <= w5346 and not w5347;
w5350 <= not w5348 and not w5349;
w5351 <= w5088 and w5125;
w5352 <= not w5088 and not w5125;
w5353 <= not w5351 and not w5352;
w5354 <= w5161 and not w5353;
w5355 <= not w5161 and w5353;
w5356 <= not w5354 and not w5355;
w5357 <= not w5144 and not w5164;
w5358 <= not w5356 and w5357;
w5359 <= w5356 and not w5357;
w5360 <= not w5358 and not w5359;
w5361 <= w5007 and w5141;
w5362 <= not w5007 and not w5141;
w5363 <= not w5361 and not w5362;
w5364 <= a(32) and a(46);
w5365 <= w708 and w5364;
w5366 <= a(45) and a(46);
w5367 <= w24 and w5366;
w5368 <= not w5365 and not w5367;
w5369 <= a(3) and a(45);
w5370 <= a(16) and a(32);
w5371 <= w5369 and w5370;
w5372 <= not w5368 and not w5371;
w5373 <= a(46) and not w5372;
w5374 <= a(2) and w5373;
w5375 <= not w5371 and not w5372;
w5376 <= not w5369 and not w5370;
w5377 <= w5375 and not w5376;
w5378 <= not w5374 and not w5377;
w5379 <= w5363 and not w5378;
w5380 <= w5363 and not w5379;
w5381 <= not w5378 and not w5379;
w5382 <= not w5380 and not w5381;
w5383 <= not w5360 and w5382;
w5384 <= w5360 and not w5382;
w5385 <= not w5383 and not w5384;
w5386 <= not w5118 and not w5167;
w5387 <= not w5171 and not w5386;
w5388 <= w5385 and not w5387;
w5389 <= not w5385 and w5387;
w5390 <= not w5388 and not w5389;
w5391 <= w5071 and w5110;
w5392 <= not w5071 and not w5110;
w5393 <= not w5391 and not w5392;
w5394 <= w5060 and not w5393;
w5395 <= not w5060 and w5393;
w5396 <= not w5394 and not w5395;
w5397 <= not w5040 and not w5045;
w5398 <= not w5077 and not w5093;
w5399 <= w5397 and w5398;
w5400 <= not w5397 and not w5398;
w5401 <= not w5399 and not w5400;
w5402 <= w5396 and w5401;
w5403 <= not w5396 and not w5401;
w5404 <= not w5402 and not w5403;
w5405 <= w5390 and w5404;
w5406 <= not w5390 and not w5404;
w5407 <= not w5405 and not w5406;
w5408 <= not w5350 and w5407;
w5409 <= not w5349 and not w5407;
w5410 <= not w5348 and w5409;
w5411 <= not w5408 and not w5410;
w5412 <= w5315 and w5411;
w5413 <= not w5315 and not w5411;
w5414 <= not w5412 and not w5413;
w5415 <= w5200 and not w5414;
w5416 <= not w5200 and w5414;
w5417 <= not w5415 and not w5416;
w5418 <= w5199 and not w5417;
w5419 <= not w5199 and not w5415;
w5420 <= not w5416 and w5419;
w5421 <= not w5418 and not w5420;
w5422 <= not w5347 and not w5408;
w5423 <= not w5388 and not w5405;
w5424 <= not w5320 and not w5344;
w5425 <= a(7) and a(42);
w5426 <= a(8) and a(41);
w5427 <= not w5425 and not w5426;
w5428 <= w186 and w5150;
w5429 <= a(36) and not w5428;
w5430 <= a(13) and w5429;
w5431 <= not w5427 and w5430;
w5432 <= not w5428 and not w5431;
w5433 <= not w5427 and w5432;
w5434 <= a(36) and not w5431;
w5435 <= a(13) and w5434;
w5436 <= not w5433 and not w5435;
w5437 <= not w1710 and not w2109;
w5438 <= w1710 and w2109;
w5439 <= a(38) and not w5438;
w5440 <= a(11) and w5439;
w5441 <= not w5437 and w5440;
w5442 <= a(38) and not w5441;
w5443 <= a(11) and w5442;
w5444 <= not w5438 and not w5441;
w5445 <= not w5437 and w5444;
w5446 <= not w5443 and not w5445;
w5447 <= not w5436 and not w5446;
w5448 <= not w5436 and not w5447;
w5449 <= not w5446 and not w5447;
w5450 <= not w5448 and not w5449;
w5451 <= a(35) and a(43);
w5452 <= w921 and w5451;
w5453 <= a(15) and a(43);
w5454 <= w3688 and w5453;
w5455 <= w701 and w3125;
w5456 <= not w5454 and not w5455;
w5457 <= not w5452 and not w5456;
w5458 <= a(34) and not w5457;
w5459 <= a(15) and w5458;
w5460 <= a(6) and a(43);
w5461 <= a(14) and a(35);
w5462 <= not w5460 and not w5461;
w5463 <= not w5452 and not w5457;
w5464 <= not w5462 and w5463;
w5465 <= not w5459 and not w5464;
w5466 <= not w5450 and not w5465;
w5467 <= not w5450 and not w5466;
w5468 <= not w5465 and not w5466;
w5469 <= not w5467 and not w5468;
w5470 <= a(2) and a(47);
w5471 <= not w4826 and not w5470;
w5472 <= a(46) and a(47);
w5473 <= w24 and w5472;
w5474 <= a(27) and not w5473;
w5475 <= a(22) and w5474;
w5476 <= not w5471 and w5475;
w5477 <= not w5473 and not w5476;
w5478 <= not w5471 and w5477;
w5479 <= a(27) and not w5476;
w5480 <= a(22) and w5479;
w5481 <= not w5478 and not w5480;
w5482 <= w1300 and w2140;
w5483 <= w1298 and w2916;
w5484 <= w1296 and w2423;
w5485 <= not w5483 and not w5484;
w5486 <= not w5482 and not w5485;
w5487 <= a(30) and not w5486;
w5488 <= a(19) and w5487;
w5489 <= not w5482 and not w5486;
w5490 <= a(20) and a(29);
w5491 <= a(21) and a(28);
w5492 <= not w5490 and not w5491;
w5493 <= w5489 and not w5492;
w5494 <= not w5488 and not w5493;
w5495 <= not w5481 and not w5494;
w5496 <= not w5481 and not w5495;
w5497 <= not w5494 and not w5495;
w5498 <= not w5496 and not w5497;
w5499 <= w286 and w5236;
w5500 <= w290 and w3977;
w5501 <= a(37) and a(40);
w5502 <= w988 and w5501;
w5503 <= not w5500 and not w5502;
w5504 <= not w5499 and not w5503;
w5505 <= a(40) and not w5504;
w5506 <= a(9) and w5505;
w5507 <= not w5499 and not w5504;
w5508 <= a(10) and a(39);
w5509 <= not w4291 and not w5508;
w5510 <= w5507 and not w5509;
w5511 <= not w5506 and not w5510;
w5512 <= not w5498 and not w5511;
w5513 <= not w5498 and not w5512;
w5514 <= not w5511 and not w5512;
w5515 <= not w5513 and not w5514;
w5516 <= a(44) and w30;
w5517 <= a(45) and w18;
w5518 <= not w5516 and not w5517;
w5519 <= a(44) and a(45);
w5520 <= w32 and w5519;
w5521 <= a(49) and not w5520;
w5522 <= not w5518 and w5521;
w5523 <= a(0) and not w5522;
w5524 <= a(49) and w5523;
w5525 <= not w5520 and not w5522;
w5526 <= a(4) and a(45);
w5527 <= a(5) and a(44);
w5528 <= not w5526 and not w5527;
w5529 <= w5525 and not w5528;
w5530 <= not w5524 and not w5529;
w5531 <= not w5323 and not w5332;
w5532 <= not w5530 and w5531;
w5533 <= w5530 and not w5531;
w5534 <= not w5532 and not w5533;
w5535 <= w858 and w3618;
w5536 <= w856 and w2404;
w5537 <= w854 and w2949;
w5538 <= not w5536 and not w5537;
w5539 <= not w5535 and not w5538;
w5540 <= a(33) and not w5539;
w5541 <= a(16) and w5540;
w5542 <= not w5535 and not w5539;
w5543 <= a(17) and a(32);
w5544 <= a(18) and a(31);
w5545 <= not w5543 and not w5544;
w5546 <= w5542 and not w5545;
w5547 <= not w5541 and not w5546;
w5548 <= not w5534 and not w5547;
w5549 <= w5534 and w5547;
w5550 <= not w5548 and not w5549;
w5551 <= w5515 and w5550;
w5552 <= not w5515 and not w5550;
w5553 <= not w5551 and not w5552;
w5554 <= not w5469 and not w5553;
w5555 <= w5469 and w5553;
w5556 <= not w5554 and not w5555;
w5557 <= not w5424 and w5556;
w5558 <= w5424 and not w5556;
w5559 <= not w5557 and not w5558;
w5560 <= not w5423 and w5559;
w5561 <= w5423 and not w5559;
w5562 <= not w5560 and not w5561;
w5563 <= not w5422 and w5562;
w5564 <= w5422 and not w5562;
w5565 <= not w5563 and not w5564;
w5566 <= not w5307 and not w5310;
w5567 <= not w5352 and not w5355;
w5568 <= not w5362 and not w5379;
w5569 <= w5567 and w5568;
w5570 <= not w5567 and not w5568;
w5571 <= not w5569 and not w5570;
w5572 <= not w5392 and not w5395;
w5573 <= not w5571 and w5572;
w5574 <= w5571 and not w5572;
w5575 <= not w5573 and not w5574;
w5576 <= not w5359 and not w5384;
w5577 <= not w5400 and not w5402;
w5578 <= not w5576 and not w5577;
w5579 <= not w5576 and not w5578;
w5580 <= not w5577 and not w5578;
w5581 <= not w5579 and not w5580;
w5582 <= not w5575 and w5581;
w5583 <= w5575 and not w5581;
w5584 <= not w5582 and not w5583;
w5585 <= not w5566 and w5584;
w5586 <= not w5566 and not w5585;
w5587 <= w5584 and not w5585;
w5588 <= not w5586 and not w5587;
w5589 <= w5211 and w5294;
w5590 <= not w5211 and not w5294;
w5591 <= not w5589 and not w5590;
w5592 <= w5227 and not w5591;
w5593 <= not w5227 and w5591;
w5594 <= not w5592 and not w5593;
w5595 <= not w5283 and not w5300;
w5596 <= not w5594 and w5595;
w5597 <= w5594 and not w5595;
w5598 <= not w5596 and not w5597;
w5599 <= not w5338 and not w5342;
w5600 <= not w5598 and w5599;
w5601 <= w5598 and not w5599;
w5602 <= not w5600 and not w5601;
w5603 <= not w5253 and not w5305;
w5604 <= w5602 and not w5603;
w5605 <= not w5602 and w5603;
w5606 <= not w5604 and not w5605;
w5607 <= w5262 and w5375;
w5608 <= not w5262 and not w5375;
w5609 <= not w5607 and not w5608;
w5610 <= w5280 and not w5609;
w5611 <= not w5280 and w5609;
w5612 <= not w5610 and not w5611;
w5613 <= not w5230 and not w5247;
w5614 <= a(48) and w1553;
w5615 <= a(1) and a(48);
w5616 <= not a(25) and not w5615;
w5617 <= not w5614 and not w5616;
w5618 <= w5328 and w5617;
w5619 <= not w5328 and not w5617;
w5620 <= not w5618 and not w5619;
w5621 <= not w5242 and w5620;
w5622 <= w5242 and not w5620;
w5623 <= not w5621 and not w5622;
w5624 <= not w5613 and w5623;
w5625 <= w5613 and not w5623;
w5626 <= not w5624 and not w5625;
w5627 <= w5612 and w5626;
w5628 <= not w5612 and not w5626;
w5629 <= not w5627 and not w5628;
w5630 <= w5606 and w5629;
w5631 <= not w5606 and not w5629;
w5632 <= not w5630 and not w5631;
w5633 <= not w5588 and w5632;
w5634 <= not w5587 and not w5632;
w5635 <= not w5586 and w5634;
w5636 <= not w5633 and not w5635;
w5637 <= w5565 and w5636;
w5638 <= not w5565 and not w5636;
w5639 <= not w5637 and not w5638;
w5640 <= not w5314 and not w5412;
w5641 <= not w5639 and w5640;
w5642 <= w5639 and not w5640;
w5643 <= not w5641 and not w5642;
w5644 <= not w5416 and not w5419;
w5645 <= not w5643 and w5644;
w5646 <= w5643 and not w5644;
w5647 <= not w5645 and not w5646;
w5648 <= not w5641 and not w5644;
w5649 <= not w5642 and not w5648;
w5650 <= not w5563 and not w5637;
w5651 <= not w5585 and not w5633;
w5652 <= not w5604 and not w5630;
w5653 <= not w5578 and not w5583;
w5654 <= a(35) and a(45);
w5655 <= w920 and w5654;
w5656 <= a(16) and a(45);
w5657 <= w3470 and w5656;
w5658 <= w697 and w3125;
w5659 <= not w5657 and not w5658;
w5660 <= not w5655 and not w5659;
w5661 <= not w5655 and not w5660;
w5662 <= a(5) and a(45);
w5663 <= a(15) and a(35);
w5664 <= not w5662 and not w5663;
w5665 <= w5661 and not w5664;
w5666 <= a(34) and not w5660;
w5667 <= a(16) and w5666;
w5668 <= not w5665 and not w5667;
w5669 <= a(28) and a(32);
w5670 <= w1275 and w5669;
w5671 <= w1725 and w2137;
w5672 <= not w5670 and not w5671;
w5673 <= a(18) and a(32);
w5674 <= a(23) and a(27);
w5675 <= w5673 and w5674;
w5676 <= not w5672 and not w5675;
w5677 <= a(28) and not w5676;
w5678 <= a(22) and w5677;
w5679 <= not w5673 and not w5674;
w5680 <= not w5675 and not w5676;
w5681 <= not w5679 and w5680;
w5682 <= not w5678 and not w5681;
w5683 <= not w5668 and not w5682;
w5684 <= not w5668 and not w5683;
w5685 <= not w5682 and not w5683;
w5686 <= not w5684 and not w5685;
w5687 <= not w5618 and not w5621;
w5688 <= w5686 and w5687;
w5689 <= not w5686 and not w5687;
w5690 <= not w5688 and not w5689;
w5691 <= a(0) and a(50);
w5692 <= a(2) and a(48);
w5693 <= not w5691 and not w5692;
w5694 <= a(48) and a(50);
w5695 <= w2 and w5694;
w5696 <= not w5693 and not w5695;
w5697 <= w5614 and w5696;
w5698 <= not w5695 and not w5697;
w5699 <= not w5693 and w5698;
w5700 <= w5614 and not w5697;
w5701 <= not w5699 and not w5700;
w5702 <= a(33) and a(46);
w5703 <= w987 and w5702;
w5704 <= w15 and w5472;
w5705 <= a(17) and a(47);
w5706 <= w2952 and w5705;
w5707 <= not w5704 and not w5706;
w5708 <= not w5703 and not w5707;
w5709 <= a(47) and not w5708;
w5710 <= a(3) and w5709;
w5711 <= not w5703 and not w5708;
w5712 <= a(4) and a(46);
w5713 <= a(17) and a(33);
w5714 <= not w5712 and not w5713;
w5715 <= w5711 and not w5714;
w5716 <= not w5710 and not w5715;
w5717 <= not w5701 and not w5716;
w5718 <= not w5701 and not w5717;
w5719 <= not w5716 and not w5717;
w5720 <= not w5718 and not w5719;
w5721 <= w1300 and w2423;
w5722 <= w1298 and w3258;
w5723 <= w1296 and w2671;
w5724 <= not w5722 and not w5723;
w5725 <= not w5721 and not w5724;
w5726 <= a(31) and not w5725;
w5727 <= a(19) and w5726;
w5728 <= not w5721 and not w5725;
w5729 <= a(20) and a(30);
w5730 <= a(21) and a(29);
w5731 <= not w5729 and not w5730;
w5732 <= w5728 and not w5731;
w5733 <= not w5727 and not w5732;
w5734 <= not w5720 and not w5733;
w5735 <= not w5720 and not w5734;
w5736 <= not w5733 and not w5734;
w5737 <= not w5735 and not w5736;
w5738 <= w141 and w5102;
w5739 <= a(36) and a(44);
w5740 <= w921 and w5739;
w5741 <= not w5738 and not w5740;
w5742 <= a(7) and a(43);
w5743 <= a(14) and a(36);
w5744 <= w5742 and w5743;
w5745 <= not w5741 and not w5744;
w5746 <= not w5744 and not w5745;
w5747 <= not w5742 and not w5743;
w5748 <= w5746 and not w5747;
w5749 <= a(44) and not w5745;
w5750 <= a(6) and w5749;
w5751 <= not w5748 and not w5750;
w5752 <= a(37) and a(41);
w5753 <= w332 and w5752;
w5754 <= w238 and w5150;
w5755 <= a(13) and a(42);
w5756 <= w4636 and w5755;
w5757 <= not w5754 and not w5756;
w5758 <= not w5753 and not w5757;
w5759 <= a(42) and not w5758;
w5760 <= a(8) and w5759;
w5761 <= not w5753 and not w5758;
w5762 <= a(9) and a(41);
w5763 <= not w3495 and not w5762;
w5764 <= w5761 and not w5763;
w5765 <= not w5760 and not w5764;
w5766 <= not w5751 and not w5765;
w5767 <= not w5751 and not w5766;
w5768 <= not w5765 and not w5766;
w5769 <= not w5767 and not w5768;
w5770 <= w529 and w3977;
w5771 <= w286 and w3609;
w5772 <= w408 and w4889;
w5773 <= not w5771 and not w5772;
w5774 <= not w5770 and not w5773;
w5775 <= a(38) and not w5774;
w5776 <= a(12) and w5775;
w5777 <= not w5770 and not w5774;
w5778 <= a(10) and a(40);
w5779 <= not w5121 and not w5778;
w5780 <= w5777 and not w5779;
w5781 <= not w5776 and not w5780;
w5782 <= not w5769 and not w5781;
w5783 <= not w5769 and not w5782;
w5784 <= not w5781 and not w5782;
w5785 <= not w5783 and not w5784;
w5786 <= not w5737 and w5785;
w5787 <= w5737 and not w5785;
w5788 <= not w5786 and not w5787;
w5789 <= w5690 and not w5788;
w5790 <= not w5690 and w5788;
w5791 <= not w5789 and not w5790;
w5792 <= not w5653 and w5791;
w5793 <= not w5653 and not w5792;
w5794 <= w5791 and not w5792;
w5795 <= not w5793 and not w5794;
w5796 <= not w5652 and not w5795;
w5797 <= w5652 and not w5794;
w5798 <= not w5793 and w5797;
w5799 <= not w5796 and not w5798;
w5800 <= not w5651 and w5799;
w5801 <= w5651 and not w5799;
w5802 <= not w5800 and not w5801;
w5803 <= not w5557 and not w5560;
w5804 <= not w5597 and not w5601;
w5805 <= not w5624 and not w5627;
w5806 <= w5804 and w5805;
w5807 <= not w5804 and not w5805;
w5808 <= not w5806 and not w5807;
w5809 <= not w5590 and not w5593;
w5810 <= not w5608 and not w5611;
w5811 <= w5809 and w5810;
w5812 <= not w5809 and not w5810;
w5813 <= not w5811 and not w5812;
w5814 <= w5477 and w5525;
w5815 <= not w5477 and not w5525;
w5816 <= not w5814 and not w5815;
w5817 <= w5463 and not w5816;
w5818 <= not w5463 and w5816;
w5819 <= not w5817 and not w5818;
w5820 <= w5813 and w5819;
w5821 <= not w5813 and not w5819;
w5822 <= not w5820 and not w5821;
w5823 <= w5808 and w5822;
w5824 <= not w5808 and not w5822;
w5825 <= not w5823 and not w5824;
w5826 <= w5803 and not w5825;
w5827 <= not w5803 and w5825;
w5828 <= not w5826 and not w5827;
w5829 <= not w5495 and not w5512;
w5830 <= not w5530 and not w5531;
w5831 <= not w5548 and not w5830;
w5832 <= w5829 and w5831;
w5833 <= not w5829 and not w5831;
w5834 <= not w5832 and not w5833;
w5835 <= a(1) and a(49);
w5836 <= w2107 and w5835;
w5837 <= not w2107 and not w5835;
w5838 <= not w5836 and not w5837;
w5839 <= w5444 and not w5838;
w5840 <= not w5444 and w5838;
w5841 <= not w5839 and not w5840;
w5842 <= not w5507 and w5841;
w5843 <= w5507 and not w5841;
w5844 <= not w5842 and not w5843;
w5845 <= w5834 and w5844;
w5846 <= not w5834 and not w5844;
w5847 <= not w5845 and not w5846;
w5848 <= w5489 and w5542;
w5849 <= not w5489 and not w5542;
w5850 <= not w5848 and not w5849;
w5851 <= w5432 and not w5850;
w5852 <= not w5432 and w5850;
w5853 <= not w5851 and not w5852;
w5854 <= not w5447 and not w5466;
w5855 <= not w5853 and w5854;
w5856 <= w5853 and not w5854;
w5857 <= not w5855 and not w5856;
w5858 <= not w5570 and not w5574;
w5859 <= not w5857 and w5858;
w5860 <= w5857 and not w5858;
w5861 <= not w5859 and not w5860;
w5862 <= not w5515 and w5550;
w5863 <= not w5554 and not w5862;
w5864 <= w5861 and not w5863;
w5865 <= not w5861 and w5863;
w5866 <= not w5864 and not w5865;
w5867 <= w5847 and w5866;
w5868 <= not w5847 and not w5866;
w5869 <= not w5867 and not w5868;
w5870 <= w5828 and w5869;
w5871 <= not w5828 and not w5869;
w5872 <= not w5870 and not w5871;
w5873 <= w5802 and w5872;
w5874 <= not w5802 and not w5872;
w5875 <= not w5873 and not w5874;
w5876 <= w5650 and not w5875;
w5877 <= not w5650 and w5875;
w5878 <= not w5876 and not w5877;
w5879 <= w5649 and not w5878;
w5880 <= not w5649 and not w5876;
w5881 <= not w5877 and w5880;
w5882 <= not w5879 and not w5881;
w5883 <= not w5877 and not w5880;
w5884 <= not w5800 and not w5873;
w5885 <= not w5827 and not w5870;
w5886 <= not w5864 and not w5867;
w5887 <= not w5807 and not w5823;
w5888 <= a(0) and a(51);
w5889 <= w5836 and w5888;
w5890 <= w5836 and not w5889;
w5891 <= not w5836 and w5888;
w5892 <= not w5890 and not w5891;
w5893 <= a(1) and a(50);
w5894 <= a(26) and w5893;
w5895 <= a(26) and not w5894;
w5896 <= w5893 and not w5894;
w5897 <= not w5895 and not w5896;
w5898 <= not w5892 and not w5897;
w5899 <= not w5892 and not w5898;
w5900 <= not w5897 and not w5898;
w5901 <= not w5899 and not w5900;
w5902 <= w1296 and w3618;
w5903 <= a(17) and not w5902;
w5904 <= a(20) and a(31);
w5905 <= a(19) and a(32);
w5906 <= not w5904 and not w5905;
w5907 <= a(34) and not w5906;
w5908 <= w5903 and w5907;
w5909 <= a(34) and not w5908;
w5910 <= a(17) and w5909;
w5911 <= not w5902 and not w5908;
w5912 <= not w5906 and w5911;
w5913 <= not w5910 and not w5912;
w5914 <= not w5901 and not w5913;
w5915 <= not w5901 and not w5914;
w5916 <= not w5913 and not w5914;
w5917 <= not w5915 and not w5916;
w5918 <= not w5849 and not w5852;
w5919 <= w5917 and w5918;
w5920 <= not w5917 and not w5918;
w5921 <= not w5919 and not w5920;
w5922 <= w1146 and w5702;
w5923 <= w856 and w2778;
w5924 <= not w5922 and not w5923;
w5925 <= a(5) and a(46);
w5926 <= a(16) and a(35);
w5927 <= w5925 and w5926;
w5928 <= not w5924 and not w5927;
w5929 <= not w5927 and not w5928;
w5930 <= not w5925 and not w5926;
w5931 <= w5929 and not w5930;
w5932 <= a(33) and not w5928;
w5933 <= a(18) and w5932;
w5934 <= not w5931 and not w5933;
w5935 <= w1725 and w2140;
w5936 <= w1173 and w2916;
w5937 <= w1380 and w2423;
w5938 <= not w5936 and not w5937;
w5939 <= not w5935 and not w5938;
w5940 <= a(30) and not w5939;
w5941 <= a(21) and w5940;
w5942 <= a(22) and a(29);
w5943 <= a(23) and a(28);
w5944 <= not w5942 and not w5943;
w5945 <= not w5935 and not w5939;
w5946 <= not w5944 and w5945;
w5947 <= not w5941 and not w5946;
w5948 <= not w5934 and not w5947;
w5949 <= not w5934 and not w5948;
w5950 <= not w5947 and not w5948;
w5951 <= not w5949 and not w5950;
w5952 <= a(37) and a(45);
w5953 <= w921 and w5952;
w5954 <= a(6) and a(45);
w5955 <= a(36) and w5954;
w5956 <= a(15) and w5955;
w5957 <= w701 and w3493;
w5958 <= not w5956 and not w5957;
w5959 <= not w5953 and not w5958;
w5960 <= a(36) and not w5959;
w5961 <= a(15) and w5960;
w5962 <= a(14) and a(37);
w5963 <= not w5954 and not w5962;
w5964 <= not w5953 and not w5959;
w5965 <= not w5963 and w5964;
w5966 <= not w5961 and not w5965;
w5967 <= not w5951 and not w5966;
w5968 <= not w5951 and not w5967;
w5969 <= not w5966 and not w5967;
w5970 <= not w5968 and not w5969;
w5971 <= a(13) and a(43);
w5972 <= w4887 and w5971;
w5973 <= w186 and w5102;
w5974 <= a(13) and a(44);
w5975 <= w4629 and w5974;
w5976 <= not w5973 and not w5975;
w5977 <= not w5972 and not w5976;
w5978 <= not w5972 and not w5977;
w5979 <= a(8) and a(43);
w5980 <= a(13) and a(38);
w5981 <= not w5979 and not w5980;
w5982 <= w5978 and not w5981;
w5983 <= a(44) and not w5977;
w5984 <= a(7) and w5983;
w5985 <= not w5982 and not w5984;
w5986 <= a(9) and a(42);
w5987 <= w286 and w3790;
w5988 <= w4556 and w5986;
w5989 <= w290 and w5150;
w5990 <= not w5988 and not w5989;
w5991 <= not w5987 and not w5990;
w5992 <= w5986 and not w5991;
w5993 <= not w5987 and not w5991;
w5994 <= a(10) and a(41);
w5995 <= not w4556 and not w5994;
w5996 <= w5993 and not w5995;
w5997 <= not w5992 and not w5996;
w5998 <= not w5985 and not w5997;
w5999 <= not w5985 and not w5998;
w6000 <= not w5997 and not w5998;
w6001 <= not w5999 and not w6000;
w6002 <= a(24) and a(27);
w6003 <= not w2269 and not w6002;
w6004 <= w1710 and w2033;
w6005 <= a(40) and not w6004;
w6006 <= a(11) and w6005;
w6007 <= not w6003 and w6006;
w6008 <= a(40) and not w6007;
w6009 <= a(11) and w6008;
w6010 <= not w6004 and not w6007;
w6011 <= not w6003 and w6010;
w6012 <= not w6009 and not w6011;
w6013 <= not w6001 and not w6012;
w6014 <= not w6001 and not w6013;
w6015 <= not w6012 and not w6013;
w6016 <= not w6014 and not w6015;
w6017 <= not w5970 and w6016;
w6018 <= w5970 and not w6016;
w6019 <= not w6017 and not w6018;
w6020 <= w5921 and not w6019;
w6021 <= not w5921 and w6019;
w6022 <= not w6020 and not w6021;
w6023 <= not w5887 and w6022;
w6024 <= w5887 and not w6022;
w6025 <= not w6023 and not w6024;
w6026 <= not w5886 and w6025;
w6027 <= w5886 and not w6025;
w6028 <= not w6026 and not w6027;
w6029 <= not w5885 and w6028;
w6030 <= w5885 and not w6028;
w6031 <= not w6029 and not w6030;
w6032 <= not w5792 and not w5796;
w6033 <= not w5856 and not w5860;
w6034 <= not w5833 and not w5845;
w6035 <= w6033 and w6034;
w6036 <= not w6033 and not w6034;
w6037 <= not w6035 and not w6036;
w6038 <= not w5815 and not w5818;
w6039 <= not w5840 and not w5842;
w6040 <= w6038 and w6039;
w6041 <= not w6038 and not w6039;
w6042 <= not w6040 and not w6041;
w6043 <= not w5717 and not w5734;
w6044 <= not w6042 and w6043;
w6045 <= w6042 and not w6043;
w6046 <= not w6044 and not w6045;
w6047 <= w6037 and w6046;
w6048 <= not w6037 and not w6046;
w6049 <= not w6047 and not w6048;
w6050 <= not w6032 and w6049;
w6051 <= w6032 and not w6049;
w6052 <= not w6050 and not w6051;
w6053 <= not w5737 and not w5785;
w6054 <= not w5789 and not w6053;
w6055 <= w5661 and w5777;
w6056 <= not w5661 and not w5777;
w6057 <= not w6055 and not w6056;
w6058 <= a(47) and a(48);
w6059 <= w15 and w6058;
w6060 <= a(47) and a(49);
w6061 <= w58 and w6060;
w6062 <= a(48) and a(49);
w6063 <= w24 and w6062;
w6064 <= not w6061 and not w6063;
w6065 <= not w6059 and not w6064;
w6066 <= a(49) and not w6065;
w6067 <= a(2) and w6066;
w6068 <= not w6059 and not w6065;
w6069 <= a(3) and a(48);
w6070 <= a(4) and a(47);
w6071 <= not w6069 and not w6070;
w6072 <= w6068 and not w6071;
w6073 <= not w6067 and not w6072;
w6074 <= w6057 and not w6073;
w6075 <= w6057 and not w6074;
w6076 <= not w6073 and not w6074;
w6077 <= not w6075 and not w6076;
w6078 <= not w5683 and not w5689;
w6079 <= w6077 and w6078;
w6080 <= not w6077 and not w6078;
w6081 <= not w6079 and not w6080;
w6082 <= not w5812 and not w5820;
w6083 <= w6081 and not w6082;
w6084 <= not w6081 and w6082;
w6085 <= not w6083 and not w6084;
w6086 <= not w6054 and w6085;
w6087 <= w6054 and not w6085;
w6088 <= not w6086 and not w6087;
w6089 <= w5746 and w5761;
w6090 <= not w5746 and not w5761;
w6091 <= not w6089 and not w6090;
w6092 <= w5680 and not w6091;
w6093 <= not w5680 and w6091;
w6094 <= not w6092 and not w6093;
w6095 <= not w5766 and not w5782;
w6096 <= not w6094 and w6095;
w6097 <= w6094 and not w6095;
w6098 <= not w6096 and not w6097;
w6099 <= w5711 and w5728;
w6100 <= not w5711 and not w5728;
w6101 <= not w6099 and not w6100;
w6102 <= w5698 and not w6101;
w6103 <= not w5698 and w6101;
w6104 <= not w6102 and not w6103;
w6105 <= w6098 and w6104;
w6106 <= not w6098 and not w6104;
w6107 <= not w6105 and not w6106;
w6108 <= w6088 and w6107;
w6109 <= not w6088 and not w6107;
w6110 <= not w6108 and not w6109;
w6111 <= w6052 and w6110;
w6112 <= not w6052 and not w6110;
w6113 <= not w6111 and not w6112;
w6114 <= w6031 and w6113;
w6115 <= not w6031 and not w6113;
w6116 <= not w6114 and not w6115;
w6117 <= not w5884 and w6116;
w6118 <= w5884 and not w6116;
w6119 <= not w6117 and not w6118;
w6120 <= not w5883 and not w6119;
w6121 <= w5883 and w6119;
w6122 <= not w6120 and not w6121;
w6123 <= not w5883 and not w6118;
w6124 <= not w6117 and not w6123;
w6125 <= not w6029 and not w6114;
w6126 <= not w6023 and not w6026;
w6127 <= not w6100 and not w6103;
w6128 <= a(2) and a(50);
w6129 <= a(3) and a(49);
w6130 <= not w6128 and not w6129;
w6131 <= a(49) and a(50);
w6132 <= w24 and w6131;
w6133 <= a(33) and not w6132;
w6134 <= a(19) and w6133;
w6135 <= not w6130 and w6134;
w6136 <= a(33) and not w6135;
w6137 <= a(19) and w6136;
w6138 <= not w6132 and not w6135;
w6139 <= not w6130 and w6138;
w6140 <= not w6137 and not w6139;
w6141 <= not w6127 and not w6140;
w6142 <= not w6127 and not w6141;
w6143 <= not w6140 and not w6141;
w6144 <= not w6142 and not w6143;
w6145 <= not w6090 and not w6093;
w6146 <= w6144 and w6145;
w6147 <= not w6144 and not w6145;
w6148 <= not w6146 and not w6147;
w6149 <= not w6080 and not w6083;
w6150 <= not w6148 and w6149;
w6151 <= w6148 and not w6149;
w6152 <= not w6150 and not w6151;
w6153 <= not w5998 and not w6013;
w6154 <= not w6056 and not w6074;
w6155 <= a(1) and a(51);
w6156 <= not w2439 and not w6155;
w6157 <= w2439 and w6155;
w6158 <= not w6156 and not w6157;
w6159 <= w5894 and w6158;
w6160 <= not w5894 and not w6158;
w6161 <= not w6159 and not w6160;
w6162 <= not w6010 and w6161;
w6163 <= w6010 and not w6161;
w6164 <= not w6162 and not w6163;
w6165 <= not w6154 and w6164;
w6166 <= w6154 and not w6164;
w6167 <= not w6165 and not w6166;
w6168 <= not w6153 and w6167;
w6169 <= w6153 and not w6167;
w6170 <= not w6168 and not w6169;
w6171 <= w6152 and w6170;
w6172 <= not w6152 and not w6170;
w6173 <= not w6171 and not w6172;
w6174 <= w6126 and not w6173;
w6175 <= not w6126 and w6173;
w6176 <= not w6174 and not w6175;
w6177 <= not w5889 and not w5898;
w6178 <= w5993 and w6177;
w6179 <= not w5993 and not w6177;
w6180 <= not w6178 and not w6179;
w6181 <= a(35) and w599;
w6182 <= a(48) and w18;
w6183 <= not w6181 and not w6182;
w6184 <= a(4) and a(48);
w6185 <= a(17) and a(35);
w6186 <= w6184 and w6185;
w6187 <= a(52) and not w6186;
w6188 <= not w6183 and w6187;
w6189 <= a(52) and not w6188;
w6190 <= a(0) and w6189;
w6191 <= not w6186 and not w6188;
w6192 <= not w6184 and not w6185;
w6193 <= w6191 and not w6192;
w6194 <= not w6190 and not w6193;
w6195 <= w6180 and not w6194;
w6196 <= w6180 and not w6195;
w6197 <= not w6194 and not w6195;
w6198 <= not w6196 and not w6197;
w6199 <= not w5914 and not w5920;
w6200 <= w6198 and w6199;
w6201 <= not w6198 and not w6199;
w6202 <= not w6200 and not w6201;
w6203 <= not w6041 and not w6045;
w6204 <= not w6202 and w6203;
w6205 <= w6202 and not w6203;
w6206 <= not w6204 and not w6205;
w6207 <= not w5970 and not w6016;
w6208 <= not w6020 and not w6207;
w6209 <= w5929 and w5978;
w6210 <= not w5929 and not w5978;
w6211 <= not w6209 and not w6210;
w6212 <= w5945 and not w6211;
w6213 <= not w5945 and w6211;
w6214 <= not w6212 and not w6213;
w6215 <= w5911 and w6068;
w6216 <= not w5911 and not w6068;
w6217 <= not w6215 and not w6216;
w6218 <= w5964 and not w6217;
w6219 <= not w5964 and w6217;
w6220 <= not w6218 and not w6219;
w6221 <= not w5948 and not w5967;
w6222 <= not w6220 and w6221;
w6223 <= w6220 and not w6221;
w6224 <= not w6222 and not w6223;
w6225 <= w6214 and w6224;
w6226 <= not w6214 and not w6224;
w6227 <= not w6225 and not w6226;
w6228 <= not w6208 and w6227;
w6229 <= not w6208 and not w6228;
w6230 <= w6227 and not w6228;
w6231 <= not w6229 and not w6230;
w6232 <= w6206 and not w6231;
w6233 <= w6206 and not w6232;
w6234 <= not w6231 and not w6232;
w6235 <= not w6233 and not w6234;
w6236 <= w6176 and not w6235;
w6237 <= w6176 and not w6236;
w6238 <= not w6235 and not w6236;
w6239 <= not w6237 and not w6238;
w6240 <= not w6086 and not w6108;
w6241 <= not w6036 and not w6047;
w6242 <= not w6097 and not w6105;
w6243 <= a(36) and a(46);
w6244 <= w527 and w6243;
w6245 <= w138 and w5472;
w6246 <= a(5) and a(47);
w6247 <= a(16) and a(36);
w6248 <= w6246 and w6247;
w6249 <= not w6245 and not w6248;
w6250 <= not w6244 and not w6249;
w6251 <= not w6244 and not w6250;
w6252 <= a(6) and a(46);
w6253 <= not w6247 and not w6252;
w6254 <= w6251 and not w6253;
w6255 <= w6246 and not w6250;
w6256 <= not w6254 and not w6255;
w6257 <= a(10) and a(42);
w6258 <= w408 and w5219;
w6259 <= a(40) and a(42);
w6260 <= w286 and w6259;
w6261 <= w529 and w5150;
w6262 <= not w6260 and not w6261;
w6263 <= not w6258 and not w6262;
w6264 <= w6257 and not w6263;
w6265 <= not w6258 and not w6263;
w6266 <= a(11) and a(41);
w6267 <= not w4998 and not w6266;
w6268 <= w6265 and not w6267;
w6269 <= not w6264 and not w6268;
w6270 <= not w6256 and not w6269;
w6271 <= not w6256 and not w6270;
w6272 <= not w6269 and not w6270;
w6273 <= not w6271 and not w6272;
w6274 <= a(7) and a(45);
w6275 <= a(8) and a(44);
w6276 <= not w6274 and not w6275;
w6277 <= w186 and w5519;
w6278 <= a(37) and not w6277;
w6279 <= a(15) and w6278;
w6280 <= not w6276 and w6279;
w6281 <= a(37) and not w6280;
w6282 <= a(15) and w6281;
w6283 <= not w6277 and not w6280;
w6284 <= not w6276 and w6283;
w6285 <= not w6282 and not w6284;
w6286 <= not w6273 and not w6285;
w6287 <= not w6273 and not w6286;
w6288 <= not w6285 and not w6286;
w6289 <= not w6287 and not w6288;
w6290 <= w1300 and w3618;
w6291 <= a(31) and a(34);
w6292 <= w3454 and w6291;
w6293 <= w1137 and w3896;
w6294 <= not w6292 and not w6293;
w6295 <= not w6290 and not w6294;
w6296 <= not w6290 and not w6295;
w6297 <= a(20) and a(32);
w6298 <= a(21) and a(31);
w6299 <= not w6297 and not w6298;
w6300 <= w6296 and not w6299;
w6301 <= a(34) and not w6295;
w6302 <= a(18) and w6301;
w6303 <= not w6300 and not w6302;
w6304 <= w1472 and w2140;
w6305 <= w1921 and w2916;
w6306 <= w1725 and w2423;
w6307 <= not w6305 and not w6306;
w6308 <= not w6304 and not w6307;
w6309 <= a(30) and not w6308;
w6310 <= a(22) and w6309;
w6311 <= a(23) and a(29);
w6312 <= a(24) and a(28);
w6313 <= not w6311 and not w6312;
w6314 <= not w6304 and not w6308;
w6315 <= not w6313 and w6314;
w6316 <= not w6310 and not w6315;
w6317 <= not w6303 and not w6316;
w6318 <= not w6303 and not w6317;
w6319 <= not w6316 and not w6317;
w6320 <= not w6318 and not w6319;
w6321 <= w5234 and w5971;
w6322 <= a(9) and a(43);
w6323 <= w4007 and w6322;
w6324 <= w551 and w4889;
w6325 <= not w6323 and not w6324;
w6326 <= not w6321 and not w6325;
w6327 <= w4007 and not w6326;
w6328 <= not w6321 and not w6326;
w6329 <= a(13) and a(39);
w6330 <= not w6322 and not w6329;
w6331 <= w6328 and not w6330;
w6332 <= not w6327 and not w6331;
w6333 <= not w6320 and not w6332;
w6334 <= not w6320 and not w6333;
w6335 <= not w6332 and not w6333;
w6336 <= not w6334 and not w6335;
w6337 <= w6289 and w6336;
w6338 <= not w6289 and not w6336;
w6339 <= not w6337 and not w6338;
w6340 <= not w6242 and w6339;
w6341 <= w6242 and not w6339;
w6342 <= not w6340 and not w6341;
w6343 <= not w6241 and w6342;
w6344 <= w6241 and not w6342;
w6345 <= not w6343 and not w6344;
w6346 <= w6240 and not w6345;
w6347 <= not w6240 and w6345;
w6348 <= not w6346 and not w6347;
w6349 <= not w6050 and not w6111;
w6350 <= w6348 and not w6349;
w6351 <= not w6348 and w6349;
w6352 <= not w6350 and not w6351;
w6353 <= not w6239 and w6352;
w6354 <= w6239 and not w6352;
w6355 <= not w6353 and not w6354;
w6356 <= w6125 and not w6355;
w6357 <= not w6125 and w6355;
w6358 <= not w6356 and not w6357;
w6359 <= w6124 and not w6358;
w6360 <= not w6124 and not w6356;
w6361 <= not w6357 and w6360;
w6362 <= not w6359 and not w6361;
w6363 <= not w6357 and not w6360;
w6364 <= not w6350 and not w6353;
w6365 <= not w6175 and not w6236;
w6366 <= not w6228 and not w6232;
w6367 <= a(2) and a(51);
w6368 <= a(3) and a(50);
w6369 <= not w6367 and not w6368;
w6370 <= a(50) and a(51);
w6371 <= w24 and w6370;
w6372 <= not w6369 and not w6371;
w6373 <= w6157 and w6372;
w6374 <= not w6371 and not w6373;
w6375 <= not w6369 and w6374;
w6376 <= w6157 and not w6373;
w6377 <= not w6375 and not w6376;
w6378 <= a(17) and a(36);
w6379 <= a(18) and a(35);
w6380 <= not w6378 and not w6379;
w6381 <= w858 and w3634;
w6382 <= a(4) and not w6381;
w6383 <= a(49) and w6382;
w6384 <= not w6380 and w6383;
w6385 <= a(49) and not w6384;
w6386 <= a(4) and w6385;
w6387 <= not w6381 and not w6384;
w6388 <= not w6380 and w6387;
w6389 <= not w6386 and not w6388;
w6390 <= not w6377 and not w6389;
w6391 <= not w6377 and not w6390;
w6392 <= not w6389 and not w6390;
w6393 <= not w6391 and not w6392;
w6394 <= w1300 and w2949;
w6395 <= w1298 and w3896;
w6396 <= w1296 and w3956;
w6397 <= not w6395 and not w6396;
w6398 <= not w6394 and not w6397;
w6399 <= a(34) and not w6398;
w6400 <= a(19) and w6399;
w6401 <= not w6394 and not w6398;
w6402 <= a(20) and a(33);
w6403 <= a(21) and a(32);
w6404 <= not w6402 and not w6403;
w6405 <= w6401 and not w6404;
w6406 <= not w6400 and not w6405;
w6407 <= not w6393 and not w6406;
w6408 <= not w6393 and not w6407;
w6409 <= not w6406 and not w6407;
w6410 <= not w6408 and not w6409;
w6411 <= not w6141 and not w6147;
w6412 <= w6410 and w6411;
w6413 <= not w6410 and not w6411;
w6414 <= not w6412 and not w6413;
w6415 <= w141 and w5472;
w6416 <= a(6) and a(47);
w6417 <= w4010 and w6416;
w6418 <= not w6415 and not w6417;
w6419 <= a(7) and a(46);
w6420 <= w4010 and w6419;
w6421 <= not w6418 and not w6420;
w6422 <= not w6420 and not w6421;
w6423 <= not w4010 and not w6419;
w6424 <= w6422 and not w6423;
w6425 <= w6416 and not w6421;
w6426 <= not w6424 and not w6425;
w6427 <= a(14) and a(44);
w6428 <= w5234 and w6427;
w6429 <= w238 and w5519;
w6430 <= a(8) and a(45);
w6431 <= a(14) and a(39);
w6432 <= w6430 and w6431;
w6433 <= not w6429 and not w6432;
w6434 <= not w6428 and not w6433;
w6435 <= not w6428 and not w6434;
w6436 <= a(9) and a(44);
w6437 <= not w6431 and not w6436;
w6438 <= w6435 and not w6437;
w6439 <= w6430 and not w6434;
w6440 <= not w6438 and not w6439;
w6441 <= not w6426 and not w6440;
w6442 <= not w6426 and not w6441;
w6443 <= not w6440 and not w6441;
w6444 <= not w6442 and not w6443;
w6445 <= a(5) and a(48);
w6446 <= a(16) and a(37);
w6447 <= not w6445 and not w6446;
w6448 <= a(16) and a(48);
w6449 <= w4048 and w6448;
w6450 <= a(0) and not w6449;
w6451 <= a(53) and w6450;
w6452 <= not w6447 and w6451;
w6453 <= a(53) and not w6452;
w6454 <= a(0) and w6453;
w6455 <= not w6449 and not w6452;
w6456 <= not w6447 and w6455;
w6457 <= not w6454 and not w6456;
w6458 <= not w6444 and not w6457;
w6459 <= not w6444 and not w6458;
w6460 <= not w6457 and not w6458;
w6461 <= not w6459 and not w6460;
w6462 <= not w6414 and w6461;
w6463 <= w6414 and not w6461;
w6464 <= not w6462 and not w6463;
w6465 <= a(10) and a(43);
w6466 <= a(12) and a(41);
w6467 <= not w6465 and not w6466;
w6468 <= w286 and w4613;
w6469 <= w5778 and w5971;
w6470 <= w554 and w5219;
w6471 <= not w6469 and not w6470;
w6472 <= not w6468 and not w6471;
w6473 <= not w6468 and not w6472;
w6474 <= not w6467 and w6473;
w6475 <= a(40) and not w6472;
w6476 <= a(13) and w6475;
w6477 <= not w6474 and not w6476;
w6478 <= w1472 and w2423;
w6479 <= w1921 and w3258;
w6480 <= w1725 and w2671;
w6481 <= not w6479 and not w6480;
w6482 <= not w6478 and not w6481;
w6483 <= w2156 and not w6482;
w6484 <= a(23) and a(30);
w6485 <= a(24) and a(29);
w6486 <= not w6484 and not w6485;
w6487 <= not w6478 and not w6482;
w6488 <= not w6486 and w6487;
w6489 <= not w6483 and not w6488;
w6490 <= not w6477 and not w6489;
w6491 <= not w6477 and not w6490;
w6492 <= not w6489 and not w6490;
w6493 <= not w6491 and not w6492;
w6494 <= a(25) and a(28);
w6495 <= not w2033 and not w6494;
w6496 <= w2137 and w2269;
w6497 <= a(42) and not w6496;
w6498 <= a(11) and w6497;
w6499 <= not w6495 and w6498;
w6500 <= a(42) and not w6499;
w6501 <= a(11) and w6500;
w6502 <= not w6496 and not w6499;
w6503 <= not w6495 and w6502;
w6504 <= not w6501 and not w6503;
w6505 <= not w6493 and not w6504;
w6506 <= not w6493 and not w6505;
w6507 <= not w6504 and not w6505;
w6508 <= not w6506 and not w6507;
w6509 <= not w6165 and not w6168;
w6510 <= w6508 and w6509;
w6511 <= not w6508 and not w6509;
w6512 <= not w6510 and not w6511;
w6513 <= not w6223 and not w6225;
w6514 <= w6512 and not w6513;
w6515 <= not w6512 and w6513;
w6516 <= not w6514 and not w6515;
w6517 <= w6464 and w6516;
w6518 <= not w6464 and not w6516;
w6519 <= not w6517 and not w6518;
w6520 <= not w6366 and w6519;
w6521 <= w6366 and not w6519;
w6522 <= not w6520 and not w6521;
w6523 <= not w6365 and w6522;
w6524 <= w6365 and not w6522;
w6525 <= not w6523 and not w6524;
w6526 <= w6251 and w6296;
w6527 <= not w6251 and not w6296;
w6528 <= not w6526 and not w6527;
w6529 <= w6283 and not w6528;
w6530 <= not w6283 and w6528;
w6531 <= not w6529 and not w6530;
w6532 <= not w6270 and not w6286;
w6533 <= a(52) and w1748;
w6534 <= a(1) and a(52);
w6535 <= not a(27) and not w6534;
w6536 <= not w6533 and not w6535;
w6537 <= w6265 and not w6536;
w6538 <= not w6265 and w6536;
w6539 <= not w6537 and not w6538;
w6540 <= not w6328 and w6539;
w6541 <= w6328 and not w6539;
w6542 <= not w6540 and not w6541;
w6543 <= not w6532 and w6542;
w6544 <= not w6532 and not w6543;
w6545 <= w6542 and not w6543;
w6546 <= not w6544 and not w6545;
w6547 <= w6531 and not w6546;
w6548 <= w6531 and not w6547;
w6549 <= not w6546 and not w6547;
w6550 <= not w6548 and not w6549;
w6551 <= w6138 and w6191;
w6552 <= not w6138 and not w6191;
w6553 <= not w6551 and not w6552;
w6554 <= w6314 and not w6553;
w6555 <= not w6314 and w6553;
w6556 <= not w6554 and not w6555;
w6557 <= not w6317 and not w6333;
w6558 <= not w6179 and not w6195;
w6559 <= w6557 and w6558;
w6560 <= not w6557 and not w6558;
w6561 <= not w6559 and not w6560;
w6562 <= w6556 and w6561;
w6563 <= not w6556 and not w6561;
w6564 <= not w6562 and not w6563;
w6565 <= not w6550 and w6564;
w6566 <= w6564 and not w6565;
w6567 <= not w6550 and not w6565;
w6568 <= not w6566 and not w6567;
w6569 <= not w6151 and not w6171;
w6570 <= w6568 and w6569;
w6571 <= not w6568 and not w6569;
w6572 <= not w6570 and not w6571;
w6573 <= not w6338 and not w6340;
w6574 <= not w6210 and not w6213;
w6575 <= not w6159 and not w6162;
w6576 <= w6574 and w6575;
w6577 <= not w6574 and not w6575;
w6578 <= not w6576 and not w6577;
w6579 <= not w6216 and not w6219;
w6580 <= not w6578 and w6579;
w6581 <= w6578 and not w6579;
w6582 <= not w6580 and not w6581;
w6583 <= not w6201 and not w6205;
w6584 <= not w6582 and w6583;
w6585 <= w6582 and not w6583;
w6586 <= not w6584 and not w6585;
w6587 <= not w6573 and w6586;
w6588 <= w6573 and not w6586;
w6589 <= not w6587 and not w6588;
w6590 <= not w6343 and not w6347;
w6591 <= not w6589 and w6590;
w6592 <= w6589 and not w6590;
w6593 <= not w6591 and not w6592;
w6594 <= w6572 and w6593;
w6595 <= not w6572 and not w6593;
w6596 <= not w6594 and not w6595;
w6597 <= w6525 and w6596;
w6598 <= not w6525 and not w6596;
w6599 <= not w6597 and not w6598;
w6600 <= not w6364 and w6599;
w6601 <= w6364 and not w6599;
w6602 <= not w6600 and not w6601;
w6603 <= not w6363 and not w6602;
w6604 <= w6363 and w6602;
w6605 <= not w6603 and not w6604;
w6606 <= not w6523 and not w6597;
w6607 <= not w6565 and not w6571;
w6608 <= not w6585 and not w6587;
w6609 <= w6607 and w6608;
w6610 <= not w6607 and not w6608;
w6611 <= not w6609 and not w6610;
w6612 <= not w6543 and not w6547;
w6613 <= not w6560 and not w6562;
w6614 <= a(0) and a(54);
w6615 <= w6533 and w6614;
w6616 <= w6533 and not w6615;
w6617 <= not w6533 and w6614;
w6618 <= not w6616 and not w6617;
w6619 <= a(1) and a(53);
w6620 <= w2606 and w6619;
w6621 <= w6619 and not w6620;
w6622 <= w2606 and not w6620;
w6623 <= not w6621 and not w6622;
w6624 <= not w6618 and not w6623;
w6625 <= not w6618 and not w6624;
w6626 <= not w6623 and not w6624;
w6627 <= not w6625 and not w6626;
w6628 <= w1380 and w2949;
w6629 <= a(32) and a(35);
w6630 <= w3842 and w6629;
w6631 <= w1298 and w2778;
w6632 <= not w6630 and not w6631;
w6633 <= not w6628 and not w6632;
w6634 <= not w6628 and not w6633;
w6635 <= a(21) and a(33);
w6636 <= a(22) and a(32);
w6637 <= not w6635 and not w6636;
w6638 <= w6634 and not w6637;
w6639 <= a(35) and not w6633;
w6640 <= a(19) and w6639;
w6641 <= not w6638 and not w6640;
w6642 <= w1710 and w2423;
w6643 <= w1353 and w3258;
w6644 <= w1472 and w2671;
w6645 <= not w6643 and not w6644;
w6646 <= not w6642 and not w6645;
w6647 <= a(31) and not w6646;
w6648 <= a(23) and w6647;
w6649 <= not w6642 and not w6646;
w6650 <= a(25) and a(29);
w6651 <= not w2425 and not w6650;
w6652 <= w6649 and not w6651;
w6653 <= not w6648 and not w6652;
w6654 <= not w6641 and not w6653;
w6655 <= not w6641 and not w6654;
w6656 <= not w6653 and not w6654;
w6657 <= not w6655 and not w6656;
w6658 <= not w6627 and w6657;
w6659 <= w6627 and not w6657;
w6660 <= not w6658 and not w6659;
w6661 <= not w6613 and not w6660;
w6662 <= not w6613 and not w6661;
w6663 <= not w6660 and not w6661;
w6664 <= not w6662 and not w6663;
w6665 <= not w6612 and not w6664;
w6666 <= not w6612 and not w6665;
w6667 <= not w6664 and not w6665;
w6668 <= not w6666 and not w6667;
w6669 <= w6611 and not w6668;
w6670 <= w6611 and not w6669;
w6671 <= not w6668 and not w6669;
w6672 <= not w6670 and not w6671;
w6673 <= not w6592 and not w6594;
w6674 <= not w6672 and not w6673;
w6675 <= not w6672 and not w6674;
w6676 <= not w6673 and not w6674;
w6677 <= not w6675 and not w6676;
w6678 <= not w6517 and not w6520;
w6679 <= not w6527 and not w6530;
w6680 <= not w6552 and not w6555;
w6681 <= w6679 and w6680;
w6682 <= not w6679 and not w6680;
w6683 <= not w6681 and not w6682;
w6684 <= not w6538 and not w6540;
w6685 <= not w6683 and w6684;
w6686 <= w6683 and not w6684;
w6687 <= not w6685 and not w6686;
w6688 <= not w6413 and not w6463;
w6689 <= w6687 and not w6688;
w6690 <= not w6687 and w6688;
w6691 <= not w6689 and not w6690;
w6692 <= w6422 and w6455;
w6693 <= not w6422 and not w6455;
w6694 <= not w6692 and not w6693;
w6695 <= w6502 and not w6694;
w6696 <= not w6502 and w6694;
w6697 <= not w6695 and not w6696;
w6698 <= w6387 and w6401;
w6699 <= not w6387 and not w6401;
w6700 <= not w6698 and not w6699;
w6701 <= w6487 and not w6700;
w6702 <= not w6487 and w6700;
w6703 <= not w6701 and not w6702;
w6704 <= not w6441 and not w6458;
w6705 <= not w6703 and w6704;
w6706 <= w6703 and not w6704;
w6707 <= not w6705 and not w6706;
w6708 <= w6697 and w6707;
w6709 <= not w6697 and not w6707;
w6710 <= not w6708 and not w6709;
w6711 <= w6691 and w6710;
w6712 <= not w6691 and not w6710;
w6713 <= not w6711 and not w6712;
w6714 <= w6678 and not w6713;
w6715 <= not w6678 and w6713;
w6716 <= not w6714 and not w6715;
w6717 <= a(5) and a(49);
w6718 <= a(18) and a(36);
w6719 <= not w6717 and not w6718;
w6720 <= a(20) and a(49);
w6721 <= w3470 and w6720;
w6722 <= w1137 and w4401;
w6723 <= not w6721 and not w6722;
w6724 <= w6717 and w6718;
w6725 <= not w6723 and not w6724;
w6726 <= not w6724 and not w6725;
w6727 <= not w6719 and w6726;
w6728 <= a(34) and not w6725;
w6729 <= a(20) and w6728;
w6730 <= not w6727 and not w6729;
w6731 <= w408 and w4824;
w6732 <= w624 and w4613;
w6733 <= w554 and w5150;
w6734 <= not w6732 and not w6733;
w6735 <= not w6731 and not w6734;
w6736 <= a(41) and not w6735;
w6737 <= a(13) and w6736;
w6738 <= not w6731 and not w6735;
w6739 <= a(11) and a(43);
w6740 <= a(12) and a(42);
w6741 <= not w6739 and not w6740;
w6742 <= w6738 and not w6741;
w6743 <= not w6737 and not w6742;
w6744 <= not w6730 and not w6743;
w6745 <= not w6730 and not w6744;
w6746 <= not w6743 and not w6744;
w6747 <= not w6745 and not w6746;
w6748 <= a(38) and a(48);
w6749 <= w527 and w6748;
w6750 <= a(17) and a(48);
w6751 <= w4294 and w6750;
w6752 <= w854 and w4371;
w6753 <= not w6751 and not w6752;
w6754 <= not w6749 and not w6753;
w6755 <= a(37) and not w6754;
w6756 <= a(17) and w6755;
w6757 <= a(6) and a(48);
w6758 <= a(16) and a(38);
w6759 <= not w6757 and not w6758;
w6760 <= not w6749 and not w6754;
w6761 <= not w6759 and w6760;
w6762 <= not w6756 and not w6761;
w6763 <= not w6747 and not w6762;
w6764 <= not w6747 and not w6763;
w6765 <= not w6762 and not w6763;
w6766 <= not w6764 and not w6765;
w6767 <= not w6577 and not w6581;
w6768 <= w6766 and w6767;
w6769 <= not w6766 and not w6767;
w6770 <= not w6768 and not w6769;
w6771 <= w15 and w6370;
w6772 <= a(50) and a(52);
w6773 <= w58 and w6772;
w6774 <= a(51) and a(52);
w6775 <= w24 and w6774;
w6776 <= not w6773 and not w6775;
w6777 <= not w6771 and not w6776;
w6778 <= not w6771 and not w6777;
w6779 <= a(3) and a(51);
w6780 <= a(4) and a(50);
w6781 <= not w6779 and not w6780;
w6782 <= w6778 and not w6781;
w6783 <= a(52) and not w6777;
w6784 <= a(2) and w6783;
w6785 <= not w6782 and not w6784;
w6786 <= a(7) and a(47);
w6787 <= a(15) and a(39);
w6788 <= w6786 and w6787;
w6789 <= w186 and w5472;
w6790 <= not w6788 and not w6789;
w6791 <= a(8) and a(46);
w6792 <= w6787 and w6791;
w6793 <= not w6790 and not w6792;
w6794 <= w6786 and not w6793;
w6795 <= not w6792 and not w6793;
w6796 <= not w6787 and not w6791;
w6797 <= w6795 and not w6796;
w6798 <= not w6794 and not w6797;
w6799 <= not w6785 and not w6798;
w6800 <= not w6785 and not w6799;
w6801 <= not w6798 and not w6799;
w6802 <= not w6800 and not w6801;
w6803 <= a(9) and a(45);
w6804 <= w5778 and w6427;
w6805 <= w290 and w5519;
w6806 <= w4661 and w6803;
w6807 <= not w6805 and not w6806;
w6808 <= not w6804 and not w6807;
w6809 <= w6803 and not w6808;
w6810 <= not w6804 and not w6808;
w6811 <= a(10) and a(44);
w6812 <= not w4661 and not w6811;
w6813 <= w6810 and not w6812;
w6814 <= not w6809 and not w6813;
w6815 <= not w6802 and not w6814;
w6816 <= not w6802 and not w6815;
w6817 <= not w6814 and not w6815;
w6818 <= not w6816 and not w6817;
w6819 <= not w6770 and w6818;
w6820 <= w6770 and not w6818;
w6821 <= not w6819 and not w6820;
w6822 <= not w6511 and not w6514;
w6823 <= w6374 and w6435;
w6824 <= not w6374 and not w6435;
w6825 <= not w6823 and not w6824;
w6826 <= w6473 and not w6825;
w6827 <= not w6473 and w6825;
w6828 <= not w6826 and not w6827;
w6829 <= not w6490 and not w6505;
w6830 <= not w6390 and not w6407;
w6831 <= w6829 and w6830;
w6832 <= not w6829 and not w6830;
w6833 <= not w6831 and not w6832;
w6834 <= w6828 and w6833;
w6835 <= not w6828 and not w6833;
w6836 <= not w6834 and not w6835;
w6837 <= not w6822 and w6836;
w6838 <= not w6822 and not w6837;
w6839 <= w6836 and not w6837;
w6840 <= not w6838 and not w6839;
w6841 <= w6821 and not w6840;
w6842 <= w6821 and not w6841;
w6843 <= not w6840 and not w6841;
w6844 <= not w6842 and not w6843;
w6845 <= w6716 and not w6844;
w6846 <= w6716 and not w6845;
w6847 <= not w6844 and not w6845;
w6848 <= not w6846 and not w6847;
w6849 <= not w6677 and w6848;
w6850 <= w6677 and not w6848;
w6851 <= not w6849 and not w6850;
w6852 <= not w6606 and not w6851;
w6853 <= w6606 and w6851;
w6854 <= not w6852 and not w6853;
w6855 <= not w6363 and not w6601;
w6856 <= not w6600 and not w6855;
w6857 <= not w6854 and w6856;
w6858 <= w6854 and not w6856;
w6859 <= not w6857 and not w6858;
w6860 <= not w6677 and not w6848;
w6861 <= not w6674 and not w6860;
w6862 <= not w6715 and not w6845;
w6863 <= not w6837 and not w6841;
w6864 <= not w6689 and not w6711;
w6865 <= not w6706 and not w6708;
w6866 <= a(6) and a(49);
w6867 <= a(17) and a(38);
w6868 <= not w6866 and not w6867;
w6869 <= a(17) and a(49);
w6870 <= w4366 and w6869;
w6871 <= a(3) and not w6870;
w6872 <= a(52) and w6871;
w6873 <= not w6868 and w6872;
w6874 <= not w6870 and not w6873;
w6875 <= not w6868 and w6874;
w6876 <= a(52) and not w6873;
w6877 <= a(3) and w6876;
w6878 <= not w6875 and not w6877;
w6879 <= a(40) and a(46);
w6880 <= w1323 and w6879;
w6881 <= w701 and w5219;
w6882 <= not w6880 and not w6881;
w6883 <= a(9) and a(46);
w6884 <= a(14) and a(41);
w6885 <= w6883 and w6884;
w6886 <= not w6882 and not w6885;
w6887 <= a(40) and not w6886;
w6888 <= a(15) and w6887;
w6889 <= not w6883 and not w6884;
w6890 <= not w6885 and not w6886;
w6891 <= not w6889 and w6890;
w6892 <= not w6888 and not w6891;
w6893 <= not w6878 and not w6892;
w6894 <= not w6878 and not w6893;
w6895 <= not w6892 and not w6893;
w6896 <= not w6894 and not w6895;
w6897 <= not w6699 and not w6702;
w6898 <= w6896 and w6897;
w6899 <= not w6896 and not w6897;
w6900 <= not w6898 and not w6899;
w6901 <= not w6832 and not w6834;
w6902 <= w6900 and not w6901;
w6903 <= not w6900 and w6901;
w6904 <= not w6902 and not w6903;
w6905 <= not w6865 and w6904;
w6906 <= w6865 and not w6904;
w6907 <= not w6905 and not w6906;
w6908 <= not w6864 and w6907;
w6909 <= not w6864 and not w6908;
w6910 <= w6907 and not w6908;
w6911 <= not w6909 and not w6910;
w6912 <= not w6863 and not w6911;
w6913 <= not w6863 and not w6912;
w6914 <= not w6911 and not w6912;
w6915 <= not w6913 and not w6914;
w6916 <= not w6862 and not w6915;
w6917 <= not w6862 and not w6916;
w6918 <= not w6915 and not w6916;
w6919 <= not w6917 and not w6918;
w6920 <= not w6693 and not w6696;
w6921 <= not w6824 and not w6827;
w6922 <= w6920 and w6921;
w6923 <= not w6920 and not w6921;
w6924 <= not w6922 and not w6923;
w6925 <= a(28) and a(54);
w6926 <= a(1) and w6925;
w6927 <= a(1) and a(54);
w6928 <= not a(28) and not w6927;
w6929 <= not w6926 and not w6928;
w6930 <= w6620 and w6929;
w6931 <= w6620 and not w6930;
w6932 <= w6929 and not w6930;
w6933 <= not w6931 and not w6932;
w6934 <= not w6738 and not w6933;
w6935 <= not w6738 and not w6934;
w6936 <= not w6933 and not w6934;
w6937 <= not w6935 and not w6936;
w6938 <= w6924 and not w6937;
w6939 <= w6924 and not w6938;
w6940 <= not w6937 and not w6938;
w6941 <= not w6939 and not w6940;
w6942 <= not w6769 and not w6820;
w6943 <= not w6941 and not w6942;
w6944 <= not w6941 and not w6943;
w6945 <= not w6942 and not w6943;
w6946 <= not w6944 and not w6945;
w6947 <= not w6615 and not w6624;
w6948 <= w6795 and w6947;
w6949 <= not w6795 and not w6947;
w6950 <= not w6948 and not w6949;
w6951 <= a(18) and a(37);
w6952 <= a(19) and a(36);
w6953 <= not w6951 and not w6952;
w6954 <= w955 and w3493;
w6955 <= a(5) and not w6954;
w6956 <= a(50) and w6955;
w6957 <= not w6953 and w6956;
w6958 <= a(50) and not w6957;
w6959 <= a(5) and w6958;
w6960 <= not w6954 and not w6957;
w6961 <= not w6953 and w6960;
w6962 <= not w6959 and not w6961;
w6963 <= w6950 and not w6962;
w6964 <= w6950 and not w6963;
w6965 <= not w6962 and not w6963;
w6966 <= not w6964 and not w6965;
w6967 <= w6778 and w6810;
w6968 <= not w6778 and not w6810;
w6969 <= not w6967 and not w6968;
w6970 <= w6726 and not w6969;
w6971 <= not w6726 and w6969;
w6972 <= not w6970 and not w6971;
w6973 <= not w6627 and not w6657;
w6974 <= not w6654 and not w6973;
w6975 <= w6972 and not w6974;
w6976 <= not w6972 and w6974;
w6977 <= not w6975 and not w6976;
w6978 <= not w6966 and w6977;
w6979 <= not w6966 and not w6978;
w6980 <= w6977 and not w6978;
w6981 <= not w6979 and not w6980;
w6982 <= not w6946 and not w6981;
w6983 <= not w6946 and not w6982;
w6984 <= not w6981 and not w6982;
w6985 <= not w6983 and not w6984;
w6986 <= not w6610 and not w6669;
w6987 <= w6985 and w6986;
w6988 <= not w6985 and not w6986;
w6989 <= not w6987 and not w6988;
w6990 <= w624 and w4445;
w6991 <= w529 and w5519;
w6992 <= a(13) and a(45);
w6993 <= w6257 and w6992;
w6994 <= not w6991 and not w6993;
w6995 <= not w6990 and not w6994;
w6996 <= not w6990 and not w6995;
w6997 <= a(11) and a(44);
w6998 <= not w5755 and not w6997;
w6999 <= w6996 and not w6998;
w7000 <= a(45) and not w6995;
w7001 <= a(10) and w7000;
w7002 <= not w6999 and not w7001;
w7003 <= a(26) and a(29);
w7004 <= not w2137 and not w7003;
w7005 <= w2137 and w7003;
w7006 <= a(43) and not w7005;
w7007 <= a(12) and w7006;
w7008 <= not w7004 and w7007;
w7009 <= a(43) and not w7008;
w7010 <= a(12) and w7009;
w7011 <= not w7005 and not w7008;
w7012 <= not w7004 and w7011;
w7013 <= not w7010 and not w7012;
w7014 <= not w7002 and not w7013;
w7015 <= not w7002 and not w7014;
w7016 <= not w7013 and not w7014;
w7017 <= not w7015 and not w7016;
w7018 <= a(7) and a(48);
w7019 <= a(8) and a(47);
w7020 <= not w7018 and not w7019;
w7021 <= w186 and w6058;
w7022 <= a(39) and not w7021;
w7023 <= a(16) and w7022;
w7024 <= not w7020 and w7023;
w7025 <= a(39) and not w7024;
w7026 <= a(16) and w7025;
w7027 <= not w7021 and not w7024;
w7028 <= not w7020 and w7027;
w7029 <= not w7026 and not w7028;
w7030 <= not w7017 and not w7029;
w7031 <= not w7017 and not w7030;
w7032 <= not w7029 and not w7030;
w7033 <= not w7031 and not w7032;
w7034 <= not w6682 and not w6686;
w7035 <= w7033 and w7034;
w7036 <= not w7033 and not w7034;
w7037 <= not w7035 and not w7036;
w7038 <= a(51) and a(53);
w7039 <= w58 and w7038;
w7040 <= a(51) and w18;
w7041 <= a(53) and w2;
w7042 <= not w7040 and not w7041;
w7043 <= a(55) and not w7039;
w7044 <= not w7042 and w7043;
w7045 <= not w7039 and not w7044;
w7046 <= a(2) and a(53);
w7047 <= a(4) and a(51);
w7048 <= not w7046 and not w7047;
w7049 <= w7045 and not w7048;
w7050 <= a(55) and not w7044;
w7051 <= a(0) and w7050;
w7052 <= not w7049 and not w7051;
w7053 <= w1380 and w3956;
w7054 <= w1499 and w2778;
w7055 <= w1300 and w3125;
w7056 <= not w7054 and not w7055;
w7057 <= not w7053 and not w7056;
w7058 <= a(35) and not w7057;
w7059 <= a(20) and w7058;
w7060 <= not w7053 and not w7057;
w7061 <= a(21) and a(34);
w7062 <= not w2401 and not w7061;
w7063 <= w7060 and not w7062;
w7064 <= not w7059 and not w7063;
w7065 <= not w7052 and not w7064;
w7066 <= not w7052 and not w7065;
w7067 <= not w7064 and not w7065;
w7068 <= not w7066 and not w7067;
w7069 <= a(23) and a(32);
w7070 <= w1710 and w2671;
w7071 <= w1353 and w2294;
w7072 <= w1472 and w3618;
w7073 <= not w7071 and not w7072;
w7074 <= not w7070 and not w7073;
w7075 <= w7069 and not w7074;
w7076 <= not w7070 and not w7074;
w7077 <= a(24) and a(31);
w7078 <= a(25) and a(30);
w7079 <= not w7077 and not w7078;
w7080 <= w7076 and not w7079;
w7081 <= not w7075 and not w7080;
w7082 <= not w7068 and not w7081;
w7083 <= not w7068 and not w7082;
w7084 <= not w7081 and not w7082;
w7085 <= not w7083 and not w7084;
w7086 <= w7037 and not w7085;
w7087 <= not w7037 and w7085;
w7088 <= not w6661 and not w6665;
w7089 <= w6634 and w6649;
w7090 <= not w6634 and not w6649;
w7091 <= not w7089 and not w7090;
w7092 <= w6760 and not w7091;
w7093 <= not w6760 and w7091;
w7094 <= not w7092 and not w7093;
w7095 <= not w6744 and not w6763;
w7096 <= not w6799 and not w6815;
w7097 <= w7095 and w7096;
w7098 <= not w7095 and not w7096;
w7099 <= not w7097 and not w7098;
w7100 <= w7094 and w7099;
w7101 <= not w7094 and not w7099;
w7102 <= not w7100 and not w7101;
w7103 <= not w7088 and w7102;
w7104 <= w7088 and not w7102;
w7105 <= not w7103 and not w7104;
w7106 <= not w7087 and w7105;
w7107 <= not w7086 and w7106;
w7108 <= w7105 and not w7107;
w7109 <= not w7087 and not w7107;
w7110 <= not w7086 and w7109;
w7111 <= not w7108 and not w7110;
w7112 <= not w6989 and w7111;
w7113 <= w6989 and not w7111;
w7114 <= not w7112 and not w7113;
w7115 <= not w6919 and w7114;
w7116 <= w6919 and not w7114;
w7117 <= not w7115 and not w7116;
w7118 <= not w6861 and w7117;
w7119 <= w6861 and not w7117;
w7120 <= not w7118 and not w7119;
w7121 <= not w6853 and not w6856;
w7122 <= not w6852 and not w7121;
w7123 <= not w7120 and w7122;
w7124 <= w7120 and not w7122;
w7125 <= not w7123 and not w7124;
w7126 <= not w6916 and not w7115;
w7127 <= a(7) and a(49);
w7128 <= a(17) and a(39);
w7129 <= not w7127 and not w7128;
w7130 <= w141 and w6131;
w7131 <= a(17) and a(50);
w7132 <= w4552 and w7131;
w7133 <= not w7130 and not w7132;
w7134 <= w7127 and w7128;
w7135 <= not w7133 and not w7134;
w7136 <= not w7134 and not w7135;
w7137 <= not w7129 and w7136;
w7138 <= a(50) and not w7135;
w7139 <= a(6) and w7138;
w7140 <= not w7137 and not w7139;
w7141 <= w554 and w5102;
w7142 <= w624 and w4617;
w7143 <= w408 and w5519;
w7144 <= not w7142 and not w7143;
w7145 <= not w7141 and not w7144;
w7146 <= a(45) and not w7145;
w7147 <= a(11) and w7146;
w7148 <= a(12) and a(44);
w7149 <= not w5971 and not w7148;
w7150 <= not w7141 and not w7145;
w7151 <= not w7149 and w7150;
w7152 <= not w7147 and not w7151;
w7153 <= not w7140 and not w7152;
w7154 <= not w7140 and not w7153;
w7155 <= not w7152 and not w7153;
w7156 <= not w7154 and not w7155;
w7157 <= a(15) and a(48);
w7158 <= w5426 and w7157;
w7159 <= a(40) and a(48);
w7160 <= w1315 and w7159;
w7161 <= w697 and w5219;
w7162 <= not w7160 and not w7161;
w7163 <= not w7158 and not w7162;
w7164 <= w3975 and not w7163;
w7165 <= not w7158 and not w7163;
w7166 <= a(8) and a(48);
w7167 <= a(15) and a(41);
w7168 <= not w7166 and not w7167;
w7169 <= w7165 and not w7168;
w7170 <= not w7164 and not w7169;
w7171 <= not w7156 and not w7170;
w7172 <= not w7156 and not w7171;
w7173 <= not w7170 and not w7171;
w7174 <= not w7172 and not w7173;
w7175 <= w1725 and w3956;
w7176 <= w1499 and w4401;
w7177 <= a(33) and a(36);
w7178 <= w4229 and w7177;
w7179 <= not w7176 and not w7178;
w7180 <= not w7175 and not w7179;
w7181 <= not w7175 and not w7180;
w7182 <= a(22) and a(34);
w7183 <= a(23) and a(33);
w7184 <= not w7182 and not w7183;
w7185 <= w7181 and not w7184;
w7186 <= a(36) and not w7180;
w7187 <= a(20) and w7186;
w7188 <= not w7185 and not w7187;
w7189 <= w2269 and w2671;
w7190 <= w2107 and w2294;
w7191 <= w1710 and w3618;
w7192 <= not w7190 and not w7191;
w7193 <= not w7189 and not w7192;
w7194 <= a(32) and not w7193;
w7195 <= a(24) and w7194;
w7196 <= not w7189 and not w7193;
w7197 <= a(25) and a(31);
w7198 <= a(26) and a(30);
w7199 <= not w7197 and not w7198;
w7200 <= w7196 and not w7199;
w7201 <= not w7195 and not w7200;
w7202 <= not w7188 and not w7201;
w7203 <= not w7188 and not w7202;
w7204 <= not w7201 and not w7202;
w7205 <= not w7203 and not w7204;
w7206 <= a(14) and a(46);
w7207 <= w6257 and w7206;
w7208 <= w290 and w5472;
w7209 <= a(14) and a(47);
w7210 <= w5986 and w7209;
w7211 <= not w7208 and not w7210;
w7212 <= not w7207 and not w7211;
w7213 <= a(47) and not w7212;
w7214 <= a(9) and w7213;
w7215 <= not w7207 and not w7212;
w7216 <= a(10) and a(46);
w7217 <= not w5152 and not w7216;
w7218 <= w7215 and not w7217;
w7219 <= not w7214 and not w7218;
w7220 <= not w7205 and not w7219;
w7221 <= not w7205 and not w7220;
w7222 <= not w7219 and not w7220;
w7223 <= not w7221 and not w7222;
w7224 <= not w7174 and w7223;
w7225 <= w7174 and not w7223;
w7226 <= not w7224 and not w7225;
w7227 <= a(54) and a(56);
w7228 <= w2 and w7227;
w7229 <= a(0) and a(56);
w7230 <= a(2) and a(54);
w7231 <= not w7229 and not w7230;
w7232 <= not w7228 and not w7231;
w7233 <= w6926 and w7232;
w7234 <= not w6926 and not w7232;
w7235 <= not w7233 and not w7234;
w7236 <= not w7027 and w7235;
w7237 <= w7027 and not w7235;
w7238 <= not w7236 and not w7237;
w7239 <= a(52) and a(53);
w7240 <= w15 and w7239;
w7241 <= a(37) and a(53);
w7242 <= w1079 and w7241;
w7243 <= not w7240 and not w7242;
w7244 <= a(4) and a(52);
w7245 <= a(19) and a(37);
w7246 <= w7244 and w7245;
w7247 <= not w7243 and not w7246;
w7248 <= a(53) and not w7247;
w7249 <= a(3) and w7248;
w7250 <= not w7246 and not w7247;
w7251 <= not w7244 and not w7245;
w7252 <= w7250 and not w7251;
w7253 <= not w7249 and not w7252;
w7254 <= w7238 and not w7253;
w7255 <= w7238 and not w7254;
w7256 <= not w7253 and not w7254;
w7257 <= not w7255 and not w7256;
w7258 <= w7226 and w7257;
w7259 <= not w7226 and not w7257;
w7260 <= not w7258 and not w7259;
w7261 <= not w6902 and not w6905;
w7262 <= w7060 and w7076;
w7263 <= not w7060 and not w7076;
w7264 <= not w7262 and not w7263;
w7265 <= w6874 and not w7264;
w7266 <= not w6874 and w7264;
w7267 <= not w7265 and not w7266;
w7268 <= not w7014 and not w7030;
w7269 <= a(1) and a(55);
w7270 <= not w1847 and not w7269;
w7271 <= w1847 and w7269;
w7272 <= not w7011 and not w7271;
w7273 <= not w7270 and w7272;
w7274 <= not w7011 and not w7273;
w7275 <= not w7271 and not w7273;
w7276 <= not w7270 and w7275;
w7277 <= not w7274 and not w7276;
w7278 <= not w6996 and not w7277;
w7279 <= w6996 and not w7276;
w7280 <= not w7274 and w7279;
w7281 <= not w7278 and not w7280;
w7282 <= not w7268 and w7281;
w7283 <= w7268 and not w7281;
w7284 <= not w7282 and not w7283;
w7285 <= w7267 and w7284;
w7286 <= not w7267 and not w7284;
w7287 <= not w7285 and not w7286;
w7288 <= not w7261 and w7287;
w7289 <= not w7261 and not w7288;
w7290 <= w7287 and not w7288;
w7291 <= not w7289 and not w7290;
w7292 <= w7260 and not w7291;
w7293 <= w7260 and not w7292;
w7294 <= not w7291 and not w7292;
w7295 <= not w7293 and not w7294;
w7296 <= not w6908 and not w6912;
w7297 <= w6960 and w7045;
w7298 <= not w6960 and not w7045;
w7299 <= not w7297 and not w7298;
w7300 <= w6890 and not w7299;
w7301 <= not w6890 and w7299;
w7302 <= not w7300 and not w7301;
w7303 <= not w6893 and not w6899;
w7304 <= not w7302 and w7303;
w7305 <= w7302 and not w7303;
w7306 <= not w7304 and not w7305;
w7307 <= not w6923 and not w6938;
w7308 <= not w7306 and w7307;
w7309 <= w7306 and not w7307;
w7310 <= not w7308 and not w7309;
w7311 <= not w7090 and not w7093;
w7312 <= not w6949 and not w6963;
w7313 <= w7311 and w7312;
w7314 <= not w7311 and not w7312;
w7315 <= not w7313 and not w7314;
w7316 <= not w7065 and not w7082;
w7317 <= not w7315 and w7316;
w7318 <= w7315 and not w7316;
w7319 <= not w7317 and not w7318;
w7320 <= not w7036 and not w7086;
w7321 <= w7319 and not w7320;
w7322 <= w7319 and not w7321;
w7323 <= not w7320 and not w7321;
w7324 <= not w7322 and not w7323;
w7325 <= w7310 and not w7324;
w7326 <= not w7310 and not w7323;
w7327 <= not w7322 and w7326;
w7328 <= not w7325 and not w7327;
w7329 <= not w7296 and w7328;
w7330 <= not w7296 and not w7329;
w7331 <= w7328 and not w7329;
w7332 <= not w7330 and not w7331;
w7333 <= not w7295 and not w7332;
w7334 <= not w7295 and not w7333;
w7335 <= not w7332 and not w7333;
w7336 <= not w7334 and not w7335;
w7337 <= not w6975 and not w6978;
w7338 <= not w6930 and not w6934;
w7339 <= a(5) and a(51);
w7340 <= a(18) and a(38);
w7341 <= not w7339 and not w7340;
w7342 <= a(38) and a(51);
w7343 <= w1146 and w7342;
w7344 <= a(35) and not w7343;
w7345 <= a(21) and w7344;
w7346 <= not w7341 and w7345;
w7347 <= a(35) and not w7346;
w7348 <= a(21) and w7347;
w7349 <= not w7343 and not w7346;
w7350 <= not w7341 and w7349;
w7351 <= not w7348 and not w7350;
w7352 <= not w7338 and not w7351;
w7353 <= not w7338 and not w7352;
w7354 <= not w7351 and not w7352;
w7355 <= not w7353 and not w7354;
w7356 <= not w6968 and not w6971;
w7357 <= w7355 and w7356;
w7358 <= not w7355 and not w7356;
w7359 <= not w7357 and not w7358;
w7360 <= not w7098 and not w7100;
w7361 <= w7359 and not w7360;
w7362 <= not w7359 and w7360;
w7363 <= not w7361 and not w7362;
w7364 <= w7337 and not w7363;
w7365 <= not w7337 and w7363;
w7366 <= not w7364 and not w7365;
w7367 <= not w6943 and not w6982;
w7368 <= not w7366 and w7367;
w7369 <= w7366 and not w7367;
w7370 <= not w7368 and not w7369;
w7371 <= not w7103 and not w7107;
w7372 <= not w7370 and w7371;
w7373 <= w7370 and not w7371;
w7374 <= not w7372 and not w7373;
w7375 <= not w6988 and not w7113;
w7376 <= w7374 and not w7375;
w7377 <= w7374 and not w7376;
w7378 <= not w7375 and not w7376;
w7379 <= not w7377 and not w7378;
w7380 <= not w7336 and not w7379;
w7381 <= w7336 and not w7378;
w7382 <= not w7377 and w7381;
w7383 <= not w7380 and not w7382;
w7384 <= not w7126 and w7383;
w7385 <= w7126 and not w7383;
w7386 <= not w7384 and not w7385;
w7387 <= not w7119 and not w7122;
w7388 <= not w7118 and not w7387;
w7389 <= not w7386 and w7388;
w7390 <= w7386 and not w7388;
w7391 <= not w7389 and not w7390;
w7392 <= not w7376 and not w7380;
w7393 <= not w7369 and not w7373;
w7394 <= not w7273 and not w7278;
w7395 <= not w7236 and not w7254;
w7396 <= w7394 and w7395;
w7397 <= not w7394 and not w7395;
w7398 <= not w7396 and not w7397;
w7399 <= not w7202 and not w7220;
w7400 <= not w7398 and w7399;
w7401 <= w7398 and not w7399;
w7402 <= not w7400 and not w7401;
w7403 <= not w7174 and not w7223;
w7404 <= not w7259 and not w7403;
w7405 <= w7402 and not w7404;
w7406 <= not w7402 and w7404;
w7407 <= not w7405 and not w7406;
w7408 <= not w7153 and not w7171;
w7409 <= w7165 and w7196;
w7410 <= not w7165 and not w7196;
w7411 <= not w7409 and not w7410;
w7412 <= w7136 and not w7411;
w7413 <= not w7136 and w7411;
w7414 <= not w7412 and not w7413;
w7415 <= w7181 and w7250;
w7416 <= not w7181 and not w7250;
w7417 <= not w7415 and not w7416;
w7418 <= not w7228 and not w7233;
w7419 <= not w7417 and w7418;
w7420 <= w7417 and not w7418;
w7421 <= not w7419 and not w7420;
w7422 <= w7414 and w7421;
w7423 <= not w7414 and not w7421;
w7424 <= not w7422 and not w7423;
w7425 <= not w7408 and w7424;
w7426 <= w7408 and not w7424;
w7427 <= not w7425 and not w7426;
w7428 <= w7407 and w7427;
w7429 <= not w7407 and not w7427;
w7430 <= not w7428 and not w7429;
w7431 <= w7393 and not w7430;
w7432 <= not w7393 and w7430;
w7433 <= not w7431 and not w7432;
w7434 <= not w7361 and not w7365;
w7435 <= w7215 and w7349;
w7436 <= not w7215 and not w7349;
w7437 <= not w7435 and not w7436;
w7438 <= w7150 and not w7437;
w7439 <= not w7150 and w7437;
w7440 <= not w7438 and not w7439;
w7441 <= not w7352 and not w7358;
w7442 <= not w7440 and w7441;
w7443 <= w7440 and not w7441;
w7444 <= not w7442 and not w7443;
w7445 <= a(16) and a(49);
w7446 <= w5426 and w7445;
w7447 <= w186 and w6131;
w7448 <= a(16) and a(50);
w7449 <= w5217 and w7448;
w7450 <= not w7447 and not w7449;
w7451 <= not w7446 and not w7450;
w7452 <= not w7446 and not w7451;
w7453 <= a(8) and a(49);
w7454 <= a(16) and a(41);
w7455 <= not w7453 and not w7454;
w7456 <= w7452 and not w7455;
w7457 <= a(50) and not w7451;
w7458 <= a(7) and w7457;
w7459 <= not w7456 and not w7458;
w7460 <= w1725 and w3125;
w7461 <= w1173 and w4401;
w7462 <= w1380 and w3634;
w7463 <= not w7461 and not w7462;
w7464 <= not w7460 and not w7463;
w7465 <= a(36) and not w7464;
w7466 <= a(21) and w7465;
w7467 <= a(22) and a(35);
w7468 <= a(23) and a(34);
w7469 <= not w7467 and not w7468;
w7470 <= not w7460 and not w7464;
w7471 <= not w7469 and w7470;
w7472 <= not w7466 and not w7471;
w7473 <= not w7459 and not w7472;
w7474 <= not w7459 and not w7473;
w7475 <= not w7472 and not w7473;
w7476 <= not w7474 and not w7475;
w7477 <= w2269 and w3618;
w7478 <= w2107 and w2404;
w7479 <= w1710 and w2949;
w7480 <= not w7478 and not w7479;
w7481 <= not w7477 and not w7480;
w7482 <= a(33) and not w7481;
w7483 <= a(24) and w7482;
w7484 <= not w7477 and not w7481;
w7485 <= a(25) and a(32);
w7486 <= a(26) and a(31);
w7487 <= not w7485 and not w7486;
w7488 <= w7484 and not w7487;
w7489 <= not w7483 and not w7488;
w7490 <= not w7476 and not w7489;
w7491 <= not w7476 and not w7490;
w7492 <= not w7489 and not w7490;
w7493 <= not w7491 and not w7492;
w7494 <= w7444 and not w7493;
w7495 <= not w7444 and w7493;
w7496 <= not w7434 and not w7495;
w7497 <= not w7494 and w7496;
w7498 <= not w7434 and not w7497;
w7499 <= not w7495 and not w7497;
w7500 <= not w7494 and w7499;
w7501 <= not w7498 and not w7500;
w7502 <= not w7314 and not w7318;
w7503 <= a(53) and a(55);
w7504 <= w58 and w7503;
w7505 <= a(53) and a(54);
w7506 <= w15 and w7505;
w7507 <= a(54) and a(55);
w7508 <= w24 and w7507;
w7509 <= not w7506 and not w7508;
w7510 <= not w7504 and not w7509;
w7511 <= not w7504 and not w7510;
w7512 <= a(2) and a(55);
w7513 <= a(4) and a(53);
w7514 <= not w7512 and not w7513;
w7515 <= w7511 and not w7514;
w7516 <= a(54) and not w7510;
w7517 <= a(3) and w7516;
w7518 <= not w7515 and not w7517;
w7519 <= a(19) and a(38);
w7520 <= a(20) and a(37);
w7521 <= not w7519 and not w7520;
w7522 <= w1296 and w4371;
w7523 <= a(5) and not w7522;
w7524 <= a(52) and w7523;
w7525 <= not w7521 and w7524;
w7526 <= a(52) and not w7525;
w7527 <= a(5) and w7526;
w7528 <= not w7522 and not w7525;
w7529 <= not w7521 and w7528;
w7530 <= not w7527 and not w7529;
w7531 <= not w7518 and not w7530;
w7532 <= not w7518 and not w7531;
w7533 <= not w7530 and not w7531;
w7534 <= not w7532 and not w7533;
w7535 <= a(9) and a(48);
w7536 <= a(10) and a(47);
w7537 <= not w7535 and not w7536;
w7538 <= w290 and w6058;
w7539 <= a(42) and not w7538;
w7540 <= a(15) and w7539;
w7541 <= not w7537 and w7540;
w7542 <= a(42) and not w7541;
w7543 <= a(15) and w7542;
w7544 <= not w7538 and not w7541;
w7545 <= not w7537 and w7544;
w7546 <= not w7543 and not w7545;
w7547 <= not w7534 and not w7546;
w7548 <= not w7534 and not w7547;
w7549 <= not w7546 and not w7547;
w7550 <= not w7548 and not w7549;
w7551 <= a(11) and a(46);
w7552 <= not w5974 and not w7551;
w7553 <= a(44) and a(46);
w7554 <= w624 and w7553;
w7555 <= w551 and w5102;
w7556 <= w6739 and w7206;
w7557 <= not w7555 and not w7556;
w7558 <= not w7554 and not w7557;
w7559 <= not w7554 and not w7558;
w7560 <= not w7552 and w7559;
w7561 <= a(43) and not w7558;
w7562 <= a(14) and w7561;
w7563 <= not w7560 and not w7562;
w7564 <= not w2140 and not w2728;
w7565 <= w2137 and w2423;
w7566 <= a(45) and not w7565;
w7567 <= a(12) and w7566;
w7568 <= not w7564 and w7567;
w7569 <= a(45) and not w7568;
w7570 <= a(12) and w7569;
w7571 <= not w7565 and not w7568;
w7572 <= not w7564 and w7571;
w7573 <= not w7570 and not w7572;
w7574 <= not w7563 and not w7573;
w7575 <= not w7563 and not w7574;
w7576 <= not w7573 and not w7574;
w7577 <= not w7575 and not w7576;
w7578 <= a(17) and a(51);
w7579 <= w4778 and w7578;
w7580 <= a(39) and a(51);
w7581 <= w1284 and w7580;
w7582 <= w858 and w3977;
w7583 <= not w7581 and not w7582;
w7584 <= not w7579 and not w7583;
w7585 <= a(39) and not w7584;
w7586 <= a(18) and w7585;
w7587 <= not w7579 and not w7584;
w7588 <= a(6) and a(51);
w7589 <= a(17) and a(40);
w7590 <= not w7588 and not w7589;
w7591 <= w7587 and not w7590;
w7592 <= not w7586 and not w7591;
w7593 <= not w7577 and not w7592;
w7594 <= not w7577 and not w7593;
w7595 <= not w7592 and not w7593;
w7596 <= not w7594 and not w7595;
w7597 <= w7550 and w7596;
w7598 <= not w7550 and not w7596;
w7599 <= not w7597 and not w7598;
w7600 <= not w7502 and w7599;
w7601 <= w7502 and not w7599;
w7602 <= not w7600 and not w7601;
w7603 <= w7501 and w7602;
w7604 <= not w7501 and not w7602;
w7605 <= not w7603 and not w7604;
w7606 <= w7433 and not w7605;
w7607 <= w7433 and not w7606;
w7608 <= not w7605 and not w7606;
w7609 <= not w7607 and not w7608;
w7610 <= not w7329 and not w7333;
w7611 <= not w7288 and not w7292;
w7612 <= not w7321 and not w7325;
w7613 <= not w7305 and not w7309;
w7614 <= not w7282 and not w7285;
w7615 <= w7613 and w7614;
w7616 <= not w7613 and not w7614;
w7617 <= not w7615 and not w7616;
w7618 <= a(0) and a(57);
w7619 <= w7271 and w7618;
w7620 <= w7271 and not w7619;
w7621 <= not w7271 and w7618;
w7622 <= not w7620 and not w7621;
w7623 <= a(1) and a(56);
w7624 <= a(29) and w7623;
w7625 <= a(29) and not w7624;
w7626 <= w7623 and not w7624;
w7627 <= not w7625 and not w7626;
w7628 <= not w7622 and not w7627;
w7629 <= not w7622 and not w7628;
w7630 <= not w7627 and not w7628;
w7631 <= not w7629 and not w7630;
w7632 <= not w7263 and not w7266;
w7633 <= w7631 and w7632;
w7634 <= not w7631 and not w7632;
w7635 <= not w7633 and not w7634;
w7636 <= not w7298 and not w7301;
w7637 <= not w7635 and w7636;
w7638 <= w7635 and not w7636;
w7639 <= not w7637 and not w7638;
w7640 <= w7617 and w7639;
w7641 <= not w7617 and not w7639;
w7642 <= not w7640 and not w7641;
w7643 <= not w7612 and w7642;
w7644 <= w7612 and not w7642;
w7645 <= not w7643 and not w7644;
w7646 <= not w7611 and w7645;
w7647 <= w7611 and not w7645;
w7648 <= not w7646 and not w7647;
w7649 <= not w7610 and w7648;
w7650 <= not w7610 and not w7649;
w7651 <= w7648 and not w7649;
w7652 <= not w7650 and not w7651;
w7653 <= not w7609 and not w7652;
w7654 <= w7609 and not w7651;
w7655 <= not w7650 and w7654;
w7656 <= not w7653 and not w7655;
w7657 <= not w7392 and w7656;
w7658 <= w7392 and not w7656;
w7659 <= not w7657 and not w7658;
w7660 <= not w7385 and not w7388;
w7661 <= not w7384 and not w7660;
w7662 <= not w7659 and w7661;
w7663 <= w7659 and not w7661;
w7664 <= not w7662 and not w7663;
w7665 <= not w7658 and not w7661;
w7666 <= not w7657 and not w7665;
w7667 <= not w7649 and not w7653;
w7668 <= not w7432 and not w7606;
w7669 <= not w7405 and not w7428;
w7670 <= not w7443 and not w7494;
w7671 <= not w7436 and not w7439;
w7672 <= not w7416 and not w7420;
w7673 <= w7671 and w7672;
w7674 <= not w7671 and not w7672;
w7675 <= not w7673 and not w7674;
w7676 <= not w7410 and not w7413;
w7677 <= not w7675 and w7676;
w7678 <= w7675 and not w7676;
w7679 <= not w7677 and not w7678;
w7680 <= not w7422 and not w7425;
w7681 <= w7679 and not w7680;
w7682 <= not w7679 and w7680;
w7683 <= not w7681 and not w7682;
w7684 <= not w7670 and w7683;
w7685 <= w7670 and not w7683;
w7686 <= not w7684 and not w7685;
w7687 <= w7669 and not w7686;
w7688 <= not w7669 and w7686;
w7689 <= not w7687 and not w7688;
w7690 <= not w7501 and w7602;
w7691 <= not w7497 and not w7690;
w7692 <= w7689 and not w7691;
w7693 <= not w7689 and w7691;
w7694 <= not w7692 and not w7693;
w7695 <= w7668 and not w7694;
w7696 <= not w7668 and w7694;
w7697 <= not w7695 and not w7696;
w7698 <= not w7643 and not w7646;
w7699 <= not w7598 and not w7600;
w7700 <= not w7574 and not w7593;
w7701 <= not w7531 and not w7547;
w7702 <= a(1) and a(57);
w7703 <= w2916 and w7702;
w7704 <= not w2916 and not w7702;
w7705 <= not w7703 and not w7704;
w7706 <= not w7624 and not w7705;
w7707 <= w7624 and w7705;
w7708 <= not w7706 and not w7707;
w7709 <= not w7571 and w7708;
w7710 <= w7571 and not w7708;
w7711 <= not w7709 and not w7710;
w7712 <= not w7701 and w7711;
w7713 <= not w7701 and not w7712;
w7714 <= w7711 and not w7712;
w7715 <= not w7713 and not w7714;
w7716 <= not w7700 and not w7715;
w7717 <= w7700 and not w7714;
w7718 <= not w7713 and w7717;
w7719 <= not w7716 and not w7718;
w7720 <= not w7699 and w7719;
w7721 <= w7699 and not w7719;
w7722 <= not w7720 and not w7721;
w7723 <= not w7473 and not w7490;
w7724 <= w7484 and w7544;
w7725 <= not w7484 and not w7544;
w7726 <= not w7724 and not w7725;
w7727 <= w7470 and not w7726;
w7728 <= not w7470 and w7726;
w7729 <= not w7727 and not w7728;
w7730 <= w7511 and w7528;
w7731 <= not w7511 and not w7528;
w7732 <= not w7730 and not w7731;
w7733 <= w7559 and not w7732;
w7734 <= not w7559 and w7732;
w7735 <= not w7733 and not w7734;
w7736 <= w7729 and w7735;
w7737 <= not w7729 and not w7735;
w7738 <= not w7736 and not w7737;
w7739 <= not w7723 and w7738;
w7740 <= w7723 and not w7738;
w7741 <= not w7739 and not w7740;
w7742 <= w7722 and w7741;
w7743 <= not w7722 and not w7741;
w7744 <= not w7742 and not w7743;
w7745 <= w7698 and not w7744;
w7746 <= not w7698 and w7744;
w7747 <= not w7745 and not w7746;
w7748 <= a(56) and a(58);
w7749 <= w2 and w7748;
w7750 <= w58 and w7227;
w7751 <= not w7749 and not w7750;
w7752 <= a(0) and a(58);
w7753 <= a(4) and a(54);
w7754 <= w7752 and w7753;
w7755 <= not w7751 and not w7754;
w7756 <= not w7754 and not w7755;
w7757 <= not w7752 and not w7753;
w7758 <= w7756 and not w7757;
w7759 <= a(2) and a(56);
w7760 <= not w7755 and w7759;
w7761 <= not w7758 and not w7760;
w7762 <= a(20) and a(38);
w7763 <= a(21) and a(37);
w7764 <= not w7762 and not w7763;
w7765 <= w1300 and w4371;
w7766 <= a(5) and not w7765;
w7767 <= a(53) and w7766;
w7768 <= not w7764 and w7767;
w7769 <= a(53) and not w7768;
w7770 <= a(5) and w7769;
w7771 <= not w7765 and not w7768;
w7772 <= not w7764 and w7771;
w7773 <= not w7770 and not w7772;
w7774 <= not w7761 and not w7773;
w7775 <= not w7761 and not w7774;
w7776 <= not w7773 and not w7774;
w7777 <= not w7775 and not w7776;
w7778 <= a(42) and a(49);
w7779 <= w653 and w7778;
w7780 <= w854 and w5150;
w7781 <= w5762 and w6869;
w7782 <= not w7780 and not w7781;
w7783 <= not w7779 and not w7782;
w7784 <= a(41) and not w7783;
w7785 <= a(17) and w7784;
w7786 <= a(9) and a(49);
w7787 <= a(16) and a(42);
w7788 <= not w7786 and not w7787;
w7789 <= not w7779 and not w7783;
w7790 <= not w7788 and w7789;
w7791 <= not w7785 and not w7790;
w7792 <= not w7777 and not w7791;
w7793 <= not w7777 and not w7792;
w7794 <= not w7791 and not w7792;
w7795 <= not w7793 and not w7794;
w7796 <= a(7) and a(51);
w7797 <= a(8) and a(50);
w7798 <= not w7796 and not w7797;
w7799 <= w186 and w6370;
w7800 <= a(40) and not w7799;
w7801 <= a(18) and w7800;
w7802 <= not w7798 and w7801;
w7803 <= not w7799 and not w7802;
w7804 <= not w7798 and w7803;
w7805 <= a(40) and not w7802;
w7806 <= a(18) and w7805;
w7807 <= not w7804 and not w7806;
w7808 <= w1472 and w3125;
w7809 <= w1921 and w4401;
w7810 <= w1725 and w3634;
w7811 <= not w7809 and not w7810;
w7812 <= not w7808 and not w7811;
w7813 <= a(36) and not w7812;
w7814 <= a(22) and w7813;
w7815 <= not w7808 and not w7812;
w7816 <= a(23) and a(35);
w7817 <= a(24) and a(34);
w7818 <= not w7816 and not w7817;
w7819 <= w7815 and not w7818;
w7820 <= not w7814 and not w7819;
w7821 <= not w7807 and not w7820;
w7822 <= not w7807 and not w7821;
w7823 <= not w7820 and not w7821;
w7824 <= not w7822 and not w7823;
w7825 <= w2033 and w3618;
w7826 <= w2404 and w2439;
w7827 <= w2269 and w2949;
w7828 <= not w7826 and not w7827;
w7829 <= not w7825 and not w7828;
w7830 <= w3107 and not w7829;
w7831 <= not w7825 and not w7829;
w7832 <= a(27) and a(31);
w7833 <= not w3072 and not w7832;
w7834 <= w7831 and not w7833;
w7835 <= not w7830 and not w7834;
w7836 <= not w7824 and not w7835;
w7837 <= not w7824 and not w7836;
w7838 <= not w7835 and not w7836;
w7839 <= not w7837 and not w7838;
w7840 <= not w7795 and w7839;
w7841 <= w7795 and not w7839;
w7842 <= not w7840 and not w7841;
w7843 <= not w7397 and not w7401;
w7844 <= w7842 and w7843;
w7845 <= not w7842 and not w7843;
w7846 <= not w7844 and not w7845;
w7847 <= not w7616 and not w7640;
w7848 <= w7452 and w7587;
w7849 <= not w7452 and not w7587;
w7850 <= not w7848 and not w7849;
w7851 <= not w7619 and not w7628;
w7852 <= not w7850 and w7851;
w7853 <= w7850 and not w7851;
w7854 <= not w7852 and not w7853;
w7855 <= not w7634 and not w7638;
w7856 <= not w7854 and w7855;
w7857 <= w7854 and not w7855;
w7858 <= not w7856 and not w7857;
w7859 <= a(43) and a(47);
w7860 <= w622 and w7859;
w7861 <= w529 and w6058;
w7862 <= w6465 and w7157;
w7863 <= not w7861 and not w7862;
w7864 <= not w7860 and not w7863;
w7865 <= not w7860 and not w7864;
w7866 <= a(11) and a(47);
w7867 <= not w5453 and not w7866;
w7868 <= w7865 and not w7867;
w7869 <= a(48) and not w7864;
w7870 <= a(10) and w7869;
w7871 <= not w7868 and not w7870;
w7872 <= w554 and w5366;
w7873 <= w412 and w7553;
w7874 <= w551 and w5519;
w7875 <= not w7873 and not w7874;
w7876 <= not w7872 and not w7875;
w7877 <= w6427 and not w7876;
w7878 <= not w7872 and not w7876;
w7879 <= a(12) and a(46);
w7880 <= not w6992 and not w7879;
w7881 <= w7878 and not w7880;
w7882 <= not w7877 and not w7881;
w7883 <= not w7871 and not w7882;
w7884 <= not w7871 and not w7883;
w7885 <= not w7882 and not w7883;
w7886 <= not w7884 and not w7885;
w7887 <= a(6) and a(52);
w7888 <= a(19) and a(39);
w7889 <= not w7887 and not w7888;
w7890 <= w7887 and w7888;
w7891 <= a(3) and not w7890;
w7892 <= a(55) and w7891;
w7893 <= not w7889 and w7892;
w7894 <= a(55) and not w7893;
w7895 <= a(3) and w7894;
w7896 <= not w7890 and not w7893;
w7897 <= not w7889 and w7896;
w7898 <= not w7895 and not w7897;
w7899 <= not w7886 and not w7898;
w7900 <= not w7886 and not w7899;
w7901 <= not w7898 and not w7899;
w7902 <= not w7900 and not w7901;
w7903 <= not w7858 and w7902;
w7904 <= w7858 and not w7902;
w7905 <= not w7903 and not w7904;
w7906 <= not w7847 and w7905;
w7907 <= not w7847 and not w7906;
w7908 <= w7905 and not w7906;
w7909 <= not w7907 and not w7908;
w7910 <= w7846 and not w7909;
w7911 <= w7846 and not w7910;
w7912 <= not w7909 and not w7910;
w7913 <= not w7911 and not w7912;
w7914 <= w7747 and not w7913;
w7915 <= w7747 and not w7914;
w7916 <= not w7913 and not w7914;
w7917 <= not w7915 and not w7916;
w7918 <= not w7697 and w7917;
w7919 <= w7697 and not w7917;
w7920 <= not w7918 and not w7919;
w7921 <= not w7667 and w7920;
w7922 <= w7667 and not w7920;
w7923 <= not w7921 and not w7922;
w7924 <= w7666 and not w7923;
w7925 <= not w7666 and not w7922;
w7926 <= not w7921 and w7925;
w7927 <= not w7924 and not w7926;
w7928 <= not w7746 and not w7914;
w7929 <= not w7906 and not w7910;
w7930 <= not w7720 and not w7742;
w7931 <= not w7857 and not w7904;
w7932 <= not w7849 and not w7853;
w7933 <= not w7731 and not w7734;
w7934 <= w7932 and w7933;
w7935 <= not w7932 and not w7933;
w7936 <= not w7934 and not w7935;
w7937 <= not w7725 and not w7728;
w7938 <= not w7936 and w7937;
w7939 <= w7936 and not w7937;
w7940 <= not w7938 and not w7939;
w7941 <= not w7736 and not w7739;
w7942 <= w7940 and not w7941;
w7943 <= not w7940 and w7941;
w7944 <= not w7942 and not w7943;
w7945 <= not w7931 and w7944;
w7946 <= w7931 and not w7944;
w7947 <= not w7945 and not w7946;
w7948 <= not w7930 and w7947;
w7949 <= w7930 and not w7947;
w7950 <= not w7948 and not w7949;
w7951 <= not w7929 and w7950;
w7952 <= w7929 and not w7950;
w7953 <= not w7951 and not w7952;
w7954 <= w7928 and not w7953;
w7955 <= not w7928 and w7953;
w7956 <= not w7954 and not w7955;
w7957 <= not w7681 and not w7684;
w7958 <= not w7712 and not w7716;
w7959 <= w412 and w5056;
w7960 <= w408 and w6058;
w7961 <= a(45) and a(48);
w7962 <= w1411 and w7961;
w7963 <= not w7960 and not w7962;
w7964 <= not w7959 and not w7963;
w7965 <= not w7959 and not w7964;
w7966 <= a(12) and a(47);
w7967 <= a(14) and a(45);
w7968 <= not w7966 and not w7967;
w7969 <= w7965 and not w7968;
w7970 <= a(48) and not w7964;
w7971 <= a(11) and w7970;
w7972 <= not w7969 and not w7971;
w7973 <= a(13) and a(46);
w7974 <= a(28) and a(31);
w7975 <= not w2423 and not w7974;
w7976 <= w2423 and w7974;
w7977 <= w7973 and not w7976;
w7978 <= not w7975 and w7977;
w7979 <= w7973 and not w7978;
w7980 <= not w7976 and not w7978;
w7981 <= not w7975 and w7980;
w7982 <= not w7979 and not w7981;
w7983 <= not w7972 and not w7982;
w7984 <= not w7972 and not w7983;
w7985 <= not w7982 and not w7983;
w7986 <= not w7984 and not w7985;
w7987 <= a(16) and a(43);
w7988 <= a(17) and a(42);
w7989 <= not w7987 and not w7988;
w7990 <= w854 and w4824;
w7991 <= a(8) and not w7990;
w7992 <= a(51) and w7991;
w7993 <= not w7989 and w7992;
w7994 <= a(51) and not w7993;
w7995 <= a(8) and w7994;
w7996 <= not w7990 and not w7993;
w7997 <= not w7989 and w7996;
w7998 <= not w7995 and not w7997;
w7999 <= not w7986 and not w7998;
w8000 <= not w7986 and not w7999;
w8001 <= not w7998 and not w7999;
w8002 <= not w8000 and not w8001;
w8003 <= a(2) and a(57);
w8004 <= a(3) and a(56);
w8005 <= not w8003 and not w8004;
w8006 <= a(56) and a(57);
w8007 <= w24 and w8006;
w8008 <= not w8005 and not w8007;
w8009 <= w7703 and w8008;
w8010 <= not w8007 and not w8009;
w8011 <= not w8005 and w8010;
w8012 <= w7703 and not w8009;
w8013 <= not w8011 and not w8012;
w8014 <= w7831 and not w8013;
w8015 <= not w7831 and w8013;
w8016 <= not w8014 and not w8015;
w8017 <= w32 and w7507;
w8018 <= a(19) and a(55);
w8019 <= w4389 and w8018;
w8020 <= not w8017 and not w8019;
w8021 <= a(5) and a(54);
w8022 <= a(19) and a(40);
w8023 <= w8021 and w8022;
w8024 <= not w8020 and not w8023;
w8025 <= a(55) and not w8024;
w8026 <= a(4) and w8025;
w8027 <= not w8023 and not w8024;
w8028 <= not w8021 and not w8022;
w8029 <= w8027 and not w8028;
w8030 <= not w8026 and not w8029;
w8031 <= not w8016 and not w8030;
w8032 <= w8016 and w8030;
w8033 <= not w8031 and not w8032;
w8034 <= w8002 and not w8033;
w8035 <= not w8002 and w8033;
w8036 <= not w8034 and not w8035;
w8037 <= not w7958 and w8036;
w8038 <= w7958 and not w8036;
w8039 <= not w8037 and not w8038;
w8040 <= w7957 and not w8039;
w8041 <= not w7957 and w8039;
w8042 <= not w8040 and not w8041;
w8043 <= a(18) and a(52);
w8044 <= w5217 and w8043;
w8045 <= a(41) and a(53);
w8046 <= w1284 and w8045;
w8047 <= w141 and w7239;
w8048 <= not w8046 and not w8047;
w8049 <= not w8044 and not w8048;
w8050 <= not w8044 and not w8049;
w8051 <= a(7) and a(52);
w8052 <= a(18) and a(41);
w8053 <= not w8051 and not w8052;
w8054 <= w8050 and not w8053;
w8055 <= a(53) and not w8049;
w8056 <= a(6) and w8055;
w8057 <= not w8054 and not w8056;
w8058 <= a(44) and a(49);
w8059 <= w491 and w8058;
w8060 <= a(44) and a(50);
w8061 <= w1323 and w8060;
w8062 <= w290 and w6131;
w8063 <= not w8061 and not w8062;
w8064 <= not w8059 and not w8063;
w8065 <= a(50) and not w8064;
w8066 <= a(9) and w8065;
w8067 <= a(10) and a(49);
w8068 <= not w5104 and not w8067;
w8069 <= not w8059 and not w8064;
w8070 <= not w8068 and w8069;
w8071 <= not w8066 and not w8070;
w8072 <= not w8057 and not w8071;
w8073 <= not w8057 and not w8072;
w8074 <= not w8071 and not w8072;
w8075 <= not w8073 and not w8074;
w8076 <= not w7707 and not w7709;
w8077 <= w8075 and w8076;
w8078 <= not w8075 and not w8076;
w8079 <= not w8077 and not w8078;
w8080 <= not w7674 and not w7678;
w8081 <= not w8079 and w8080;
w8082 <= w8079 and not w8080;
w8083 <= not w8081 and not w8082;
w8084 <= w1380 and w4371;
w8085 <= w1499 and w5236;
w8086 <= w1300 and w4889;
w8087 <= not w8085 and not w8086;
w8088 <= not w8084 and not w8087;
w8089 <= not w8084 and not w8088;
w8090 <= a(21) and a(38);
w8091 <= a(22) and a(37);
w8092 <= not w8090 and not w8091;
w8093 <= w8089 and not w8092;
w8094 <= a(39) and not w8088;
w8095 <= a(20) and w8094;
w8096 <= not w8093 and not w8095;
w8097 <= w1710 and w3125;
w8098 <= w1353 and w4401;
w8099 <= w1472 and w3634;
w8100 <= not w8098 and not w8099;
w8101 <= not w8097 and not w8100;
w8102 <= a(36) and not w8101;
w8103 <= a(23) and w8102;
w8104 <= a(24) and a(35);
w8105 <= a(25) and a(34);
w8106 <= not w8104 and not w8105;
w8107 <= not w8097 and not w8101;
w8108 <= not w8106 and w8107;
w8109 <= not w8103 and not w8108;
w8110 <= not w8096 and not w8109;
w8111 <= not w8096 and not w8110;
w8112 <= not w8109 and not w8110;
w8113 <= not w8111 and not w8112;
w8114 <= a(32) and a(59);
w8115 <= w1618 and w8114;
w8116 <= w2033 and w2949;
w8117 <= a(26) and a(59);
w8118 <= w2411 and w8117;
w8119 <= not w8116 and not w8118;
w8120 <= not w8115 and not w8119;
w8121 <= a(33) and not w8120;
w8122 <= a(26) and w8121;
w8123 <= not w8115 and not w8120;
w8124 <= a(0) and a(59);
w8125 <= a(27) and a(32);
w8126 <= not w8124 and not w8125;
w8127 <= w8123 and not w8126;
w8128 <= not w8122 and not w8127;
w8129 <= not w8113 and not w8128;
w8130 <= not w8113 and not w8129;
w8131 <= not w8128 and not w8129;
w8132 <= not w8130 and not w8131;
w8133 <= w8083 and not w8132;
w8134 <= not w8083 and w8132;
w8135 <= w8042 and not w8134;
w8136 <= not w8133 and w8135;
w8137 <= w8042 and not w8136;
w8138 <= not w8134 and not w8136;
w8139 <= not w8133 and w8138;
w8140 <= not w8137 and not w8139;
w8141 <= not w7688 and not w7692;
w8142 <= not w7883 and not w7899;
w8143 <= not w7821 and not w7836;
w8144 <= w8142 and w8143;
w8145 <= not w8142 and not w8143;
w8146 <= not w8144 and not w8145;
w8147 <= not w7774 and not w7792;
w8148 <= not w8146 and w8147;
w8149 <= w8146 and not w8147;
w8150 <= not w8148 and not w8149;
w8151 <= not w7795 and not w7839;
w8152 <= not w7845 and not w8151;
w8153 <= w7756 and w7896;
w8154 <= not w7756 and not w7896;
w8155 <= not w8153 and not w8154;
w8156 <= w7789 and not w8155;
w8157 <= not w7789 and w8155;
w8158 <= not w8156 and not w8157;
w8159 <= w7771 and w7815;
w8160 <= not w7771 and not w7815;
w8161 <= not w8159 and not w8160;
w8162 <= w7803 and not w8161;
w8163 <= not w7803 and w8161;
w8164 <= not w8162 and not w8163;
w8165 <= a(58) and w2208;
w8166 <= a(1) and a(58);
w8167 <= not a(30) and not w8166;
w8168 <= not w8165 and not w8167;
w8169 <= w7878 and not w8168;
w8170 <= not w7878 and w8168;
w8171 <= not w8169 and not w8170;
w8172 <= not w7865 and w8171;
w8173 <= w7865 and not w8171;
w8174 <= not w8172 and not w8173;
w8175 <= w8164 and w8174;
w8176 <= w8164 and not w8175;
w8177 <= w8174 and not w8175;
w8178 <= not w8176 and not w8177;
w8179 <= w8158 and not w8178;
w8180 <= not w8158 and not w8177;
w8181 <= not w8176 and w8180;
w8182 <= not w8179 and not w8181;
w8183 <= not w8152 and w8182;
w8184 <= not w8152 and not w8183;
w8185 <= w8182 and not w8183;
w8186 <= not w8184 and not w8185;
w8187 <= w8150 and not w8186;
w8188 <= not w8150 and not w8185;
w8189 <= not w8184 and w8188;
w8190 <= not w8187 and not w8189;
w8191 <= not w8141 and w8190;
w8192 <= w8141 and not w8190;
w8193 <= not w8191 and not w8192;
w8194 <= not w8140 and w8193;
w8195 <= w8140 and not w8193;
w8196 <= not w8194 and not w8195;
w8197 <= w7956 and w8196;
w8198 <= not w7956 and not w8196;
w8199 <= not w8197 and not w8198;
w8200 <= not w7696 and not w7919;
w8201 <= not w8199 and w8200;
w8202 <= w8199 and not w8200;
w8203 <= not w8201 and not w8202;
w8204 <= not w7921 and not w7925;
w8205 <= not w8203 and w8204;
w8206 <= w8203 and not w8204;
w8207 <= not w8205 and not w8206;
w8208 <= not w7955 and not w8197;
w8209 <= not w8191 and not w8194;
w8210 <= not w8041 and not w8136;
w8211 <= not w8183 and not w8187;
w8212 <= not w8160 and not w8163;
w8213 <= not w8154 and not w8157;
w8214 <= w8212 and w8213;
w8215 <= not w8212 and not w8213;
w8216 <= not w8214 and not w8215;
w8217 <= not w7831 and not w8013;
w8218 <= not w8031 and not w8217;
w8219 <= not w8216 and w8218;
w8220 <= w8216 and not w8218;
w8221 <= not w8219 and not w8220;
w8222 <= not w8145 and not w8149;
w8223 <= not w8221 and w8222;
w8224 <= w8221 and not w8222;
w8225 <= not w8223 and not w8224;
w8226 <= not w8082 and not w8133;
w8227 <= w8225 and not w8226;
w8228 <= not w8225 and w8226;
w8229 <= not w8227 and not w8228;
w8230 <= not w8211 and w8229;
w8231 <= w8211 and not w8229;
w8232 <= not w8230 and not w8231;
w8233 <= not w8210 and w8232;
w8234 <= w8210 and not w8232;
w8235 <= not w8233 and not w8234;
w8236 <= w8209 and not w8235;
w8237 <= not w8209 and w8235;
w8238 <= not w8236 and not w8237;
w8239 <= not w7942 and not w7945;
w8240 <= w15 and w8006;
w8241 <= w58 and w7748;
w8242 <= a(57) and a(58);
w8243 <= w24 and w8242;
w8244 <= not w8241 and not w8243;
w8245 <= not w8240 and not w8244;
w8246 <= not w8240 and not w8245;
w8247 <= a(3) and a(57);
w8248 <= a(4) and a(56);
w8249 <= not w8247 and not w8248;
w8250 <= w8246 and not w8249;
w8251 <= a(58) and not w8245;
w8252 <= a(2) and w8251;
w8253 <= not w8250 and not w8252;
w8254 <= w1380 and w4889;
w8255 <= w1499 and w3609;
w8256 <= w1300 and w3977;
w8257 <= not w8255 and not w8256;
w8258 <= not w8254 and not w8257;
w8259 <= a(40) and not w8258;
w8260 <= a(20) and w8259;
w8261 <= a(21) and a(39);
w8262 <= a(22) and a(38);
w8263 <= not w8261 and not w8262;
w8264 <= not w8254 and not w8258;
w8265 <= not w8263 and w8264;
w8266 <= not w8260 and not w8265;
w8267 <= not w8253 and not w8266;
w8268 <= not w8253 and not w8267;
w8269 <= not w8266 and not w8267;
w8270 <= not w8268 and not w8269;
w8271 <= w2269 and w3125;
w8272 <= w2107 and w4401;
w8273 <= w1710 and w3634;
w8274 <= not w8272 and not w8273;
w8275 <= not w8271 and not w8274;
w8276 <= a(36) and not w8275;
w8277 <= a(24) and w8276;
w8278 <= not w8271 and not w8275;
w8279 <= a(25) and a(35);
w8280 <= a(26) and a(34);
w8281 <= not w8279 and not w8280;
w8282 <= w8278 and not w8281;
w8283 <= not w8277 and not w8282;
w8284 <= not w8270 and not w8283;
w8285 <= not w8270 and not w8284;
w8286 <= not w8283 and not w8284;
w8287 <= not w8285 and not w8286;
w8288 <= not w7935 and not w7939;
w8289 <= w8287 and w8288;
w8290 <= not w8287 and not w8288;
w8291 <= not w8289 and not w8290;
w8292 <= a(44) and a(51);
w8293 <= w653 and w8292;
w8294 <= w854 and w5102;
w8295 <= w6322 and w7578;
w8296 <= not w8294 and not w8295;
w8297 <= not w8293 and not w8296;
w8298 <= a(43) and not w8297;
w8299 <= a(17) and w8298;
w8300 <= not w8293 and not w8297;
w8301 <= a(9) and a(51);
w8302 <= a(16) and a(44);
w8303 <= not w8301 and not w8302;
w8304 <= w8300 and not w8303;
w8305 <= not w8299 and not w8304;
w8306 <= w7965 and not w8305;
w8307 <= not w7965 and w8305;
w8308 <= not w8306 and not w8307;
w8309 <= a(45) and a(49);
w8310 <= w622 and w8309;
w8311 <= w529 and w6131;
w8312 <= a(45) and a(50);
w8313 <= w491 and w8312;
w8314 <= not w8311 and not w8313;
w8315 <= not w8310 and not w8314;
w8316 <= a(50) and not w8315;
w8317 <= a(10) and w8316;
w8318 <= a(11) and a(49);
w8319 <= a(15) and a(45);
w8320 <= not w8318 and not w8319;
w8321 <= not w8310 and not w8315;
w8322 <= not w8320 and w8321;
w8323 <= not w8317 and not w8322;
w8324 <= not w8308 and not w8323;
w8325 <= w8308 and w8323;
w8326 <= not w8324 and not w8325;
w8327 <= not w8291 and not w8326;
w8328 <= w8291 and w8326;
w8329 <= not w8327 and not w8328;
w8330 <= not w8239 and w8329;
w8331 <= not w8239 and not w8330;
w8332 <= w8329 and not w8330;
w8333 <= not w8331 and not w8332;
w8334 <= not w8175 and not w8179;
w8335 <= a(0) and a(60);
w8336 <= w8165 and w8335;
w8337 <= w8165 and not w8336;
w8338 <= not w8165 and w8335;
w8339 <= not w8337 and not w8338;
w8340 <= a(1) and a(59);
w8341 <= w3258 and w8340;
w8342 <= w8340 and not w8341;
w8343 <= w3258 and not w8341;
w8344 <= not w8342 and not w8343;
w8345 <= not w8339 and not w8344;
w8346 <= not w8339 and not w8345;
w8347 <= not w8344 and not w8345;
w8348 <= not w8346 and not w8347;
w8349 <= w2137 and w2949;
w8350 <= w3865 and w7183;
w8351 <= not w8349 and not w8350;
w8352 <= a(23) and a(37);
w8353 <= w5669 and w8352;
w8354 <= not w8351 and not w8353;
w8355 <= a(33) and not w8354;
w8356 <= a(27) and w8355;
w8357 <= not w8353 and not w8354;
w8358 <= not w5669 and not w8352;
w8359 <= w8357 and not w8358;
w8360 <= not w8356 and not w8359;
w8361 <= not w8348 and not w8360;
w8362 <= not w8348 and not w8361;
w8363 <= not w8360 and not w8361;
w8364 <= not w8362 and not w8363;
w8365 <= not w8170 and not w8172;
w8366 <= w8364 and w8365;
w8367 <= not w8364 and not w8365;
w8368 <= not w8366 and not w8367;
w8369 <= w186 and w7239;
w8370 <= a(18) and a(53);
w8371 <= w5425 and w8370;
w8372 <= not w8369 and not w8371;
w8373 <= a(8) and a(52);
w8374 <= a(18) and a(42);
w8375 <= w8373 and w8374;
w8376 <= not w8372 and not w8375;
w8377 <= not w8375 and not w8376;
w8378 <= not w8373 and not w8374;
w8379 <= w8377 and not w8378;
w8380 <= a(53) and not w8376;
w8381 <= a(7) and w8380;
w8382 <= not w8379 and not w8381;
w8383 <= w554 and w6058;
w8384 <= a(46) and a(48);
w8385 <= w412 and w8384;
w8386 <= w551 and w5472;
w8387 <= not w8385 and not w8386;
w8388 <= not w8383 and not w8387;
w8389 <= w7206 and not w8388;
w8390 <= not w8383 and not w8388;
w8391 <= a(12) and a(48);
w8392 <= a(13) and a(47);
w8393 <= not w8391 and not w8392;
w8394 <= w8390 and not w8393;
w8395 <= not w8389 and not w8394;
w8396 <= not w8382 and not w8395;
w8397 <= not w8382 and not w8396;
w8398 <= not w8395 and not w8396;
w8399 <= not w8397 and not w8398;
w8400 <= a(41) and a(55);
w8401 <= w1308 and w8400;
w8402 <= w138 and w7507;
w8403 <= not w8401 and not w8402;
w8404 <= a(6) and a(54);
w8405 <= a(19) and a(41);
w8406 <= w8404 and w8405;
w8407 <= not w8403 and not w8406;
w8408 <= a(55) and not w8407;
w8409 <= a(5) and w8408;
w8410 <= not w8406 and not w8407;
w8411 <= not w8404 and not w8405;
w8412 <= w8410 and not w8411;
w8413 <= not w8409 and not w8412;
w8414 <= not w8399 and not w8413;
w8415 <= not w8399 and not w8414;
w8416 <= not w8413 and not w8414;
w8417 <= not w8415 and not w8416;
w8418 <= not w8368 and w8417;
w8419 <= w8368 and not w8417;
w8420 <= not w8418 and not w8419;
w8421 <= not w8334 and w8420;
w8422 <= w8334 and not w8420;
w8423 <= not w8421 and not w8422;
w8424 <= not w8333 and w8423;
w8425 <= w8423 and not w8424;
w8426 <= not w8333 and not w8424;
w8427 <= not w8425 and not w8426;
w8428 <= not w7948 and not w7951;
w8429 <= w7996 and w8050;
w8430 <= not w7996 and not w8050;
w8431 <= not w8429 and not w8430;
w8432 <= w7980 and not w8431;
w8433 <= not w7980 and w8431;
w8434 <= not w8432 and not w8433;
w8435 <= not w8110 and not w8129;
w8436 <= not w8434 and w8435;
w8437 <= w8434 and not w8435;
w8438 <= not w8436 and not w8437;
w8439 <= not w7983 and not w7999;
w8440 <= not w8438 and w8439;
w8441 <= w8438 and not w8439;
w8442 <= not w8440 and not w8441;
w8443 <= not w8035 and not w8037;
w8444 <= not w8072 and not w8078;
w8445 <= w8027 and w8089;
w8446 <= not w8027 and not w8089;
w8447 <= not w8445 and not w8446;
w8448 <= w8107 and not w8447;
w8449 <= not w8107 and w8447;
w8450 <= not w8448 and not w8449;
w8451 <= w8010 and w8123;
w8452 <= not w8010 and not w8123;
w8453 <= not w8451 and not w8452;
w8454 <= w8069 and not w8453;
w8455 <= not w8069 and w8453;
w8456 <= not w8454 and not w8455;
w8457 <= w8450 and w8456;
w8458 <= not w8450 and not w8456;
w8459 <= not w8457 and not w8458;
w8460 <= not w8444 and w8459;
w8461 <= w8444 and not w8459;
w8462 <= not w8460 and not w8461;
w8463 <= not w8443 and w8462;
w8464 <= not w8443 and not w8463;
w8465 <= w8462 and not w8463;
w8466 <= not w8464 and not w8465;
w8467 <= w8442 and not w8466;
w8468 <= not w8442 and not w8465;
w8469 <= not w8464 and w8468;
w8470 <= not w8467 and not w8469;
w8471 <= not w8428 and w8470;
w8472 <= not w8428 and not w8471;
w8473 <= w8470 and not w8471;
w8474 <= not w8472 and not w8473;
w8475 <= not w8427 and not w8474;
w8476 <= w8427 and not w8473;
w8477 <= not w8472 and w8476;
w8478 <= not w8475 and not w8477;
w8479 <= w8238 and w8478;
w8480 <= not w8238 and not w8478;
w8481 <= not w8479 and not w8480;
w8482 <= w8208 and not w8481;
w8483 <= not w8208 and w8481;
w8484 <= not w8482 and not w8483;
w8485 <= not w8201 and not w8204;
w8486 <= not w8202 and not w8485;
w8487 <= not w8484 and w8486;
w8488 <= w8484 and not w8486;
w8489 <= not w8487 and not w8488;
w8490 <= not w8237 and not w8479;
w8491 <= not w8471 and not w8475;
w8492 <= not w8330 and not w8424;
w8493 <= not w8437 and not w8441;
w8494 <= a(7) and a(54);
w8495 <= a(8) and a(53);
w8496 <= not w8494 and not w8495;
w8497 <= w186 and w7505;
w8498 <= a(42) and not w8497;
w8499 <= a(19) and w8498;
w8500 <= not w8496 and w8499;
w8501 <= not w8497 and not w8500;
w8502 <= not w8496 and w8501;
w8503 <= a(42) and not w8500;
w8504 <= a(19) and w8503;
w8505 <= not w8502 and not w8504;
w8506 <= a(44) and a(52);
w8507 <= w1482 and w8506;
w8508 <= w6322 and w8043;
w8509 <= w858 and w5102;
w8510 <= not w8508 and not w8509;
w8511 <= not w8507 and not w8510;
w8512 <= a(43) and not w8511;
w8513 <= a(18) and w8512;
w8514 <= not w8507 and not w8511;
w8515 <= a(9) and a(52);
w8516 <= a(17) and a(44);
w8517 <= not w8515 and not w8516;
w8518 <= w8514 and not w8517;
w8519 <= not w8513 and not w8518;
w8520 <= not w8505 and not w8519;
w8521 <= not w8505 and not w8520;
w8522 <= not w8519 and not w8520;
w8523 <= not w8521 and not w8522;
w8524 <= w2137 and w3956;
w8525 <= w2606 and w2778;
w8526 <= w2033 and w3125;
w8527 <= not w8525 and not w8526;
w8528 <= not w8524 and not w8527;
w8529 <= a(35) and not w8528;
w8530 <= a(26) and w8529;
w8531 <= not w8524 and not w8528;
w8532 <= a(28) and a(33);
w8533 <= not w3309 and not w8532;
w8534 <= w8531 and not w8533;
w8535 <= not w8530 and not w8534;
w8536 <= not w8523 and not w8535;
w8537 <= not w8523 and not w8536;
w8538 <= not w8535 and not w8536;
w8539 <= not w8537 and not w8538;
w8540 <= not w8457 and not w8460;
w8541 <= not w8539 and not w8540;
w8542 <= not w8539 and not w8541;
w8543 <= not w8540 and not w8541;
w8544 <= not w8542 and not w8543;
w8545 <= not w8493 and not w8544;
w8546 <= not w8493 and not w8545;
w8547 <= not w8544 and not w8545;
w8548 <= not w8546 and not w8547;
w8549 <= not w8290 and not w8328;
w8550 <= not w8452 and not w8455;
w8551 <= not w8430 and not w8433;
w8552 <= a(3) and a(58);
w8553 <= a(4) and a(57);
w8554 <= not w8552 and not w8553;
w8555 <= w15 and w8242;
w8556 <= a(38) and not w8555;
w8557 <= a(23) and w8556;
w8558 <= not w8554 and w8557;
w8559 <= a(38) and not w8558;
w8560 <= a(23) and w8559;
w8561 <= not w8555 and not w8558;
w8562 <= not w8554 and w8561;
w8563 <= not w8560 and not w8562;
w8564 <= not w8551 and not w8563;
w8565 <= not w8551 and not w8564;
w8566 <= not w8563 and not w8564;
w8567 <= not w8565 and not w8566;
w8568 <= not w8550 and not w8567;
w8569 <= not w8550 and not w8568;
w8570 <= not w8567 and not w8568;
w8571 <= not w8569 and not w8570;
w8572 <= not w7965 and not w8305;
w8573 <= not w8324 and not w8572;
w8574 <= not w8446 and not w8449;
w8575 <= a(1) and a(60);
w8576 <= a(31) and w8575;
w8577 <= not a(31) and not w8575;
w8578 <= not w8576 and not w8577;
w8579 <= w8341 and w8578;
w8580 <= not w8341 and not w8578;
w8581 <= not w8579 and not w8580;
w8582 <= not w8390 and w8581;
w8583 <= w8390 and not w8581;
w8584 <= not w8582 and not w8583;
w8585 <= not w8574 and w8584;
w8586 <= w8574 and not w8584;
w8587 <= not w8585 and not w8586;
w8588 <= not w8573 and w8587;
w8589 <= w8573 and not w8587;
w8590 <= not w8588 and not w8589;
w8591 <= not w8571 and w8590;
w8592 <= not w8571 and not w8591;
w8593 <= w8590 and not w8591;
w8594 <= not w8592 and not w8593;
w8595 <= not w8549 and not w8594;
w8596 <= w8549 and not w8593;
w8597 <= not w8592 and w8596;
w8598 <= not w8595 and not w8597;
w8599 <= not w8548 and w8598;
w8600 <= not w8548 and not w8599;
w8601 <= w8598 and not w8599;
w8602 <= not w8600 and not w8601;
w8603 <= not w8492 and not w8602;
w8604 <= w8492 and not w8601;
w8605 <= not w8600 and w8604;
w8606 <= not w8603 and not w8605;
w8607 <= not w8491 and w8606;
w8608 <= not w8491 and not w8607;
w8609 <= w8606 and not w8607;
w8610 <= not w8608 and not w8609;
w8611 <= not w8419 and not w8421;
w8612 <= w8300 and w8377;
w8613 <= not w8300 and not w8377;
w8614 <= not w8612 and not w8613;
w8615 <= not w8336 and not w8345;
w8616 <= not w8614 and w8615;
w8617 <= w8614 and not w8615;
w8618 <= not w8616 and not w8617;
w8619 <= not w8396 and not w8414;
w8620 <= not w8618 and w8619;
w8621 <= w8618 and not w8619;
w8622 <= not w8620 and not w8621;
w8623 <= not w8361 and not w8367;
w8624 <= not w8622 and w8623;
w8625 <= w8622 and not w8623;
w8626 <= not w8624 and not w8625;
w8627 <= not w8267 and not w8284;
w8628 <= w8278 and w8357;
w8629 <= not w8278 and not w8357;
w8630 <= not w8628 and not w8629;
w8631 <= w8264 and not w8630;
w8632 <= not w8264 and w8630;
w8633 <= not w8631 and not w8632;
w8634 <= w8246 and w8410;
w8635 <= not w8246 and not w8410;
w8636 <= not w8634 and not w8635;
w8637 <= w8321 and not w8636;
w8638 <= not w8321 and w8636;
w8639 <= not w8637 and not w8638;
w8640 <= not w8633 and not w8639;
w8641 <= w8633 and w8639;
w8642 <= not w8640 and not w8641;
w8643 <= not w8627 and w8642;
w8644 <= w8627 and not w8642;
w8645 <= not w8643 and not w8644;
w8646 <= w8626 and w8645;
w8647 <= not w8626 and not w8645;
w8648 <= not w8611 and not w8647;
w8649 <= not w8646 and w8648;
w8650 <= not w8611 and not w8649;
w8651 <= not w8646 and not w8649;
w8652 <= not w8647 and w8651;
w8653 <= not w8650 and not w8652;
w8654 <= not w8230 and not w8233;
w8655 <= w8653 and w8654;
w8656 <= not w8653 and not w8654;
w8657 <= not w8655 and not w8656;
w8658 <= not w8463 and not w8467;
w8659 <= not w8224 and not w8227;
w8660 <= a(46) and a(51);
w8661 <= w491 and w8660;
w8662 <= w697 and w5366;
w8663 <= a(10) and a(51);
w8664 <= w5656 and w8663;
w8665 <= not w8662 and not w8664;
w8666 <= not w8661 and not w8665;
w8667 <= not w8661 and not w8666;
w8668 <= a(15) and a(46);
w8669 <= not w8663 and not w8668;
w8670 <= w8667 and not w8669;
w8671 <= w5656 and not w8666;
w8672 <= not w8670 and not w8671;
w8673 <= w412 and w6060;
w8674 <= a(14) and a(50);
w8675 <= w7866 and w8674;
w8676 <= w408 and w6131;
w8677 <= not w8675 and not w8676;
w8678 <= not w8673 and not w8677;
w8679 <= a(50) and not w8678;
w8680 <= a(11) and w8679;
w8681 <= not w8673 and not w8678;
w8682 <= a(12) and a(49);
w8683 <= not w7209 and not w8682;
w8684 <= w8681 and not w8683;
w8685 <= not w8680 and not w8684;
w8686 <= not w8672 and not w8685;
w8687 <= not w8672 and not w8686;
w8688 <= not w8685 and not w8686;
w8689 <= not w8687 and not w8688;
w8690 <= a(29) and a(32);
w8691 <= not w2671 and not w8690;
w8692 <= w2423 and w3618;
w8693 <= a(48) and not w8692;
w8694 <= a(13) and w8693;
w8695 <= not w8691 and w8694;
w8696 <= a(48) and not w8695;
w8697 <= a(13) and w8696;
w8698 <= not w8692 and not w8695;
w8699 <= not w8691 and w8698;
w8700 <= not w8697 and not w8699;
w8701 <= not w8689 and not w8700;
w8702 <= not w8689 and not w8701;
w8703 <= not w8700 and not w8701;
w8704 <= not w8702 and not w8703;
w8705 <= not w8215 and not w8220;
w8706 <= w8704 and w8705;
w8707 <= not w8704 and not w8705;
w8708 <= not w8706 and not w8707;
w8709 <= a(5) and a(59);
w8710 <= w7759 and w8709;
w8711 <= a(59) and a(61);
w8712 <= w2 and w8711;
w8713 <= a(5) and a(61);
w8714 <= w7229 and w8713;
w8715 <= not w8712 and not w8714;
w8716 <= not w8710 and not w8715;
w8717 <= not w8710 and not w8716;
w8718 <= a(2) and a(59);
w8719 <= a(5) and a(56);
w8720 <= not w8718 and not w8719;
w8721 <= w8717 and not w8720;
w8722 <= a(61) and not w8716;
w8723 <= a(0) and w8722;
w8724 <= not w8721 and not w8723;
w8725 <= a(20) and a(41);
w8726 <= a(21) and a(40);
w8727 <= not w8725 and not w8726;
w8728 <= w1300 and w5219;
w8729 <= a(6) and not w8728;
w8730 <= a(55) and w8729;
w8731 <= not w8727 and w8730;
w8732 <= a(55) and not w8731;
w8733 <= a(6) and w8732;
w8734 <= not w8728 and not w8731;
w8735 <= not w8727 and w8734;
w8736 <= not w8733 and not w8735;
w8737 <= not w8724 and not w8736;
w8738 <= not w8724 and not w8737;
w8739 <= not w8736 and not w8737;
w8740 <= not w8738 and not w8739;
w8741 <= w1710 and w3493;
w8742 <= a(36) and a(39);
w8743 <= w5133 and w8742;
w8744 <= w1921 and w5236;
w8745 <= not w8743 and not w8744;
w8746 <= not w8741 and not w8745;
w8747 <= a(39) and not w8746;
w8748 <= a(22) and w8747;
w8749 <= a(24) and a(37);
w8750 <= a(25) and a(36);
w8751 <= not w8749 and not w8750;
w8752 <= not w8741 and not w8746;
w8753 <= not w8751 and w8752;
w8754 <= not w8748 and not w8753;
w8755 <= not w8740 and not w8754;
w8756 <= not w8740 and not w8755;
w8757 <= not w8754 and not w8755;
w8758 <= not w8756 and not w8757;
w8759 <= not w8708 and w8758;
w8760 <= w8708 and not w8758;
w8761 <= not w8759 and not w8760;
w8762 <= not w8659 and w8761;
w8763 <= w8659 and not w8761;
w8764 <= not w8762 and not w8763;
w8765 <= not w8658 and w8764;
w8766 <= w8658 and not w8764;
w8767 <= not w8765 and not w8766;
w8768 <= w8657 and w8767;
w8769 <= not w8657 and not w8767;
w8770 <= not w8768 and not w8769;
w8771 <= not w8610 and w8770;
w8772 <= not w8609 and not w8770;
w8773 <= not w8608 and w8772;
w8774 <= not w8771 and not w8773;
w8775 <= not w8490 and w8774;
w8776 <= w8490 and not w8774;
w8777 <= not w8775 and not w8776;
w8778 <= not w8482 and not w8486;
w8779 <= not w8483 and not w8778;
w8780 <= not w8777 and w8779;
w8781 <= w8777 and not w8779;
w8782 <= not w8780 and not w8781;
w8783 <= not w8776 and not w8779;
w8784 <= not w8775 and not w8783;
w8785 <= not w8607 and not w8771;
w8786 <= not w8599 and not w8603;
w8787 <= w8514 and w8667;
w8788 <= not w8514 and not w8667;
w8789 <= not w8787 and not w8788;
w8790 <= w32 and w8242;
w8791 <= a(57) and a(59);
w8792 <= w106 and w8791;
w8793 <= a(58) and a(59);
w8794 <= w15 and w8793;
w8795 <= not w8792 and not w8794;
w8796 <= not w8790 and not w8795;
w8797 <= a(59) and not w8796;
w8798 <= a(3) and w8797;
w8799 <= not w8790 and not w8796;
w8800 <= a(4) and a(58);
w8801 <= a(5) and a(57);
w8802 <= not w8800 and not w8801;
w8803 <= w8799 and not w8802;
w8804 <= not w8798 and not w8803;
w8805 <= w8789 and not w8804;
w8806 <= w8789 and not w8805;
w8807 <= not w8804 and not w8805;
w8808 <= not w8806 and not w8807;
w8809 <= not w8520 and not w8536;
w8810 <= w8808 and w8809;
w8811 <= not w8808 and not w8809;
w8812 <= not w8810 and not w8811;
w8813 <= not w8564 and not w8568;
w8814 <= not w8812 and w8813;
w8815 <= w8812 and not w8813;
w8816 <= not w8814 and not w8815;
w8817 <= not w8613 and not w8617;
w8818 <= not w8579 and not w8582;
w8819 <= w8817 and w8818;
w8820 <= not w8817 and not w8818;
w8821 <= not w8819 and not w8820;
w8822 <= not w8629 and not w8632;
w8823 <= not w8821 and w8822;
w8824 <= w8821 and not w8822;
w8825 <= not w8823 and not w8824;
w8826 <= not w8707 and not w8760;
w8827 <= w8825 and not w8826;
w8828 <= w8825 and not w8827;
w8829 <= not w8826 and not w8827;
w8830 <= not w8828 and not w8829;
w8831 <= w8816 and not w8830;
w8832 <= not w8816 and not w8829;
w8833 <= not w8828 and w8832;
w8834 <= not w8831 and not w8833;
w8835 <= not w8786 and w8834;
w8836 <= w8786 and not w8834;
w8837 <= not w8835 and not w8836;
w8838 <= not w8591 and not w8595;
w8839 <= a(8) and a(54);
w8840 <= a(18) and a(44);
w8841 <= not w8839 and not w8840;
w8842 <= a(18) and a(54);
w8843 <= w6275 and w8842;
w8844 <= w955 and w5102;
w8845 <= a(19) and a(54);
w8846 <= w5979 and w8845;
w8847 <= not w8844 and not w8846;
w8848 <= not w8843 and not w8847;
w8849 <= not w8843 and not w8848;
w8850 <= not w8841 and w8849;
w8851 <= a(43) and not w8848;
w8852 <= a(19) and w8851;
w8853 <= not w8850 and not w8852;
w8854 <= w2140 and w3956;
w8855 <= w1847 and w2778;
w8856 <= w2137 and w3125;
w8857 <= not w8855 and not w8856;
w8858 <= not w8854 and not w8857;
w8859 <= a(35) and not w8858;
w8860 <= a(27) and w8859;
w8861 <= not w8854 and not w8858;
w8862 <= a(28) and a(34);
w8863 <= a(29) and a(33);
w8864 <= not w8862 and not w8863;
w8865 <= w8861 and not w8864;
w8866 <= not w8860 and not w8865;
w8867 <= not w8853 and not w8866;
w8868 <= not w8853 and not w8867;
w8869 <= not w8866 and not w8867;
w8870 <= not w8868 and not w8869;
w8871 <= w1472 and w4889;
w8872 <= w1921 and w3609;
w8873 <= w1725 and w3977;
w8874 <= not w8872 and not w8873;
w8875 <= not w8871 and not w8874;
w8876 <= a(40) and not w8875;
w8877 <= a(22) and w8876;
w8878 <= not w8871 and not w8875;
w8879 <= a(23) and a(39);
w8880 <= a(24) and a(38);
w8881 <= not w8879 and not w8880;
w8882 <= w8878 and not w8881;
w8883 <= not w8877 and not w8882;
w8884 <= not w8870 and not w8883;
w8885 <= not w8870 and not w8884;
w8886 <= not w8883 and not w8884;
w8887 <= not w8885 and not w8886;
w8888 <= a(0) and a(62);
w8889 <= a(2) and a(60);
w8890 <= not w8888 and not w8889;
w8891 <= a(60) and a(62);
w8892 <= w2 and w8891;
w8893 <= not w8890 and not w8892;
w8894 <= w8576 and w8893;
w8895 <= not w8892 and not w8894;
w8896 <= not w8890 and w8895;
w8897 <= w8576 and not w8894;
w8898 <= not w8896 and not w8897;
w8899 <= a(21) and a(41);
w8900 <= a(25) and a(37);
w8901 <= a(26) and a(36);
w8902 <= not w8900 and not w8901;
w8903 <= w2269 and w3493;
w8904 <= w8899 and not w8903;
w8905 <= not w8902 and w8904;
w8906 <= w8899 and not w8905;
w8907 <= not w8903 and not w8905;
w8908 <= not w8902 and w8907;
w8909 <= not w8906 and not w8908;
w8910 <= not w8898 and not w8909;
w8911 <= not w8898 and not w8910;
w8912 <= not w8909 and not w8910;
w8913 <= not w8911 and not w8912;
w8914 <= a(45) and a(52);
w8915 <= w1664 and w8914;
w8916 <= w290 and w7239;
w8917 <= a(17) and a(53);
w8918 <= w6803 and w8917;
w8919 <= not w8916 and not w8918;
w8920 <= not w8915 and not w8919;
w8921 <= a(53) and not w8920;
w8922 <= a(9) and w8921;
w8923 <= not w8915 and not w8920;
w8924 <= a(10) and a(52);
w8925 <= a(17) and a(45);
w8926 <= not w8924 and not w8925;
w8927 <= w8923 and not w8926;
w8928 <= not w8922 and not w8927;
w8929 <= not w8913 and not w8928;
w8930 <= not w8913 and not w8929;
w8931 <= not w8928 and not w8929;
w8932 <= not w8930 and not w8931;
w8933 <= a(47) and a(51);
w8934 <= w622 and w8933;
w8935 <= w1649 and w8660;
w8936 <= w697 and w5472;
w8937 <= not w8935 and not w8936;
w8938 <= not w8934 and not w8937;
w8939 <= not w8934 and not w8938;
w8940 <= a(11) and a(51);
w8941 <= a(15) and a(47);
w8942 <= not w8940 and not w8941;
w8943 <= w8939 and not w8942;
w8944 <= a(46) and not w8938;
w8945 <= a(16) and w8944;
w8946 <= not w8943 and not w8945;
w8947 <= w551 and w6062;
w8948 <= w412 and w5694;
w8949 <= w554 and w6131;
w8950 <= not w8948 and not w8949;
w8951 <= not w8947 and not w8950;
w8952 <= a(50) and not w8951;
w8953 <= a(12) and w8952;
w8954 <= a(13) and a(49);
w8955 <= a(14) and a(48);
w8956 <= not w8954 and not w8955;
w8957 <= not w8947 and not w8951;
w8958 <= not w8956 and w8957;
w8959 <= not w8953 and not w8958;
w8960 <= not w8946 and not w8959;
w8961 <= not w8946 and not w8960;
w8962 <= not w8959 and not w8960;
w8963 <= not w8961 and not w8962;
w8964 <= a(6) and a(56);
w8965 <= a(7) and a(55);
w8966 <= not w8964 and not w8965;
w8967 <= a(55) and a(56);
w8968 <= w141 and w8967;
w8969 <= a(42) and not w8968;
w8970 <= a(20) and w8969;
w8971 <= not w8966 and w8970;
w8972 <= a(42) and not w8971;
w8973 <= a(20) and w8972;
w8974 <= not w8968 and not w8971;
w8975 <= not w8966 and w8974;
w8976 <= not w8973 and not w8975;
w8977 <= not w8963 and not w8976;
w8978 <= not w8963 and not w8977;
w8979 <= not w8976 and not w8977;
w8980 <= not w8978 and not w8979;
w8981 <= not w8932 and w8980;
w8982 <= w8932 and not w8980;
w8983 <= not w8981 and not w8982;
w8984 <= not w8887 and not w8983;
w8985 <= w8887 and w8983;
w8986 <= not w8984 and not w8985;
w8987 <= not w8838 and w8986;
w8988 <= not w8838 and not w8987;
w8989 <= w8986 and not w8987;
w8990 <= not w8988 and not w8989;
w8991 <= not w8651 and not w8990;
w8992 <= not w8651 and not w8991;
w8993 <= not w8990 and not w8991;
w8994 <= not w8992 and not w8993;
w8995 <= not w8837 and w8994;
w8996 <= w8837 and not w8994;
w8997 <= not w8995 and not w8996;
w8998 <= not w8656 and not w8768;
w8999 <= not w8635 and not w8638;
w9000 <= not w8737 and not w8755;
w9001 <= w8999 and w9000;
w9002 <= not w8999 and not w9000;
w9003 <= not w9001 and not w9002;
w9004 <= not w8686 and not w8701;
w9005 <= not w9003 and w9004;
w9006 <= w9003 and not w9004;
w9007 <= not w9005 and not w9006;
w9008 <= w8717 and w8734;
w9009 <= not w8717 and not w8734;
w9010 <= not w9008 and not w9009;
w9011 <= w8501 and not w9010;
w9012 <= not w8501 and w9010;
w9013 <= not w9011 and not w9012;
w9014 <= w8531 and w8561;
w9015 <= not w8531 and not w8561;
w9016 <= not w9014 and not w9015;
w9017 <= w8752 and not w9016;
w9018 <= not w8752 and w9016;
w9019 <= not w9017 and not w9018;
w9020 <= a(1) and a(61);
w9021 <= w2294 and w9020;
w9022 <= not w2294 and not w9020;
w9023 <= not w9021 and not w9022;
w9024 <= w8698 and not w9023;
w9025 <= not w8698 and w9023;
w9026 <= not w9024 and not w9025;
w9027 <= not w8681 and w9026;
w9028 <= w8681 and not w9026;
w9029 <= not w9027 and not w9028;
w9030 <= w9019 and w9029;
w9031 <= w9019 and not w9030;
w9032 <= w9029 and not w9030;
w9033 <= not w9031 and not w9032;
w9034 <= w9013 and not w9033;
w9035 <= w9013 and not w9034;
w9036 <= not w9033 and not w9034;
w9037 <= not w9035 and not w9036;
w9038 <= w9007 and not w9037;
w9039 <= w9007 and not w9038;
w9040 <= not w9037 and not w9038;
w9041 <= not w9039 and not w9040;
w9042 <= not w8541 and not w8545;
w9043 <= w9041 and w9042;
w9044 <= not w9041 and not w9042;
w9045 <= not w9043 and not w9044;
w9046 <= not w8641 and not w8643;
w9047 <= not w8585 and not w8588;
w9048 <= w9046 and w9047;
w9049 <= not w9046 and not w9047;
w9050 <= not w9048 and not w9049;
w9051 <= not w8621 and not w8625;
w9052 <= not w9050 and w9051;
w9053 <= w9050 and not w9051;
w9054 <= not w9052 and not w9053;
w9055 <= not w8762 and not w8765;
w9056 <= not w9054 and w9055;
w9057 <= w9054 and not w9055;
w9058 <= not w9056 and not w9057;
w9059 <= w9045 and w9058;
w9060 <= not w9045 and not w9058;
w9061 <= not w9059 and not w9060;
w9062 <= not w8998 and w9061;
w9063 <= not w8998 and not w9062;
w9064 <= w9061 and not w9062;
w9065 <= not w9063 and not w9064;
w9066 <= w8997 and not w9065;
w9067 <= not w8997 and not w9064;
w9068 <= not w9063 and w9067;
w9069 <= not w9066 and not w9068;
w9070 <= not w8785 and w9069;
w9071 <= w8785 and not w9069;
w9072 <= not w9070 and not w9071;
w9073 <= w8784 and not w9072;
w9074 <= not w8784 and not w9071;
w9075 <= not w9070 and w9074;
w9076 <= not w9073 and not w9075;
w9077 <= not w9070 and not w9074;
w9078 <= not w9062 and not w9066;
w9079 <= not w8987 and not w8991;
w9080 <= not w9030 and not w9034;
w9081 <= not w9002 and not w9006;
w9082 <= w9080 and w9081;
w9083 <= not w9080 and not w9081;
w9084 <= not w9082 and not w9083;
w9085 <= not w8811 and not w8815;
w9086 <= not w9084 and w9085;
w9087 <= w9084 and not w9085;
w9088 <= not w9086 and not w9087;
w9089 <= not w8788 and not w8805;
w9090 <= not w9015 and not w9018;
w9091 <= w9089 and w9090;
w9092 <= not w9089 and not w9090;
w9093 <= not w9091 and not w9092;
w9094 <= not w9025 and not w9027;
w9095 <= not w9093 and w9094;
w9096 <= w9093 and not w9094;
w9097 <= not w9095 and not w9096;
w9098 <= not w8932 and not w8980;
w9099 <= not w8984 and not w9098;
w9100 <= w9097 and not w9099;
w9101 <= not w9097 and w9099;
w9102 <= not w9100 and not w9101;
w9103 <= w8878 and w8974;
w9104 <= not w8878 and not w8974;
w9105 <= not w9103 and not w9104;
w9106 <= w8957 and not w9105;
w9107 <= not w8957 and w9105;
w9108 <= not w9106 and not w9107;
w9109 <= w8799 and w8907;
w9110 <= not w8799 and not w8907;
w9111 <= not w9109 and not w9110;
w9112 <= w8895 and not w9111;
w9113 <= not w8895 and w9111;
w9114 <= not w9112 and not w9113;
w9115 <= not w9009 and not w9012;
w9116 <= not w9114 and w9115;
w9117 <= w9114 and not w9115;
w9118 <= not w9116 and not w9117;
w9119 <= w9108 and w9118;
w9120 <= not w9108 and not w9118;
w9121 <= not w9119 and not w9120;
w9122 <= w9102 and w9121;
w9123 <= not w9102 and not w9121;
w9124 <= not w9122 and not w9123;
w9125 <= w9088 and w9124;
w9126 <= not w9088 and not w9124;
w9127 <= not w9079 and not w9126;
w9128 <= not w9125 and w9127;
w9129 <= not w9079 and not w9128;
w9130 <= not w9125 and not w9128;
w9131 <= not w9126 and w9130;
w9132 <= not w9129 and not w9131;
w9133 <= not w8835 and not w8996;
w9134 <= w9132 and w9133;
w9135 <= not w9132 and not w9133;
w9136 <= not w9134 and not w9135;
w9137 <= not w9057 and not w9059;
w9138 <= not w9049 and not w9053;
w9139 <= w8861 and w8923;
w9140 <= not w8861 and not w8923;
w9141 <= not w9139 and not w9140;
w9142 <= w8849 and not w9141;
w9143 <= not w8849 and w9141;
w9144 <= not w9142 and not w9143;
w9145 <= not w8867 and not w8884;
w9146 <= not w9144 and w9145;
w9147 <= w9144 and not w9145;
w9148 <= not w9146 and not w9147;
w9149 <= not w8960 and not w8977;
w9150 <= not w9148 and w9149;
w9151 <= w9148 and not w9149;
w9152 <= not w9150 and not w9151;
w9153 <= not w8820 and not w8824;
w9154 <= not w8910 and not w8929;
w9155 <= w9153 and w9154;
w9156 <= not w9153 and not w9154;
w9157 <= not w9155 and not w9156;
w9158 <= a(0) and a(63);
w9159 <= w9021 and w9158;
w9160 <= w9021 and not w9159;
w9161 <= not w9021 and w9158;
w9162 <= not w9160 and not w9161;
w9163 <= a(62) and w2493;
w9164 <= a(32) and not w9163;
w9165 <= a(1) and not w9163;
w9166 <= a(62) and w9165;
w9167 <= not w9164 and not w9166;
w9168 <= not w9162 and not w9167;
w9169 <= not w9162 and not w9168;
w9170 <= not w9167 and not w9168;
w9171 <= not w9169 and not w9170;
w9172 <= w2269 and w4371;
w9173 <= w2107 and w5236;
w9174 <= w1710 and w4889;
w9175 <= not w9173 and not w9174;
w9176 <= not w9172 and not w9175;
w9177 <= not w9172 and not w9176;
w9178 <= a(25) and a(38);
w9179 <= a(26) and a(37);
w9180 <= not w9178 and not w9179;
w9181 <= w9177 and not w9180;
w9182 <= a(39) and not w9176;
w9183 <= a(24) and w9182;
w9184 <= not w9181 and not w9183;
w9185 <= w2140 and w3125;
w9186 <= w1847 and w4401;
w9187 <= w2137 and w3634;
w9188 <= not w9186 and not w9187;
w9189 <= not w9185 and not w9188;
w9190 <= a(36) and not w9189;
w9191 <= a(27) and w9190;
w9192 <= a(28) and a(35);
w9193 <= a(29) and a(34);
w9194 <= not w9192 and not w9193;
w9195 <= not w9185 and not w9189;
w9196 <= not w9194 and w9195;
w9197 <= not w9191 and not w9196;
w9198 <= not w9184 and not w9197;
w9199 <= not w9184 and not w9198;
w9200 <= not w9197 and not w9198;
w9201 <= not w9199 and not w9200;
w9202 <= not w9171 and w9201;
w9203 <= w9171 and not w9201;
w9204 <= not w9202 and not w9203;
w9205 <= w9157 and not w9204;
w9206 <= w9157 and not w9205;
w9207 <= not w9204 and not w9205;
w9208 <= not w9206 and not w9207;
w9209 <= not w9152 and w9208;
w9210 <= w9152 and not w9208;
w9211 <= not w9209 and not w9210;
w9212 <= not w9138 and w9211;
w9213 <= w9138 and not w9211;
w9214 <= not w9212 and not w9213;
w9215 <= not w9137 and w9214;
w9216 <= w9137 and not w9214;
w9217 <= not w9215 and not w9216;
w9218 <= not w9038 and not w9044;
w9219 <= not w8827 and not w8831;
w9220 <= a(46) and a(54);
w9221 <= w1482 and w9220;
w9222 <= w6803 and w8842;
w9223 <= w858 and w5366;
w9224 <= not w9222 and not w9223;
w9225 <= not w9221 and not w9224;
w9226 <= not w9221 and not w9225;
w9227 <= a(9) and a(54);
w9228 <= a(17) and a(46);
w9229 <= not w9227 and not w9228;
w9230 <= w9226 and not w9229;
w9231 <= a(45) and not w9225;
w9232 <= a(18) and w9231;
w9233 <= not w9230 and not w9232;
w9234 <= a(47) and a(52);
w9235 <= w1649 and w9234;
w9236 <= w529 and w7239;
w9237 <= a(16) and a(53);
w9238 <= w7536 and w9237;
w9239 <= not w9236 and not w9238;
w9240 <= not w9235 and not w9239;
w9241 <= a(53) and not w9240;
w9242 <= a(10) and w9241;
w9243 <= a(11) and a(52);
w9244 <= a(16) and a(47);
w9245 <= not w9243 and not w9244;
w9246 <= not w9235 and not w9240;
w9247 <= not w9245 and w9246;
w9248 <= not w9242 and not w9247;
w9249 <= not w9233 and not w9248;
w9250 <= not w9233 and not w9249;
w9251 <= not w9248 and not w9249;
w9252 <= not w9250 and not w9251;
w9253 <= w554 and w6370;
w9254 <= w627 and w5694;
w9255 <= a(12) and a(51);
w9256 <= w7157 and w9255;
w9257 <= not w9254 and not w9256;
w9258 <= not w9253 and not w9257;
w9259 <= w7157 and not w9258;
w9260 <= not w9253 and not w9258;
w9261 <= a(13) and a(50);
w9262 <= not w9255 and not w9261;
w9263 <= w9260 and not w9262;
w9264 <= not w9259 and not w9263;
w9265 <= not w9252 and not w9264;
w9266 <= not w9252 and not w9265;
w9267 <= not w9264 and not w9265;
w9268 <= not w9266 and not w9267;
w9269 <= a(6) and a(57);
w9270 <= a(20) and a(43);
w9271 <= not w9269 and not w9270;
w9272 <= w9269 and w9270;
w9273 <= a(40) and not w9272;
w9274 <= a(23) and w9273;
w9275 <= not w9271 and w9274;
w9276 <= not w9272 and not w9275;
w9277 <= not w9271 and w9276;
w9278 <= a(40) and not w9275;
w9279 <= a(23) and w9278;
w9280 <= not w9277 and not w9279;
w9281 <= a(30) and a(33);
w9282 <= not w3618 and not w9281;
w9283 <= w3618 and w9281;
w9284 <= a(49) and not w9283;
w9285 <= a(14) and w9284;
w9286 <= not w9282 and w9285;
w9287 <= a(49) and not w9286;
w9288 <= a(14) and w9287;
w9289 <= not w9283 and not w9286;
w9290 <= not w9282 and w9289;
w9291 <= not w9288 and not w9290;
w9292 <= not w9280 and not w9291;
w9293 <= not w9280 and not w9292;
w9294 <= not w9291 and not w9292;
w9295 <= not w9293 and not w9294;
w9296 <= a(44) and a(55);
w9297 <= w1662 and w9296;
w9298 <= w186 and w8967;
w9299 <= a(44) and a(56);
w9300 <= w1468 and w9299;
w9301 <= not w9298 and not w9300;
w9302 <= not w9297 and not w9301;
w9303 <= a(56) and not w9302;
w9304 <= a(7) and w9303;
w9305 <= a(8) and a(55);
w9306 <= a(19) and a(44);
w9307 <= not w9305 and not w9306;
w9308 <= not w9297 and not w9302;
w9309 <= not w9307 and w9308;
w9310 <= not w9304 and not w9309;
w9311 <= not w9295 and not w9310;
w9312 <= not w9295 and not w9311;
w9313 <= not w9310 and not w9311;
w9314 <= not w9312 and not w9313;
w9315 <= a(59) and a(60);
w9316 <= w15 and w9315;
w9317 <= w58 and w8711;
w9318 <= a(60) and a(61);
w9319 <= w24 and w9318;
w9320 <= not w9317 and not w9319;
w9321 <= not w9316 and not w9320;
w9322 <= a(2) and not w9321;
w9323 <= a(61) and w9322;
w9324 <= not w9316 and not w9321;
w9325 <= a(3) and a(60);
w9326 <= a(4) and a(59);
w9327 <= not w9325 and not w9326;
w9328 <= w9324 and not w9327;
w9329 <= not w9323 and not w9328;
w9330 <= w8939 and not w9329;
w9331 <= not w8939 and w9329;
w9332 <= not w9330 and not w9331;
w9333 <= a(21) and a(42);
w9334 <= a(22) and a(41);
w9335 <= not w9333 and not w9334;
w9336 <= w1380 and w5150;
w9337 <= a(5) and not w9336;
w9338 <= a(58) and w9337;
w9339 <= not w9335 and w9338;
w9340 <= a(58) and not w9339;
w9341 <= a(5) and w9340;
w9342 <= not w9336 and not w9339;
w9343 <= not w9335 and w9342;
w9344 <= not w9341 and not w9343;
w9345 <= not w9332 and not w9344;
w9346 <= w9332 and w9344;
w9347 <= not w9345 and not w9346;
w9348 <= w9314 and w9347;
w9349 <= not w9314 and not w9347;
w9350 <= not w9348 and not w9349;
w9351 <= not w9268 and not w9350;
w9352 <= w9268 and w9350;
w9353 <= not w9351 and not w9352;
w9354 <= not w9219 and w9353;
w9355 <= not w9219 and not w9354;
w9356 <= w9353 and not w9354;
w9357 <= not w9355 and not w9356;
w9358 <= not w9218 and not w9357;
w9359 <= not w9218 and not w9358;
w9360 <= not w9357 and not w9358;
w9361 <= not w9359 and not w9360;
w9362 <= w9217 and not w9361;
w9363 <= w9217 and not w9362;
w9364 <= not w9361 and not w9362;
w9365 <= not w9363 and not w9364;
w9366 <= not w9136 and w9365;
w9367 <= w9136 and not w9365;
w9368 <= not w9366 and not w9367;
w9369 <= w9078 and not w9368;
w9370 <= not w9078 and w9368;
w9371 <= not w9369 and not w9370;
w9372 <= not w9077 and not w9371;
w9373 <= w9077 and w9371;
w9374 <= not w9372 and not w9373;
w9375 <= not w9077 and not w9369;
w9376 <= not w9370 and not w9375;
w9377 <= not w9215 and not w9362;
w9378 <= not w9354 and not w9358;
w9379 <= not w9210 and not w9212;
w9380 <= not w9314 and w9347;
w9381 <= not w9351 and not w9380;
w9382 <= not w9156 and not w9205;
w9383 <= w9381 and w9382;
w9384 <= not w9381 and not w9382;
w9385 <= not w9383 and not w9384;
w9386 <= not w9171 and not w9201;
w9387 <= not w9198 and not w9386;
w9388 <= w9226 and w9276;
w9389 <= not w9226 and not w9276;
w9390 <= not w9388 and not w9389;
w9391 <= w9195 and not w9390;
w9392 <= not w9195 and w9390;
w9393 <= not w9391 and not w9392;
w9394 <= w9324 and w9342;
w9395 <= not w9324 and not w9342;
w9396 <= not w9394 and not w9395;
w9397 <= w9308 and not w9396;
w9398 <= not w9308 and w9396;
w9399 <= not w9397 and not w9398;
w9400 <= not w9393 and not w9399;
w9401 <= w9393 and w9399;
w9402 <= not w9400 and not w9401;
w9403 <= not w9387 and w9402;
w9404 <= w9387 and not w9402;
w9405 <= not w9403 and not w9404;
w9406 <= not w9385 and not w9405;
w9407 <= w9385 and w9405;
w9408 <= not w9406 and not w9407;
w9409 <= not w9379 and w9408;
w9410 <= not w9379 and not w9409;
w9411 <= w9408 and not w9409;
w9412 <= not w9410 and not w9411;
w9413 <= not w9378 and not w9412;
w9414 <= not w9378 and not w9413;
w9415 <= not w9412 and not w9413;
w9416 <= not w9414 and not w9415;
w9417 <= not w9377 and not w9416;
w9418 <= not w9377 and not w9417;
w9419 <= not w9416 and not w9417;
w9420 <= not w9418 and not w9419;
w9421 <= not w9100 and not w9122;
w9422 <= a(7) and a(57);
w9423 <= not w5705 and not w9422;
w9424 <= a(17) and a(57);
w9425 <= w6786 and w9424;
w9426 <= a(58) and w6416;
w9427 <= a(17) and w9426;
w9428 <= w141 and w8242;
w9429 <= not w9427 and not w9428;
w9430 <= not w9425 and not w9429;
w9431 <= not w9425 and not w9430;
w9432 <= not w9423 and w9431;
w9433 <= a(58) and not w9430;
w9434 <= a(6) and w9433;
w9435 <= not w9432 and not w9434;
w9436 <= w1380 and w4824;
w9437 <= w1499 and w4445;
w9438 <= w1300 and w5102;
w9439 <= not w9437 and not w9438;
w9440 <= not w9436 and not w9439;
w9441 <= a(44) and not w9440;
w9442 <= a(20) and w9441;
w9443 <= not w9436 and not w9440;
w9444 <= a(21) and a(43);
w9445 <= a(22) and a(42);
w9446 <= not w9444 and not w9445;
w9447 <= w9443 and not w9446;
w9448 <= not w9442 and not w9447;
w9449 <= not w9435 and not w9448;
w9450 <= not w9435 and not w9449;
w9451 <= not w9448 and not w9449;
w9452 <= not w9450 and not w9451;
w9453 <= w1710 and w3977;
w9454 <= w1353 and w3790;
w9455 <= w1472 and w5219;
w9456 <= not w9454 and not w9455;
w9457 <= not w9453 and not w9456;
w9458 <= a(41) and not w9457;
w9459 <= a(23) and w9458;
w9460 <= not w9453 and not w9457;
w9461 <= a(24) and a(40);
w9462 <= a(25) and a(39);
w9463 <= not w9461 and not w9462;
w9464 <= w9460 and not w9463;
w9465 <= not w9459 and not w9464;
w9466 <= not w9452 and not w9465;
w9467 <= not w9452 and not w9466;
w9468 <= not w9465 and not w9466;
w9469 <= not w9467 and not w9468;
w9470 <= a(8) and a(56);
w9471 <= not w6448 and not w9470;
w9472 <= a(48) and a(56);
w9473 <= w1315 and w9472;
w9474 <= a(38) and not w9473;
w9475 <= a(26) and w9474;
w9476 <= not w9471 and w9475;
w9477 <= not w9473 and not w9476;
w9478 <= not w9471 and w9477;
w9479 <= a(38) and not w9476;
w9480 <= a(26) and w9479;
w9481 <= not w9478 and not w9480;
w9482 <= w2140 and w3634;
w9483 <= w1847 and w4837;
w9484 <= w2137 and w3493;
w9485 <= not w9483 and not w9484;
w9486 <= not w9482 and not w9485;
w9487 <= w3865 and not w9486;
w9488 <= not w9482 and not w9486;
w9489 <= a(28) and a(36);
w9490 <= a(29) and a(35);
w9491 <= not w9489 and not w9490;
w9492 <= w9488 and not w9491;
w9493 <= not w9487 and not w9492;
w9494 <= not w9481 and not w9493;
w9495 <= not w9481 and not w9494;
w9496 <= not w9493 and not w9494;
w9497 <= not w9495 and not w9496;
w9498 <= a(30) and a(34);
w9499 <= not w2404 and not w9498;
w9500 <= w2671 and w3956;
w9501 <= w8674 and not w9500;
w9502 <= not w9499 and w9501;
w9503 <= w8674 and not w9502;
w9504 <= not w9500 and not w9502;
w9505 <= not w9499 and w9504;
w9506 <= not w9503 and not w9505;
w9507 <= not w9497 and not w9506;
w9508 <= not w9497 and not w9507;
w9509 <= not w9506 and not w9507;
w9510 <= not w9508 and not w9509;
w9511 <= w955 and w5366;
w9512 <= a(18) and a(46);
w9513 <= a(19) and a(45);
w9514 <= not w9512 and not w9513;
w9515 <= not w9511 and not w9514;
w9516 <= w8709 and w9515;
w9517 <= w8709 and not w9516;
w9518 <= not w9511 and not w9516;
w9519 <= not w9514 and w9518;
w9520 <= not w9517 and not w9519;
w9521 <= not w9159 and not w9168;
w9522 <= not w9520 and w9521;
w9523 <= w9520 and not w9521;
w9524 <= not w9522 and not w9523;
w9525 <= w15 and w9318;
w9526 <= w58 and w8891;
w9527 <= a(61) and a(62);
w9528 <= w24 and w9527;
w9529 <= not w9526 and not w9528;
w9530 <= not w9525 and not w9529;
w9531 <= a(62) and not w9530;
w9532 <= a(2) and w9531;
w9533 <= not w9525 and not w9530;
w9534 <= a(3) and a(61);
w9535 <= a(4) and a(60);
w9536 <= not w9534 and not w9535;
w9537 <= w9533 and not w9536;
w9538 <= not w9532 and not w9537;
w9539 <= not w9524 and not w9538;
w9540 <= w9524 and w9538;
w9541 <= not w9539 and not w9540;
w9542 <= w9510 and w9541;
w9543 <= not w9510 and not w9541;
w9544 <= not w9542 and not w9543;
w9545 <= not w9469 and not w9544;
w9546 <= w9469 and w9544;
w9547 <= not w9545 and not w9546;
w9548 <= not w9421 and w9547;
w9549 <= w9421 and not w9547;
w9550 <= not w9548 and not w9549;
w9551 <= not w9104 and not w9107;
w9552 <= not w9140 and not w9143;
w9553 <= w9551 and w9552;
w9554 <= not w9551 and not w9552;
w9555 <= not w9553 and not w9554;
w9556 <= not w9110 and not w9113;
w9557 <= not w9555 and w9556;
w9558 <= w9555 and not w9556;
w9559 <= not w9557 and not w9558;
w9560 <= not w9147 and not w9151;
w9561 <= not w9117 and not w9119;
w9562 <= not w9560 and not w9561;
w9563 <= not w9560 and not w9562;
w9564 <= not w9561 and not w9562;
w9565 <= not w9563 and not w9564;
w9566 <= w9559 and not w9565;
w9567 <= not w9559 and w9565;
w9568 <= w9550 and not w9567;
w9569 <= not w9566 and w9568;
w9570 <= w9550 and not w9569;
w9571 <= not w9567 and not w9569;
w9572 <= not w9566 and w9571;
w9573 <= not w9570 and not w9572;
w9574 <= w9177 and w9260;
w9575 <= not w9177 and not w9260;
w9576 <= not w9574 and not w9575;
w9577 <= w9246 and not w9576;
w9578 <= not w9246 and w9576;
w9579 <= not w9577 and not w9578;
w9580 <= not w9292 and not w9311;
w9581 <= not w9579 and w9580;
w9582 <= w9579 and not w9580;
w9583 <= not w9581 and not w9582;
w9584 <= not w9249 and not w9265;
w9585 <= not w9583 and w9584;
w9586 <= w9583 and not w9584;
w9587 <= not w9585 and not w9586;
w9588 <= not w9083 and not w9087;
w9589 <= not w9587 and w9588;
w9590 <= w9587 and not w9588;
w9591 <= not w9589 and not w9590;
w9592 <= not w9092 and not w9096;
w9593 <= not w8939 and not w9329;
w9594 <= not w9345 and not w9593;
w9595 <= w9592 and w9594;
w9596 <= not w9592 and not w9594;
w9597 <= not w9595 and not w9596;
w9598 <= a(62) and a(63);
w9599 <= w2493 and w9598;
w9600 <= w9163 and not w9599;
w9601 <= a(63) and w9165;
w9602 <= not w9600 and not w9601;
w9603 <= not w9289 and not w9602;
w9604 <= not w9289 and not w9603;
w9605 <= not w9602 and not w9603;
w9606 <= not w9604 and not w9605;
w9607 <= a(49) and a(55);
w9608 <= w1323 and w9607;
w9609 <= w290 and w7507;
w9610 <= not w9608 and not w9609;
w9611 <= a(10) and a(54);
w9612 <= a(15) and a(49);
w9613 <= w9611 and w9612;
w9614 <= not w9610 and not w9613;
w9615 <= not w9613 and not w9614;
w9616 <= not w9611 and not w9612;
w9617 <= w9615 and not w9616;
w9618 <= a(55) and not w9614;
w9619 <= a(9) and w9618;
w9620 <= not w9617 and not w9619;
w9621 <= w408 and w7239;
w9622 <= w624 and w7038;
w9623 <= w554 and w6774;
w9624 <= not w9622 and not w9623;
w9625 <= not w9621 and not w9624;
w9626 <= a(51) and not w9625;
w9627 <= a(13) and w9626;
w9628 <= a(11) and a(53);
w9629 <= a(12) and a(52);
w9630 <= not w9628 and not w9629;
w9631 <= not w9621 and not w9625;
w9632 <= not w9630 and w9631;
w9633 <= not w9627 and not w9632;
w9634 <= not w9620 and not w9633;
w9635 <= not w9620 and not w9634;
w9636 <= not w9633 and not w9634;
w9637 <= not w9635 and not w9636;
w9638 <= not w9606 and w9637;
w9639 <= w9606 and not w9637;
w9640 <= not w9638 and not w9639;
w9641 <= w9597 and not w9640;
w9642 <= w9597 and not w9641;
w9643 <= not w9640 and not w9641;
w9644 <= not w9642 and not w9643;
w9645 <= not w9591 and w9644;
w9646 <= w9591 and not w9644;
w9647 <= not w9645 and not w9646;
w9648 <= not w9130 and w9647;
w9649 <= w9130 and not w9647;
w9650 <= not w9648 and not w9649;
w9651 <= not w9573 and w9650;
w9652 <= w9573 and not w9650;
w9653 <= not w9651 and not w9652;
w9654 <= not w9420 and w9653;
w9655 <= w9420 and not w9653;
w9656 <= not w9654 and not w9655;
w9657 <= not w9135 and not w9367;
w9658 <= not w9656 and w9657;
w9659 <= w9656 and not w9657;
w9660 <= not w9658 and not w9659;
w9661 <= w9376 and not w9660;
w9662 <= not w9376 and not w9658;
w9663 <= not w9659 and w9662;
w9664 <= not w9661 and not w9663;
w9665 <= not w9659 and not w9662;
w9666 <= not w9417 and not w9654;
w9667 <= not w9648 and not w9651;
w9668 <= not w9548 and not w9569;
w9669 <= not w9590 and not w9646;
w9670 <= not w9510 and w9541;
w9671 <= not w9545 and not w9670;
w9672 <= not w9596 and not w9641;
w9673 <= w9671 and w9672;
w9674 <= not w9671 and not w9672;
w9675 <= not w9673 and not w9674;
w9676 <= not w9606 and not w9637;
w9677 <= not w9634 and not w9676;
w9678 <= w9460 and w9615;
w9679 <= not w9460 and not w9615;
w9680 <= not w9678 and not w9679;
w9681 <= w9431 and not w9680;
w9682 <= not w9431 and w9680;
w9683 <= not w9681 and not w9682;
w9684 <= w9518 and w9533;
w9685 <= not w9518 and not w9533;
w9686 <= not w9684 and not w9685;
w9687 <= w9477 and not w9686;
w9688 <= not w9477 and w9686;
w9689 <= not w9687 and not w9688;
w9690 <= not w9683 and not w9689;
w9691 <= w9683 and w9689;
w9692 <= not w9690 and not w9691;
w9693 <= not w9677 and w9692;
w9694 <= w9677 and not w9692;
w9695 <= not w9693 and not w9694;
w9696 <= not w9675 and not w9695;
w9697 <= w9675 and w9695;
w9698 <= not w9696 and not w9697;
w9699 <= not w9669 and w9698;
w9700 <= w9669 and not w9698;
w9701 <= not w9699 and not w9700;
w9702 <= not w9668 and w9701;
w9703 <= w9668 and not w9701;
w9704 <= not w9702 and not w9703;
w9705 <= w9667 and not w9704;
w9706 <= not w9667 and w9704;
w9707 <= not w9705 and not w9706;
w9708 <= not w9409 and not w9413;
w9709 <= not w9554 and not w9558;
w9710 <= not w9520 and not w9521;
w9711 <= not w9539 and not w9710;
w9712 <= w9709 and w9711;
w9713 <= not w9709 and not w9711;
w9714 <= not w9712 and not w9713;
w9715 <= a(61) and a(63);
w9716 <= w58 and w9715;
w9717 <= a(61) and not w9716;
w9718 <= a(4) and w9717;
w9719 <= a(2) and not w9716;
w9720 <= a(63) and w9719;
w9721 <= not w9718 and not w9720;
w9722 <= not w9504 and not w9721;
w9723 <= not w9504 and not w9722;
w9724 <= not w9721 and not w9722;
w9725 <= not w9723 and not w9724;
w9726 <= w554 and w7239;
w9727 <= w7966 and w8370;
w9728 <= not w9726 and not w9727;
w9729 <= a(13) and a(52);
w9730 <= a(18) and a(47);
w9731 <= w9729 and w9730;
w9732 <= not w9728 and not w9731;
w9733 <= not w9731 and not w9732;
w9734 <= not w9729 and not w9730;
w9735 <= w9733 and not w9734;
w9736 <= a(53) and not w9732;
w9737 <= a(12) and w9736;
w9738 <= not w9735 and not w9737;
w9739 <= w701 and w6370;
w9740 <= a(49) and a(51);
w9741 <= w699 and w9740;
w9742 <= w697 and w6131;
w9743 <= not w9741 and not w9742;
w9744 <= not w9739 and not w9743;
w9745 <= w7445 and not w9744;
w9746 <= a(14) and a(51);
w9747 <= a(15) and a(50);
w9748 <= not w9746 and not w9747;
w9749 <= not w9739 and not w9744;
w9750 <= not w9748 and w9749;
w9751 <= not w9745 and not w9750;
w9752 <= not w9738 and not w9751;
w9753 <= not w9738 and not w9752;
w9754 <= not w9751 and not w9752;
w9755 <= not w9753 and not w9754;
w9756 <= not w9725 and w9755;
w9757 <= w9725 and not w9755;
w9758 <= not w9756 and not w9757;
w9759 <= w9714 and not w9758;
w9760 <= w9714 and not w9759;
w9761 <= not w9758 and not w9759;
w9762 <= not w9760 and not w9761;
w9763 <= w9443 and w9488;
w9764 <= not w9443 and not w9488;
w9765 <= not w9763 and not w9764;
w9766 <= w9631 and not w9765;
w9767 <= not w9631 and w9765;
w9768 <= not w9766 and not w9767;
w9769 <= not w9494 and not w9507;
w9770 <= not w9768 and w9769;
w9771 <= w9768 and not w9769;
w9772 <= not w9770 and not w9771;
w9773 <= not w9449 and not w9466;
w9774 <= not w9772 and w9773;
w9775 <= w9772 and not w9773;
w9776 <= not w9774 and not w9775;
w9777 <= not w9562 and not w9566;
w9778 <= w9776 and not w9777;
w9779 <= w9776 and not w9778;
w9780 <= not w9777 and not w9778;
w9781 <= not w9779 and not w9780;
w9782 <= not w9762 and not w9781;
w9783 <= not w9762 and not w9782;
w9784 <= not w9781 and not w9782;
w9785 <= not w9783 and not w9784;
w9786 <= not w9708 and not w9785;
w9787 <= not w9708 and not w9786;
w9788 <= not w9785 and not w9786;
w9789 <= not w9787 and not w9788;
w9790 <= not w9384 and not w9407;
w9791 <= a(20) and a(56);
w9792 <= w6803 and w9791;
w9793 <= w290 and w8967;
w9794 <= not w9792 and not w9793;
w9795 <= a(10) and a(55);
w9796 <= a(20) and a(45);
w9797 <= w9795 and w9796;
w9798 <= not w9794 and not w9797;
w9799 <= not w9797 and not w9798;
w9800 <= not w9795 and not w9796;
w9801 <= w9799 and not w9800;
w9802 <= a(56) and not w9798;
w9803 <= a(9) and w9802;
w9804 <= not w9801 and not w9803;
w9805 <= w1710 and w5219;
w9806 <= w1353 and w6259;
w9807 <= w1472 and w5150;
w9808 <= not w9806 and not w9807;
w9809 <= not w9805 and not w9808;
w9810 <= a(42) and not w9809;
w9811 <= a(23) and w9810;
w9812 <= a(24) and a(41);
w9813 <= a(25) and a(40);
w9814 <= not w9812 and not w9813;
w9815 <= not w9805 and not w9809;
w9816 <= not w9814 and w9815;
w9817 <= not w9811 and not w9816;
w9818 <= not w9804 and not w9817;
w9819 <= not w9804 and not w9818;
w9820 <= not w9817 and not w9818;
w9821 <= not w9819 and not w9820;
w9822 <= w2137 and w4371;
w9823 <= w2606 and w5236;
w9824 <= w2033 and w4889;
w9825 <= not w9823 and not w9824;
w9826 <= not w9822 and not w9825;
w9827 <= a(39) and not w9826;
w9828 <= a(26) and w9827;
w9829 <= not w9822 and not w9826;
w9830 <= a(27) and a(38);
w9831 <= a(28) and a(37);
w9832 <= not w9830 and not w9831;
w9833 <= w9829 and not w9832;
w9834 <= not w9828 and not w9833;
w9835 <= not w9821 and not w9834;
w9836 <= not w9821 and not w9835;
w9837 <= not w9834 and not w9835;
w9838 <= not w9836 and not w9837;
w9839 <= a(11) and a(54);
w9840 <= a(19) and a(46);
w9841 <= not w9839 and not w9840;
w9842 <= w9839 and w9840;
w9843 <= a(29) and not w9842;
w9844 <= a(36) and w9843;
w9845 <= not w9841 and w9844;
w9846 <= not w9842 and not w9845;
w9847 <= not w9841 and w9846;
w9848 <= a(36) and not w9845;
w9849 <= a(29) and w9848;
w9850 <= not w9847 and not w9849;
w9851 <= w3618 and w3956;
w9852 <= w2949 and w3830;
w9853 <= w2671 and w3125;
w9854 <= not w9852 and not w9853;
w9855 <= not w9851 and not w9854;
w9856 <= w3830 and not w9855;
w9857 <= not w9851 and not w9855;
w9858 <= not w2949 and not w6291;
w9859 <= w9857 and not w9858;
w9860 <= not w9856 and not w9859;
w9861 <= not w9850 and not w9860;
w9862 <= not w9850 and not w9861;
w9863 <= not w9860 and not w9861;
w9864 <= not w9862 and not w9863;
w9865 <= a(3) and a(62);
w9866 <= not a(33) and not w9865;
w9867 <= a(33) and w9865;
w9868 <= w6750 and not w9867;
w9869 <= not w9866 and w9868;
w9870 <= w6750 and not w9869;
w9871 <= not w9867 and not w9869;
w9872 <= not w9866 and w9871;
w9873 <= not w9870 and not w9872;
w9874 <= not w9864 and not w9873;
w9875 <= not w9864 and not w9874;
w9876 <= not w9873 and not w9874;
w9877 <= not w9875 and not w9876;
w9878 <= a(21) and a(44);
w9879 <= a(22) and a(43);
w9880 <= not w9878 and not w9879;
w9881 <= w1380 and w5102;
w9882 <= a(8) and not w9881;
w9883 <= a(57) and w9882;
w9884 <= not w9880 and w9883;
w9885 <= a(8) and not w9884;
w9886 <= a(57) and w9885;
w9887 <= not w9881 and not w9884;
w9888 <= not w9880 and w9887;
w9889 <= not w9886 and not w9888;
w9890 <= not w9599 and not w9603;
w9891 <= not w9889 and w9890;
w9892 <= w9889 and not w9890;
w9893 <= not w9891 and not w9892;
w9894 <= w141 and w8793;
w9895 <= a(58) and a(60);
w9896 <= w74 and w9895;
w9897 <= w138 and w9315;
w9898 <= not w9896 and not w9897;
w9899 <= not w9894 and not w9898;
w9900 <= a(60) and not w9899;
w9901 <= a(5) and w9900;
w9902 <= not w9894 and not w9899;
w9903 <= a(6) and a(59);
w9904 <= a(7) and a(58);
w9905 <= not w9903 and not w9904;
w9906 <= w9902 and not w9905;
w9907 <= not w9901 and not w9906;
w9908 <= not w9893 and not w9907;
w9909 <= w9893 and w9907;
w9910 <= not w9908 and not w9909;
w9911 <= w9877 and w9910;
w9912 <= not w9877 and not w9910;
w9913 <= not w9911 and not w9912;
w9914 <= not w9838 and not w9913;
w9915 <= not w9838 and not w9914;
w9916 <= not w9913 and not w9914;
w9917 <= not w9915 and not w9916;
w9918 <= not w9790 and not w9917;
w9919 <= not w9790 and not w9918;
w9920 <= not w9917 and not w9918;
w9921 <= not w9919 and not w9920;
w9922 <= not w9575 and not w9578;
w9923 <= not w9389 and not w9392;
w9924 <= w9922 and w9923;
w9925 <= not w9922 and not w9923;
w9926 <= not w9924 and not w9925;
w9927 <= not w9395 and not w9398;
w9928 <= not w9926 and w9927;
w9929 <= w9926 and not w9927;
w9930 <= not w9928 and not w9929;
w9931 <= not w9401 and not w9403;
w9932 <= not w9582 and not w9586;
w9933 <= not w9931 and w9932;
w9934 <= w9931 and not w9932;
w9935 <= not w9933 and not w9934;
w9936 <= w9930 and not w9935;
w9937 <= not w9930 and w9935;
w9938 <= not w9936 and not w9937;
w9939 <= not w9921 and w9938;
w9940 <= not w9921 and not w9939;
w9941 <= w9938 and not w9939;
w9942 <= not w9940 and not w9941;
w9943 <= not w9789 and w9942;
w9944 <= w9789 and not w9942;
w9945 <= not w9943 and not w9944;
w9946 <= w9707 and not w9945;
w9947 <= not w9707 and w9945;
w9948 <= not w9946 and not w9947;
w9949 <= not w9666 and w9948;
w9950 <= w9666 and not w9948;
w9951 <= not w9949 and not w9950;
w9952 <= not w9665 and not w9951;
w9953 <= w9665 and w9951;
w9954 <= not w9952 and not w9953;
w9955 <= not w9665 and not w9950;
w9956 <= not w9949 and not w9955;
w9957 <= not w9706 and not w9946;
w9958 <= not w9789 and not w9942;
w9959 <= not w9786 and not w9958;
w9960 <= not w9778 and not w9782;
w9961 <= w9733 and w9799;
w9962 <= not w9733 and not w9799;
w9963 <= not w9961 and not w9962;
w9964 <= w9815 and not w9963;
w9965 <= not w9815 and w9963;
w9966 <= not w9964 and not w9965;
w9967 <= not w9889 and not w9890;
w9968 <= not w9908 and not w9967;
w9969 <= not w9966 and w9968;
w9970 <= w9966 and not w9968;
w9971 <= not w9969 and not w9970;
w9972 <= not w9818 and not w9835;
w9973 <= not w9971 and w9972;
w9974 <= w9971 and not w9972;
w9975 <= not w9973 and not w9974;
w9976 <= not w9877 and w9910;
w9977 <= not w9914 and not w9976;
w9978 <= not w9713 and not w9759;
w9979 <= w9977 and w9978;
w9980 <= not w9977 and not w9978;
w9981 <= not w9979 and not w9980;
w9982 <= w9975 and w9981;
w9983 <= not w9975 and not w9981;
w9984 <= not w9982 and not w9983;
w9985 <= not w9960 and w9984;
w9986 <= not w9960 and not w9985;
w9987 <= w9984 and not w9985;
w9988 <= not w9986 and not w9987;
w9989 <= not w9931 and not w9932;
w9990 <= not w9936 and not w9989;
w9991 <= not w9716 and not w9722;
w9992 <= w9829 and w9991;
w9993 <= not w9829 and not w9991;
w9994 <= not w9992 and not w9993;
w9995 <= w186 and w8793;
w9996 <= w118 and w9895;
w9997 <= w141 and w9315;
w9998 <= not w9996 and not w9997;
w9999 <= not w9995 and not w9998;
w10000 <= a(60) and not w9999;
w10001 <= a(6) and w10000;
w10002 <= not w9995 and not w9999;
w10003 <= a(7) and a(59);
w10004 <= a(8) and a(58);
w10005 <= not w10003 and not w10004;
w10006 <= w10002 and not w10005;
w10007 <= not w10001 and not w10006;
w10008 <= w9994 and not w10007;
w10009 <= w9994 and not w10008;
w10010 <= not w10007 and not w10008;
w10011 <= not w10009 and not w10010;
w10012 <= not w9725 and not w9755;
w10013 <= not w9752 and not w10012;
w10014 <= not w10011 and not w10013;
w10015 <= not w10011 and not w10014;
w10016 <= not w10013 and not w10014;
w10017 <= not w10015 and not w10016;
w10018 <= not w9925 and not w9929;
w10019 <= w10017 and w10018;
w10020 <= not w10017 and not w10018;
w10021 <= not w10019 and not w10020;
w10022 <= w9857 and w9871;
w10023 <= not w9857 and not w9871;
w10024 <= not w10022 and not w10023;
w10025 <= w9749 and not w10024;
w10026 <= not w9749 and w10024;
w10027 <= not w10025 and not w10026;
w10028 <= w9887 and w9902;
w10029 <= not w9887 and not w9902;
w10030 <= not w10028 and not w10029;
w10031 <= w9846 and not w10030;
w10032 <= not w9846 and w10030;
w10033 <= not w10031 and not w10032;
w10034 <= not w9861 and not w9874;
w10035 <= not w10033 and w10034;
w10036 <= w10033 and not w10034;
w10037 <= not w10035 and not w10036;
w10038 <= w10027 and w10037;
w10039 <= not w10027 and not w10037;
w10040 <= not w10038 and not w10039;
w10041 <= w10021 and w10040;
w10042 <= not w10021 and not w10040;
w10043 <= not w10041 and not w10042;
w10044 <= not w9990 and w10043;
w10045 <= w9990 and not w10043;
w10046 <= not w10044 and not w10045;
w10047 <= not w9988 and w10046;
w10048 <= w10046 and not w10047;
w10049 <= not w9988 and not w10047;
w10050 <= not w10048 and not w10049;
w10051 <= not w9959 and not w10050;
w10052 <= not w9959 and not w10051;
w10053 <= not w10050 and not w10051;
w10054 <= not w10052 and not w10053;
w10055 <= not w9699 and not w9702;
w10056 <= not w9918 and not w9939;
w10057 <= w10055 and w10056;
w10058 <= not w10055 and not w10056;
w10059 <= not w10057 and not w10058;
w10060 <= not w9674 and not w9697;
w10061 <= w32 and w9527;
w10062 <= w106 and w9715;
w10063 <= w15 and w9598;
w10064 <= not w10062 and not w10063;
w10065 <= not w10061 and not w10064;
w10066 <= not w10061 and not w10065;
w10067 <= a(4) and a(62);
w10068 <= not w8713 and not w10067;
w10069 <= w10066 and not w10068;
w10070 <= a(63) and not w10065;
w10071 <= a(3) and w10070;
w10072 <= not w10069 and not w10071;
w10073 <= w2140 and w4371;
w10074 <= w1847 and w5236;
w10075 <= w2137 and w4889;
w10076 <= not w10074 and not w10075;
w10077 <= not w10073 and not w10076;
w10078 <= a(39) and not w10077;
w10079 <= a(27) and w10078;
w10080 <= a(28) and a(38);
w10081 <= a(29) and a(37);
w10082 <= not w10080 and not w10081;
w10083 <= not w10073 and not w10077;
w10084 <= not w10082 and w10083;
w10085 <= not w10079 and not w10084;
w10086 <= not w10072 and not w10085;
w10087 <= not w10072 and not w10086;
w10088 <= not w10085 and not w10086;
w10089 <= not w10087 and not w10088;
w10090 <= a(19) and a(47);
w10091 <= a(12) and a(54);
w10092 <= w10090 and w10091;
w10093 <= w408 and w7507;
w10094 <= w7866 and w8018;
w10095 <= not w10093 and not w10094;
w10096 <= not w10092 and not w10095;
w10097 <= a(55) and not w10096;
w10098 <= a(11) and w10097;
w10099 <= not w10092 and not w10096;
w10100 <= not w10090 and not w10091;
w10101 <= w10099 and not w10100;
w10102 <= not w10098 and not w10101;
w10103 <= not w10089 and not w10102;
w10104 <= not w10089 and not w10103;
w10105 <= not w10102 and not w10103;
w10106 <= not w10104 and not w10105;
w10107 <= a(24) and a(57);
w10108 <= w5986 and w10107;
w10109 <= a(43) and a(57);
w10110 <= a(23) and w10109;
w10111 <= a(9) and w10110;
w10112 <= w1472 and w4824;
w10113 <= not w10111 and not w10112;
w10114 <= not w10108 and not w10113;
w10115 <= not w10108 and not w10114;
w10116 <= a(9) and a(57);
w10117 <= a(24) and a(42);
w10118 <= not w10116 and not w10117;
w10119 <= w10115 and not w10118;
w10120 <= a(43) and not w10114;
w10121 <= a(23) and w10120;
w10122 <= not w10119 and not w10121;
w10123 <= w1380 and w5519;
w10124 <= w1499 and w7553;
w10125 <= w1300 and w5366;
w10126 <= not w10124 and not w10125;
w10127 <= not w10123 and not w10126;
w10128 <= a(46) and not w10127;
w10129 <= a(20) and w10128;
w10130 <= a(21) and a(45);
w10131 <= a(22) and a(44);
w10132 <= not w10130 and not w10131;
w10133 <= not w10123 and not w10127;
w10134 <= not w10132 and w10133;
w10135 <= not w10129 and not w10134;
w10136 <= not w10122 and not w10135;
w10137 <= not w10122 and not w10136;
w10138 <= not w10135 and not w10136;
w10139 <= not w10137 and not w10138;
w10140 <= a(25) and a(41);
w10141 <= a(26) and a(40);
w10142 <= not w10140 and not w10141;
w10143 <= w2269 and w5219;
w10144 <= a(56) and not w10143;
w10145 <= a(10) and w10144;
w10146 <= not w10142 and w10145;
w10147 <= a(56) and not w10146;
w10148 <= a(10) and w10147;
w10149 <= not w10143 and not w10146;
w10150 <= not w10142 and w10149;
w10151 <= not w10148 and not w10150;
w10152 <= not w10139 and not w10151;
w10153 <= not w10139 and not w10152;
w10154 <= not w10151 and not w10152;
w10155 <= not w10153 and not w10154;
w10156 <= a(13) and a(53);
w10157 <= a(15) and a(51);
w10158 <= not w10156 and not w10157;
w10159 <= w627 and w7038;
w10160 <= a(48) and not w10159;
w10161 <= a(18) and w10160;
w10162 <= not w10158 and w10161;
w10163 <= not w10159 and not w10162;
w10164 <= not w10158 and w10163;
w10165 <= a(48) and not w10162;
w10166 <= a(18) and w10165;
w10167 <= not w10164 and not w10166;
w10168 <= a(31) and a(35);
w10169 <= not w3833 and not w10168;
w10170 <= w2671 and w3634;
w10171 <= a(52) and not w10170;
w10172 <= a(14) and w10171;
w10173 <= not w10169 and w10172;
w10174 <= a(52) and not w10173;
w10175 <= a(14) and w10174;
w10176 <= not w10170 and not w10173;
w10177 <= not w10169 and w10176;
w10178 <= not w10175 and not w10177;
w10179 <= not w10167 and not w10178;
w10180 <= not w10167 and not w10179;
w10181 <= not w10178 and not w10179;
w10182 <= not w10180 and not w10181;
w10183 <= not w6869 and not w7448;
w10184 <= w854 and w6131;
w10185 <= w3896 and not w10184;
w10186 <= not w10183 and w10185;
w10187 <= w3896 and not w10186;
w10188 <= not w10184 and not w10186;
w10189 <= not w10183 and w10188;
w10190 <= not w10187 and not w10189;
w10191 <= not w10182 and not w10190;
w10192 <= not w10182 and not w10191;
w10193 <= not w10190 and not w10191;
w10194 <= not w10192 and not w10193;
w10195 <= not w10155 and w10194;
w10196 <= w10155 and not w10194;
w10197 <= not w10195 and not w10196;
w10198 <= not w10106 and not w10197;
w10199 <= w10106 and w10197;
w10200 <= not w10198 and not w10199;
w10201 <= not w10060 and w10200;
w10202 <= w10060 and not w10200;
w10203 <= not w10201 and not w10202;
w10204 <= not w9679 and not w9682;
w10205 <= not w9685 and not w9688;
w10206 <= w10204 and w10205;
w10207 <= not w10204 and not w10205;
w10208 <= not w10206 and not w10207;
w10209 <= not w9764 and not w9767;
w10210 <= not w10208 and w10209;
w10211 <= w10208 and not w10209;
w10212 <= not w10210 and not w10211;
w10213 <= not w9691 and not w9693;
w10214 <= not w9771 and not w9775;
w10215 <= not w10213 and w10214;
w10216 <= w10213 and not w10214;
w10217 <= not w10215 and not w10216;
w10218 <= w10212 and not w10217;
w10219 <= not w10212 and w10217;
w10220 <= not w10218 and not w10219;
w10221 <= w10203 and w10220;
w10222 <= not w10203 and not w10220;
w10223 <= not w10221 and not w10222;
w10224 <= w10059 and w10223;
w10225 <= not w10059 and not w10223;
w10226 <= not w10054 and not w10225;
w10227 <= not w10224 and w10226;
w10228 <= not w10054 and not w10227;
w10229 <= not w10225 and not w10227;
w10230 <= not w10224 and w10229;
w10231 <= not w10228 and not w10230;
w10232 <= not w9957 and not w10231;
w10233 <= w9957 and w10231;
w10234 <= not w10232 and not w10233;
w10235 <= not w9956 and w10234;
w10236 <= w9956 and not w10234;
w10237 <= not w10235 and not w10236;
w10238 <= not w10051 and not w10227;
w10239 <= not w9985 and not w10047;
w10240 <= not w10201 and not w10221;
w10241 <= w10239 and w10240;
w10242 <= not w10239 and not w10240;
w10243 <= not w10241 and not w10242;
w10244 <= not w9980 and not w9982;
w10245 <= a(48) and a(53);
w10246 <= a(14) and w10245;
w10247 <= a(17) and w5694;
w10248 <= not w10246 and not w10247;
w10249 <= a(14) and a(53);
w10250 <= w7131 and w10249;
w10251 <= a(19) and not w10250;
w10252 <= not w10248 and w10251;
w10253 <= not w10250 and not w10252;
w10254 <= not w7131 and not w10249;
w10255 <= w10253 and not w10254;
w10256 <= a(48) and not w10252;
w10257 <= a(19) and w10256;
w10258 <= not w10255 and not w10257;
w10259 <= w2269 and w5150;
w10260 <= a(25) and a(46);
w10261 <= w9333 and w10260;
w10262 <= not w10259 and not w10261;
w10263 <= a(21) and a(46);
w10264 <= a(26) and a(41);
w10265 <= w10263 and w10264;
w10266 <= not w10262 and not w10265;
w10267 <= a(42) and not w10266;
w10268 <= a(25) and w10267;
w10269 <= not w10265 and not w10266;
w10270 <= not w10263 and not w10264;
w10271 <= w10269 and not w10270;
w10272 <= not w10268 and not w10271;
w10273 <= not w10258 and not w10272;
w10274 <= not w10258 and not w10273;
w10275 <= not w10272 and not w10273;
w10276 <= not w10274 and not w10275;
w10277 <= a(27) and a(40);
w10278 <= a(28) and a(39);
w10279 <= not w10277 and not w10278;
w10280 <= w2137 and w3977;
w10281 <= a(4) and not w10280;
w10282 <= a(63) and w10281;
w10283 <= not w10279 and w10282;
w10284 <= a(63) and not w10283;
w10285 <= a(4) and w10284;
w10286 <= not w10280 and not w10283;
w10287 <= not w10279 and w10286;
w10288 <= not w10285 and not w10287;
w10289 <= not w10276 and not w10288;
w10290 <= not w10276 and not w10289;
w10291 <= not w10288 and not w10289;
w10292 <= not w10290 and not w10291;
w10293 <= a(5) and a(62);
w10294 <= not a(34) and not w10293;
w10295 <= a(62) and w3470;
w10296 <= a(18) and a(49);
w10297 <= not w10294 and not w10295;
w10298 <= w10296 and w10297;
w10299 <= not w10295 and not w10298;
w10300 <= not w10294 and w10299;
w10301 <= w10296 and not w10298;
w10302 <= not w10300 and not w10301;
w10303 <= w2949 and w3125;
w10304 <= w3942 and w3956;
w10305 <= w3618 and w3634;
w10306 <= not w10304 and not w10305;
w10307 <= not w10303 and not w10306;
w10308 <= w3942 and not w10307;
w10309 <= not w10303 and not w10307;
w10310 <= not w3956 and not w6629;
w10311 <= w10309 and not w10310;
w10312 <= not w10308 and not w10311;
w10313 <= not w10302 and not w10312;
w10314 <= not w10302 and not w10313;
w10315 <= not w10312 and not w10313;
w10316 <= not w10314 and not w10315;
w10317 <= a(29) and a(38);
w10318 <= a(12) and a(55);
w10319 <= a(13) and a(54);
w10320 <= not w10318 and not w10319;
w10321 <= w554 and w7507;
w10322 <= w10317 and not w10321;
w10323 <= not w10320 and w10322;
w10324 <= w10317 and not w10323;
w10325 <= not w10321 and not w10323;
w10326 <= not w10320 and w10325;
w10327 <= not w10324 and not w10326;
w10328 <= not w10316 and not w10327;
w10329 <= not w10316 and not w10328;
w10330 <= not w10327 and not w10328;
w10331 <= not w10329 and not w10330;
w10332 <= a(8) and a(59);
w10333 <= a(9) and a(58);
w10334 <= not w10332 and not w10333;
w10335 <= w238 and w8793;
w10336 <= w569 and w9895;
w10337 <= w186 and w9315;
w10338 <= not w10336 and not w10337;
w10339 <= not w10335 and not w10338;
w10340 <= not w10335 and not w10339;
w10341 <= not w10334 and w10340;
w10342 <= a(60) and not w10339;
w10343 <= a(7) and w10342;
w10344 <= not w10341 and not w10343;
w10345 <= w1472 and w5102;
w10346 <= w1921 and w4617;
w10347 <= w1725 and w5519;
w10348 <= not w10346 and not w10347;
w10349 <= not w10345 and not w10348;
w10350 <= a(45) and not w10349;
w10351 <= a(22) and w10350;
w10352 <= not w10345 and not w10349;
w10353 <= a(23) and a(44);
w10354 <= a(24) and a(43);
w10355 <= not w10353 and not w10354;
w10356 <= w10352 and not w10355;
w10357 <= not w10351 and not w10356;
w10358 <= not w10344 and not w10357;
w10359 <= not w10344 and not w10358;
w10360 <= not w10357 and not w10358;
w10361 <= not w10359 and not w10360;
w10362 <= a(37) and a(52);
w10363 <= a(30) and w10362;
w10364 <= a(15) and w10363;
w10365 <= w697 and w6774;
w10366 <= not w10364 and not w10365;
w10367 <= a(16) and a(51);
w10368 <= a(30) and a(37);
w10369 <= w10367 and w10368;
w10370 <= not w10366 and not w10369;
w10371 <= a(52) and not w10370;
w10372 <= a(15) and w10371;
w10373 <= not w10367 and not w10368;
w10374 <= not w10369 and not w10370;
w10375 <= not w10373 and w10374;
w10376 <= not w10372 and not w10375;
w10377 <= not w10361 and not w10376;
w10378 <= not w10361 and not w10377;
w10379 <= not w10376 and not w10377;
w10380 <= not w10378 and not w10379;
w10381 <= not w10331 and w10380;
w10382 <= w10331 and not w10380;
w10383 <= not w10381 and not w10382;
w10384 <= not w10292 and not w10383;
w10385 <= w10292 and w10383;
w10386 <= not w10384 and not w10385;
w10387 <= not w10244 and w10386;
w10388 <= w10244 and not w10386;
w10389 <= not w10387 and not w10388;
w10390 <= not w10029 and not w10032;
w10391 <= not w9962 and not w9965;
w10392 <= w10390 and w10391;
w10393 <= not w10390 and not w10391;
w10394 <= not w10392 and not w10393;
w10395 <= not w10023 and not w10026;
w10396 <= not w10394 and w10395;
w10397 <= w10394 and not w10395;
w10398 <= not w10396 and not w10397;
w10399 <= not w10036 and not w10038;
w10400 <= not w9970 and not w9974;
w10401 <= w10399 and w10400;
w10402 <= not w10399 and not w10400;
w10403 <= not w10401 and not w10402;
w10404 <= w10398 and w10403;
w10405 <= not w10398 and not w10403;
w10406 <= not w10404 and not w10405;
w10407 <= w10389 and w10406;
w10408 <= not w10389 and not w10406;
w10409 <= not w10407 and not w10408;
w10410 <= w10243 and w10409;
w10411 <= not w10243 and not w10409;
w10412 <= not w10058 and not w10224;
w10413 <= not w10041 and not w10044;
w10414 <= not w10213 and not w10214;
w10415 <= not w10218 and not w10414;
w10416 <= not w10136 and not w10152;
w10417 <= not w9993 and not w10008;
w10418 <= w10416 and w10417;
w10419 <= not w10416 and not w10417;
w10420 <= not w10418 and not w10419;
w10421 <= not w10086 and not w10103;
w10422 <= not w10420 and w10421;
w10423 <= w10420 and not w10421;
w10424 <= not w10422 and not w10423;
w10425 <= w10002 and w10066;
w10426 <= not w10002 and not w10066;
w10427 <= not w10425 and not w10426;
w10428 <= w10083 and not w10427;
w10429 <= not w10083 and w10427;
w10430 <= not w10428 and not w10429;
w10431 <= w10115 and w10149;
w10432 <= not w10115 and not w10149;
w10433 <= not w10431 and not w10432;
w10434 <= w10133 and not w10433;
w10435 <= not w10133 and w10433;
w10436 <= not w10434 and not w10435;
w10437 <= a(6) and a(61);
w10438 <= not w10188 and w10437;
w10439 <= w10188 and not w10437;
w10440 <= not w10438 and not w10439;
w10441 <= w10176 and not w10440;
w10442 <= not w10176 and w10440;
w10443 <= not w10441 and not w10442;
w10444 <= w10436 and w10443;
w10445 <= not w10436 and not w10443;
w10446 <= not w10444 and not w10445;
w10447 <= w10430 and w10446;
w10448 <= not w10430 and not w10446;
w10449 <= not w10447 and not w10448;
w10450 <= w10424 and w10449;
w10451 <= not w10424 and not w10449;
w10452 <= not w10450 and not w10451;
w10453 <= not w10415 and w10452;
w10454 <= w10415 and not w10452;
w10455 <= not w10453 and not w10454;
w10456 <= w10413 and not w10455;
w10457 <= not w10413 and w10455;
w10458 <= not w10456 and not w10457;
w10459 <= w10099 and w10163;
w10460 <= not w10099 and not w10163;
w10461 <= not w10459 and not w10460;
w10462 <= w7866 and w9791;
w10463 <= w529 and w8006;
w10464 <= a(20) and a(57);
w10465 <= w7536 and w10464;
w10466 <= not w10463 and not w10465;
w10467 <= not w10462 and not w10466;
w10468 <= a(57) and not w10467;
w10469 <= a(10) and w10468;
w10470 <= not w10462 and not w10467;
w10471 <= a(11) and a(56);
w10472 <= a(20) and a(47);
w10473 <= not w10471 and not w10472;
w10474 <= w10470 and not w10473;
w10475 <= not w10469 and not w10474;
w10476 <= w10461 and not w10475;
w10477 <= w10461 and not w10476;
w10478 <= not w10475 and not w10476;
w10479 <= not w10477 and not w10478;
w10480 <= not w10179 and not w10191;
w10481 <= w10479 and w10480;
w10482 <= not w10479 and not w10480;
w10483 <= not w10481 and not w10482;
w10484 <= not w10207 and not w10211;
w10485 <= not w10483 and w10484;
w10486 <= w10483 and not w10484;
w10487 <= not w10485 and not w10486;
w10488 <= not w10155 and not w10194;
w10489 <= not w10198 and not w10488;
w10490 <= not w10014 and not w10020;
w10491 <= w10489 and w10490;
w10492 <= not w10489 and not w10490;
w10493 <= not w10491 and not w10492;
w10494 <= w10487 and w10493;
w10495 <= not w10487 and not w10493;
w10496 <= not w10494 and not w10495;
w10497 <= w10458 and w10496;
w10498 <= not w10458 and not w10496;
w10499 <= not w10497 and not w10498;
w10500 <= not w10412 and w10499;
w10501 <= w10412 and not w10499;
w10502 <= not w10500 and not w10501;
w10503 <= not w10411 and w10502;
w10504 <= not w10410 and w10503;
w10505 <= w10502 and not w10504;
w10506 <= not w10411 and not w10504;
w10507 <= not w10410 and w10506;
w10508 <= not w10505 and not w10507;
w10509 <= not w10238 and not w10508;
w10510 <= w10238 and w10508;
w10511 <= not w10509 and not w10510;
w10512 <= not w9956 and not w10233;
w10513 <= not w10232 and not w10512;
w10514 <= not w10511 and w10513;
w10515 <= w10511 and not w10513;
w10516 <= not w10514 and not w10515;
w10517 <= not w10242 and not w10410;
w10518 <= not w10450 and not w10453;
w10519 <= not w10331 and not w10380;
w10520 <= not w10384 and not w10519;
w10521 <= not w10460 and not w10476;
w10522 <= not w10432 and not w10435;
w10523 <= w10521 and w10522;
w10524 <= not w10521 and not w10522;
w10525 <= not w10523 and not w10524;
w10526 <= not w10358 and not w10377;
w10527 <= not w10525 and w10526;
w10528 <= w10525 and not w10526;
w10529 <= not w10527 and not w10528;
w10530 <= w186 and w9318;
w10531 <= a(60) and not w10530;
w10532 <= a(8) and w10531;
w10533 <= a(7) and not w10530;
w10534 <= a(61) and w10533;
w10535 <= not w10532 and not w10534;
w10536 <= not w10299 and not w10535;
w10537 <= not w10299 and not w10536;
w10538 <= not w10535 and not w10536;
w10539 <= not w10537 and not w10538;
w10540 <= not w10438 and not w10442;
w10541 <= w10539 and w10540;
w10542 <= not w10539 and not w10540;
w10543 <= not w10541 and not w10542;
w10544 <= not w10426 and not w10429;
w10545 <= not w10543 and w10544;
w10546 <= w10543 and not w10544;
w10547 <= not w10545 and not w10546;
w10548 <= w10529 and w10547;
w10549 <= not w10529 and not w10547;
w10550 <= not w10548 and not w10549;
w10551 <= not w10520 and w10550;
w10552 <= w10520 and not w10550;
w10553 <= not w10551 and not w10552;
w10554 <= not w10518 and w10553;
w10555 <= not w10518 and not w10554;
w10556 <= w10553 and not w10554;
w10557 <= not w10555 and not w10556;
w10558 <= not w10402 and not w10404;
w10559 <= w10253 and w10269;
w10560 <= not w10253 and not w10269;
w10561 <= not w10559 and not w10560;
w10562 <= w10325 and not w10561;
w10563 <= not w10325 and w10561;
w10564 <= not w10562 and not w10563;
w10565 <= not w10273 and not w10289;
w10566 <= not w10313 and not w10328;
w10567 <= w10565 and w10566;
w10568 <= not w10565 and not w10566;
w10569 <= not w10567 and not w10568;
w10570 <= w10564 and w10569;
w10571 <= not w10564 and not w10569;
w10572 <= not w10570 and not w10571;
w10573 <= not w10393 and not w10397;
w10574 <= w10352 and w10470;
w10575 <= not w10352 and not w10470;
w10576 <= not w10574 and not w10575;
w10577 <= w10340 and not w10576;
w10578 <= not w10340 and w10576;
w10579 <= not w10577 and not w10578;
w10580 <= w10286 and w10309;
w10581 <= not w10286 and not w10309;
w10582 <= not w10580 and not w10581;
w10583 <= w10374 and not w10582;
w10584 <= not w10374 and w10582;
w10585 <= not w10583 and not w10584;
w10586 <= w10579 and w10585;
w10587 <= not w10579 and not w10585;
w10588 <= not w10586 and not w10587;
w10589 <= not w10573 and w10588;
w10590 <= w10573 and not w10588;
w10591 <= not w10589 and not w10590;
w10592 <= w10572 and w10591;
w10593 <= not w10572 and not w10591;
w10594 <= not w10592 and not w10593;
w10595 <= not w10558 and w10594;
w10596 <= w10558 and not w10594;
w10597 <= not w10595 and not w10596;
w10598 <= not w10557 and w10597;
w10599 <= w10597 and not w10598;
w10600 <= not w10557 and not w10598;
w10601 <= not w10599 and not w10600;
w10602 <= not w10517 and not w10601;
w10603 <= not w10517 and not w10602;
w10604 <= not w10601 and not w10602;
w10605 <= not w10603 and not w10604;
w10606 <= not w10457 and not w10497;
w10607 <= not w10387 and not w10407;
w10608 <= not w10492 and not w10494;
w10609 <= not w10444 and not w10447;
w10610 <= not w10419 and not w10423;
w10611 <= w10609 and w10610;
w10612 <= not w10609 and not w10610;
w10613 <= not w10611 and not w10612;
w10614 <= not w10482 and not w10486;
w10615 <= not w10613 and w10614;
w10616 <= w10613 and not w10614;
w10617 <= not w10615 and not w10616;
w10618 <= w529 and w8242;
w10619 <= w882 and w8791;
w10620 <= w290 and w8793;
w10621 <= not w10619 and not w10620;
w10622 <= not w10618 and not w10621;
w10623 <= not w10618 and not w10622;
w10624 <= a(10) and a(58);
w10625 <= a(11) and a(57);
w10626 <= not w10624 and not w10625;
w10627 <= w10623 and not w10626;
w10628 <= a(59) and not w10622;
w10629 <= a(9) and w10628;
w10630 <= not w10627 and not w10629;
w10631 <= w2140 and w3977;
w10632 <= w1847 and w3790;
w10633 <= w2137 and w5219;
w10634 <= not w10632 and not w10633;
w10635 <= not w10631 and not w10634;
w10636 <= a(41) and not w10635;
w10637 <= a(27) and w10636;
w10638 <= a(28) and a(40);
w10639 <= a(29) and a(39);
w10640 <= not w10638 and not w10639;
w10641 <= not w10631 and not w10635;
w10642 <= not w10640 and w10641;
w10643 <= not w10637 and not w10642;
w10644 <= not w10630 and not w10643;
w10645 <= not w10630 and not w10644;
w10646 <= not w10643 and not w10644;
w10647 <= not w10645 and not w10646;
w10648 <= a(5) and a(63);
w10649 <= a(6) and a(62);
w10650 <= not w10648 and not w10649;
w10651 <= w138 and w9598;
w10652 <= a(47) and not w10651;
w10653 <= a(21) and w10652;
w10654 <= not w10650 and w10653;
w10655 <= a(47) and not w10654;
w10656 <= a(21) and w10655;
w10657 <= not w10651 and not w10654;
w10658 <= not w10650 and w10657;
w10659 <= not w10656 and not w10658;
w10660 <= not w10647 and not w10659;
w10661 <= not w10647 and not w10660;
w10662 <= not w10659 and not w10660;
w10663 <= not w10661 and not w10662;
w10664 <= a(18) and a(50);
w10665 <= a(19) and a(49);
w10666 <= not w10664 and not w10665;
w10667 <= w955 and w6131;
w10668 <= w2778 and not w10667;
w10669 <= not w10666 and w10668;
w10670 <= not w10667 and not w10669;
w10671 <= not w10666 and w10670;
w10672 <= w2778 and not w10669;
w10673 <= not w10671 and not w10672;
w10674 <= w3493 and w3618;
w10675 <= w2294 and w3336;
w10676 <= w2671 and w4371;
w10677 <= not w10675 and not w10676;
w10678 <= not w10674 and not w10677;
w10679 <= a(38) and not w10678;
w10680 <= a(30) and w10679;
w10681 <= not w10674 and not w10678;
w10682 <= a(31) and a(37);
w10683 <= a(32) and a(36);
w10684 <= not w10682 and not w10683;
w10685 <= w10681 and not w10684;
w10686 <= not w10680 and not w10685;
w10687 <= not w10673 and not w10686;
w10688 <= not w10673 and not w10687;
w10689 <= not w10686 and not w10687;
w10690 <= not w10688 and not w10689;
w10691 <= a(12) and a(56);
w10692 <= w7578 and w10691;
w10693 <= w554 and w8967;
w10694 <= not w10692 and not w10693;
w10695 <= a(13) and a(55);
w10696 <= w7578 and w10695;
w10697 <= not w10694 and not w10696;
w10698 <= w10691 and not w10697;
w10699 <= not w10696 and not w10697;
w10700 <= not w7578 and not w10695;
w10701 <= w10699 and not w10700;
w10702 <= not w10698 and not w10701;
w10703 <= not w10690 and not w10702;
w10704 <= not w10690 and not w10703;
w10705 <= not w10702 and not w10703;
w10706 <= not w10704 and not w10705;
w10707 <= a(15) and a(53);
w10708 <= a(16) and a(52);
w10709 <= not w10707 and not w10708;
w10710 <= w697 and w7239;
w10711 <= a(52) and a(54);
w10712 <= w699 and w10711;
w10713 <= w701 and w7505;
w10714 <= not w10712 and not w10713;
w10715 <= not w10710 and not w10714;
w10716 <= not w10710 and not w10715;
w10717 <= not w10709 and w10716;
w10718 <= a(54) and not w10715;
w10719 <= a(14) and w10718;
w10720 <= not w10717 and not w10719;
w10721 <= w1725 and w5366;
w10722 <= a(48) and not w10721;
w10723 <= a(23) and a(45);
w10724 <= a(22) and a(46);
w10725 <= not w10723 and not w10724;
w10726 <= a(20) and not w10725;
w10727 <= w10722 and w10726;
w10728 <= a(48) and not w10727;
w10729 <= a(20) and w10728;
w10730 <= not w10721 and not w10727;
w10731 <= not w10725 and w10730;
w10732 <= not w10729 and not w10731;
w10733 <= not w10720 and not w10732;
w10734 <= not w10720 and not w10733;
w10735 <= not w10732 and not w10733;
w10736 <= not w10734 and not w10735;
w10737 <= w2269 and w4824;
w10738 <= w2107 and w4445;
w10739 <= w1710 and w5102;
w10740 <= not w10738 and not w10739;
w10741 <= not w10737 and not w10740;
w10742 <= a(44) and not w10741;
w10743 <= a(24) and w10742;
w10744 <= not w10737 and not w10741;
w10745 <= a(25) and a(43);
w10746 <= a(26) and a(42);
w10747 <= not w10745 and not w10746;
w10748 <= w10744 and not w10747;
w10749 <= not w10743 and not w10748;
w10750 <= not w10736 and not w10749;
w10751 <= not w10736 and not w10750;
w10752 <= not w10749 and not w10750;
w10753 <= not w10751 and not w10752;
w10754 <= not w10706 and w10753;
w10755 <= w10706 and not w10753;
w10756 <= not w10754 and not w10755;
w10757 <= not w10663 and not w10756;
w10758 <= w10663 and w10756;
w10759 <= not w10757 and not w10758;
w10760 <= w10617 and w10759;
w10761 <= not w10617 and not w10759;
w10762 <= not w10760 and not w10761;
w10763 <= not w10608 and w10762;
w10764 <= w10608 and not w10762;
w10765 <= not w10763 and not w10764;
w10766 <= not w10607 and w10765;
w10767 <= w10607 and not w10765;
w10768 <= not w10766 and not w10767;
w10769 <= not w10606 and w10768;
w10770 <= w10606 and not w10768;
w10771 <= not w10769 and not w10770;
w10772 <= not w10605 and not w10771;
w10773 <= w10605 and w10771;
w10774 <= not w10772 and not w10773;
w10775 <= not w10500 and not w10504;
w10776 <= w10774 and w10775;
w10777 <= not w10774 and not w10775;
w10778 <= not w10776 and not w10777;
w10779 <= not w10510 and not w10513;
w10780 <= not w10509 and not w10779;
w10781 <= not w10778 and w10780;
w10782 <= w10778 and not w10780;
w10783 <= not w10781 and not w10782;
w10784 <= not w10554 and not w10598;
w10785 <= not w10760 and not w10763;
w10786 <= w10784 and w10785;
w10787 <= not w10784 and not w10785;
w10788 <= not w10786 and not w10787;
w10789 <= not w10568 and not w10570;
w10790 <= w858 and w6774;
w10791 <= w2940 and w6772;
w10792 <= w955 and w6370;
w10793 <= not w10791 and not w10792;
w10794 <= not w10790 and not w10793;
w10795 <= not w10790 and not w10794;
w10796 <= a(17) and a(52);
w10797 <= a(18) and a(51);
w10798 <= not w10796 and not w10797;
w10799 <= w10795 and not w10798;
w10800 <= a(50) and not w10794;
w10801 <= a(19) and w10800;
w10802 <= not w10799 and not w10801;
w10803 <= w2423 and w3977;
w10804 <= w2916 and w3790;
w10805 <= w2140 and w5219;
w10806 <= not w10804 and not w10805;
w10807 <= not w10803 and not w10806;
w10808 <= a(41) and not w10807;
w10809 <= a(28) and w10808;
w10810 <= not w10803 and not w10807;
w10811 <= a(29) and a(40);
w10812 <= a(30) and a(39);
w10813 <= not w10811 and not w10812;
w10814 <= w10810 and not w10813;
w10815 <= not w10809 and not w10814;
w10816 <= not w10802 and not w10815;
w10817 <= not w10802 and not w10816;
w10818 <= not w10815 and not w10816;
w10819 <= not w10817 and not w10818;
w10820 <= not w10575 and not w10578;
w10821 <= w10819 and w10820;
w10822 <= not w10819 and not w10820;
w10823 <= not w10821 and not w10822;
w10824 <= a(62) and w3939;
w10825 <= w3125 and not w10824;
w10826 <= not w10824 and not w10825;
w10827 <= a(7) and a(62);
w10828 <= not a(35) and not w10827;
w10829 <= w10826 and not w10828;
w10830 <= w3125 and not w10825;
w10831 <= not w10829 and not w10830;
w10832 <= w2949 and w3493;
w10833 <= w2404 and w3336;
w10834 <= w3618 and w4371;
w10835 <= not w10833 and not w10834;
w10836 <= not w10832 and not w10835;
w10837 <= a(38) and not w10836;
w10838 <= a(31) and w10837;
w10839 <= not w10832 and not w10836;
w10840 <= a(32) and a(37);
w10841 <= not w7177 and not w10840;
w10842 <= w10839 and not w10841;
w10843 <= not w10838 and not w10842;
w10844 <= not w10831 and not w10843;
w10845 <= not w10831 and not w10844;
w10846 <= not w10843 and not w10844;
w10847 <= not w10845 and not w10846;
w10848 <= w697 and w7505;
w10849 <= a(20) and a(54);
w10850 <= w9612 and w10849;
w10851 <= not w10848 and not w10850;
w10852 <= w6720 and w9237;
w10853 <= not w10851 and not w10852;
w10854 <= a(54) and not w10853;
w10855 <= a(15) and w10854;
w10856 <= not w10852 and not w10853;
w10857 <= not w6720 and not w9237;
w10858 <= w10856 and not w10857;
w10859 <= not w10855 and not w10858;
w10860 <= not w10847 and not w10859;
w10861 <= not w10847 and not w10860;
w10862 <= not w10859 and not w10860;
w10863 <= not w10861 and not w10862;
w10864 <= w10823 and not w10863;
w10865 <= not w10823 and w10863;
w10866 <= not w10789 and not w10865;
w10867 <= not w10864 and w10866;
w10868 <= not w10789 and not w10867;
w10869 <= not w10864 and not w10867;
w10870 <= not w10865 and w10869;
w10871 <= not w10868 and not w10870;
w10872 <= not w10548 and not w10551;
w10873 <= not w10871 and not w10872;
w10874 <= not w10871 and not w10873;
w10875 <= not w10872 and not w10873;
w10876 <= not w10874 and not w10875;
w10877 <= w290 and w9315;
w10878 <= w184 and w8711;
w10879 <= w238 and w9318;
w10880 <= not w10878 and not w10879;
w10881 <= not w10877 and not w10880;
w10882 <= not w10877 and not w10881;
w10883 <= a(9) and a(60);
w10884 <= a(10) and a(59);
w10885 <= not w10883 and not w10884;
w10886 <= w10882 and not w10885;
w10887 <= a(61) and not w10881;
w10888 <= a(8) and w10887;
w10889 <= not w10886 and not w10888;
w10890 <= w1710 and w5519;
w10891 <= w1353 and w7553;
w10892 <= w1472 and w5366;
w10893 <= not w10891 and not w10892;
w10894 <= not w10890 and not w10893;
w10895 <= a(46) and not w10894;
w10896 <= a(23) and w10895;
w10897 <= a(24) and a(45);
w10898 <= a(25) and a(44);
w10899 <= not w10897 and not w10898;
w10900 <= not w10890 and not w10894;
w10901 <= not w10899 and w10900;
w10902 <= not w10896 and not w10901;
w10903 <= not w10889 and not w10902;
w10904 <= not w10889 and not w10903;
w10905 <= not w10902 and not w10903;
w10906 <= not w10904 and not w10905;
w10907 <= a(26) and a(43);
w10908 <= a(27) and a(42);
w10909 <= not w10907 and not w10908;
w10910 <= w2033 and w4824;
w10911 <= a(6) and not w10910;
w10912 <= a(63) and w10911;
w10913 <= not w10909 and w10912;
w10914 <= a(63) and not w10913;
w10915 <= a(6) and w10914;
w10916 <= not w10910 and not w10913;
w10917 <= not w10909 and w10916;
w10918 <= not w10915 and not w10917;
w10919 <= not w10906 and not w10918;
w10920 <= not w10906 and not w10919;
w10921 <= not w10918 and not w10919;
w10922 <= not w10920 and not w10921;
w10923 <= not w10524 and not w10528;
w10924 <= w10922 and w10923;
w10925 <= not w10922 and not w10923;
w10926 <= not w10924 and not w10925;
w10927 <= w554 and w8006;
w10928 <= w624 and w7748;
w10929 <= w408 and w8242;
w10930 <= not w10928 and not w10929;
w10931 <= not w10927 and not w10930;
w10932 <= a(58) and not w10931;
w10933 <= a(11) and w10932;
w10934 <= not w10927 and not w10931;
w10935 <= a(12) and a(57);
w10936 <= a(13) and a(56);
w10937 <= not w10935 and not w10936;
w10938 <= w10934 and not w10937;
w10939 <= not w10933 and not w10938;
w10940 <= not w10530 and not w10536;
w10941 <= not w10939 and w10940;
w10942 <= w10939 and not w10940;
w10943 <= not w10941 and not w10942;
w10944 <= a(21) and a(48);
w10945 <= a(22) and a(47);
w10946 <= not w10944 and not w10945;
w10947 <= w1380 and w6058;
w10948 <= a(55) and not w10947;
w10949 <= a(14) and w10948;
w10950 <= not w10946 and w10949;
w10951 <= a(55) and not w10950;
w10952 <= a(14) and w10951;
w10953 <= not w10947 and not w10950;
w10954 <= not w10946 and w10953;
w10955 <= not w10952 and not w10954;
w10956 <= not w10943 and not w10955;
w10957 <= w10943 and w10955;
w10958 <= not w10956 and not w10957;
w10959 <= w10926 and w10958;
w10960 <= not w10926 and not w10958;
w10961 <= not w10876 and not w10960;
w10962 <= not w10959 and w10961;
w10963 <= not w10876 and not w10962;
w10964 <= not w10960 and not w10962;
w10965 <= not w10959 and w10964;
w10966 <= not w10963 and not w10965;
w10967 <= w10788 and not w10966;
w10968 <= not w10788 and w10966;
w10969 <= not w10766 and not w10769;
w10970 <= not w10592 and not w10595;
w10971 <= not w10706 and not w10753;
w10972 <= not w10757 and not w10971;
w10973 <= not w10586 and not w10589;
w10974 <= w10699 and w10744;
w10975 <= not w10699 and not w10744;
w10976 <= not w10974 and not w10975;
w10977 <= w10641 and not w10976;
w10978 <= not w10641 and w10976;
w10979 <= not w10977 and not w10978;
w10980 <= not w10581 and not w10584;
w10981 <= not w10560 and not w10563;
w10982 <= w10980 and w10981;
w10983 <= not w10980 and not w10981;
w10984 <= not w10982 and not w10983;
w10985 <= w10979 and w10984;
w10986 <= not w10979 and not w10984;
w10987 <= not w10985 and not w10986;
w10988 <= not w10973 and w10987;
w10989 <= w10973 and not w10987;
w10990 <= not w10988 and not w10989;
w10991 <= not w10972 and w10990;
w10992 <= w10972 and not w10990;
w10993 <= not w10991 and not w10992;
w10994 <= w10970 and not w10993;
w10995 <= not w10970 and w10993;
w10996 <= not w10994 and not w10995;
w10997 <= not w10612 and not w10616;
w10998 <= not w10687 and not w10703;
w10999 <= not w10733 and not w10750;
w11000 <= w10998 and w10999;
w11001 <= not w10998 and not w10999;
w11002 <= not w11000 and not w11001;
w11003 <= not w10542 and not w10546;
w11004 <= not w11002 and w11003;
w11005 <= w11002 and not w11003;
w11006 <= not w11004 and not w11005;
w11007 <= w10623 and w10657;
w11008 <= not w10623 and not w10657;
w11009 <= not w11007 and not w11008;
w11010 <= w10730 and not w11009;
w11011 <= not w10730 and w11009;
w11012 <= not w11010 and not w11011;
w11013 <= w10670 and w10681;
w11014 <= not w10670 and not w10681;
w11015 <= not w11013 and not w11014;
w11016 <= w10716 and not w11015;
w11017 <= not w10716 and w11015;
w11018 <= not w11016 and not w11017;
w11019 <= not w10644 and not w10660;
w11020 <= not w11018 and w11019;
w11021 <= w11018 and not w11019;
w11022 <= not w11020 and not w11021;
w11023 <= w11012 and w11022;
w11024 <= not w11012 and not w11022;
w11025 <= not w11023 and not w11024;
w11026 <= w11006 and w11025;
w11027 <= not w11006 and not w11025;
w11028 <= not w11026 and not w11027;
w11029 <= w10997 and not w11028;
w11030 <= not w10997 and w11028;
w11031 <= not w11029 and not w11030;
w11032 <= w10996 and w11031;
w11033 <= not w10996 and not w11031;
w11034 <= not w11032 and not w11033;
w11035 <= not w10969 and w11034;
w11036 <= w10969 and not w11034;
w11037 <= not w11035 and not w11036;
w11038 <= not w10968 and w11037;
w11039 <= not w10967 and w11038;
w11040 <= w11037 and not w11039;
w11041 <= not w10968 and not w11039;
w11042 <= not w10967 and w11041;
w11043 <= not w11040 and not w11042;
w11044 <= not w10605 and w10771;
w11045 <= not w10602 and not w11044;
w11046 <= not w11043 and not w11045;
w11047 <= w11043 and w11045;
w11048 <= not w11046 and not w11047;
w11049 <= not w10776 and not w10780;
w11050 <= not w10777 and not w11049;
w11051 <= not w11048 and w11050;
w11052 <= w11048 and not w11050;
w11053 <= not w11051 and not w11052;
w11054 <= not w11047 and not w11050;
w11055 <= not w11046 and not w11054;
w11056 <= not w11035 and not w11039;
w11057 <= not w10995 and not w11032;
w11058 <= w10810 and w10916;
w11059 <= not w10810 and not w10916;
w11060 <= not w11058 and not w11059;
w11061 <= w10900 and not w11060;
w11062 <= not w10900 and w11060;
w11063 <= not w11061 and not w11062;
w11064 <= a(8) and a(62);
w11065 <= w10826 and not w11064;
w11066 <= not w10826 and w11064;
w11067 <= not w10839 and not w11066;
w11068 <= not w11065 and w11067;
w11069 <= not w10839 and not w11068;
w11070 <= not w11066 and not w11068;
w11071 <= not w11065 and w11070;
w11072 <= not w11069 and not w11071;
w11073 <= w11063 and not w11072;
w11074 <= w11063 and not w11073;
w11075 <= not w11072 and not w11073;
w11076 <= not w11074 and not w11075;
w11077 <= not w10816 and not w10822;
w11078 <= w11076 and w11077;
w11079 <= not w11076 and not w11077;
w11080 <= not w11078 and not w11079;
w11081 <= not w10903 and not w10919;
w11082 <= not w10939 and not w10940;
w11083 <= not w10956 and not w11082;
w11084 <= w11081 and w11083;
w11085 <= not w11081 and not w11083;
w11086 <= not w11084 and not w11085;
w11087 <= not w10844 and not w10860;
w11088 <= not w11086 and w11087;
w11089 <= w11086 and not w11087;
w11090 <= not w11088 and not w11089;
w11091 <= not w10869 and w11090;
w11092 <= w10869 and not w11090;
w11093 <= not w11091 and not w11092;
w11094 <= not w11080 and not w11093;
w11095 <= w11080 and w11093;
w11096 <= not w11057 and not w11095;
w11097 <= not w11094 and w11096;
w11098 <= not w11057 and not w11097;
w11099 <= not w11095 and not w11097;
w11100 <= not w11094 and w11099;
w11101 <= not w11098 and not w11100;
w11102 <= not w11021 and not w11023;
w11103 <= a(7) and a(63);
w11104 <= a(23) and a(47);
w11105 <= not w11103 and not w11104;
w11106 <= w11103 and w11104;
w11107 <= a(42) and not w11106;
w11108 <= a(28) and w11107;
w11109 <= not w11105 and w11108;
w11110 <= not w11106 and not w11109;
w11111 <= not w11105 and w11110;
w11112 <= a(42) and not w11109;
w11113 <= a(28) and w11112;
w11114 <= not w11111 and not w11113;
w11115 <= w2671 and w3977;
w11116 <= w3258 and w3790;
w11117 <= w2423 and w5219;
w11118 <= not w11116 and not w11117;
w11119 <= not w11115 and not w11118;
w11120 <= a(41) and not w11119;
w11121 <= a(29) and w11120;
w11122 <= not w11115 and not w11119;
w11123 <= a(30) and a(40);
w11124 <= a(31) and a(39);
w11125 <= not w11123 and not w11124;
w11126 <= w11122 and not w11125;
w11127 <= not w11121 and not w11126;
w11128 <= not w11114 and not w11127;
w11129 <= not w11114 and not w11128;
w11130 <= not w11127 and not w11128;
w11131 <= not w11129 and not w11130;
w11132 <= not w11014 and not w11017;
w11133 <= w11131 and w11132;
w11134 <= not w11131 and not w11132;
w11135 <= not w11133 and not w11134;
w11136 <= a(14) and a(56);
w11137 <= a(15) and a(55);
w11138 <= not w11136 and not w11137;
w11139 <= w701 and w8967;
w11140 <= a(48) and not w11139;
w11141 <= a(22) and w11140;
w11142 <= not w11138 and w11141;
w11143 <= not w11139 and not w11142;
w11144 <= not w11138 and w11143;
w11145 <= a(48) and not w11142;
w11146 <= a(22) and w11145;
w11147 <= not w11144 and not w11146;
w11148 <= w2033 and w5102;
w11149 <= w2439 and w4617;
w11150 <= w2269 and w5519;
w11151 <= not w11149 and not w11150;
w11152 <= not w11148 and not w11151;
w11153 <= a(45) and not w11152;
w11154 <= a(25) and w11153;
w11155 <= a(26) and a(44);
w11156 <= a(27) and a(43);
w11157 <= not w11155 and not w11156;
w11158 <= not w11148 and not w11152;
w11159 <= not w11157 and w11158;
w11160 <= not w11154 and not w11159;
w11161 <= not w11147 and not w11160;
w11162 <= not w11147 and not w11161;
w11163 <= not w11160 and not w11161;
w11164 <= not w11162 and not w11163;
w11165 <= w1296 and w6370;
w11166 <= w1298 and w9740;
w11167 <= w1300 and w6131;
w11168 <= not w11166 and not w11167;
w11169 <= not w11165 and not w11168;
w11170 <= a(49) and not w11169;
w11171 <= a(21) and w11170;
w11172 <= not w11165 and not w11169;
w11173 <= a(19) and a(51);
w11174 <= a(20) and a(50);
w11175 <= not w11173 and not w11174;
w11176 <= w11172 and not w11175;
w11177 <= not w11171 and not w11176;
w11178 <= not w11164 and not w11177;
w11179 <= not w11164 and not w11178;
w11180 <= not w11177 and not w11178;
w11181 <= not w11179 and not w11180;
w11182 <= w11135 and not w11181;
w11183 <= not w11135 and w11181;
w11184 <= not w11102 and not w11183;
w11185 <= not w11182 and w11184;
w11186 <= not w11102 and not w11185;
w11187 <= not w11182 and not w11185;
w11188 <= not w11183 and w11187;
w11189 <= not w11186 and not w11188;
w11190 <= not w10988 and not w10991;
w11191 <= w529 and w9315;
w11192 <= w882 and w8711;
w11193 <= w290 and w9318;
w11194 <= not w11192 and not w11193;
w11195 <= not w11191 and not w11194;
w11196 <= not w11191 and not w11195;
w11197 <= a(10) and a(60);
w11198 <= a(11) and a(59);
w11199 <= not w11197 and not w11198;
w11200 <= w11196 and not w11199;
w11201 <= a(61) and not w11195;
w11202 <= a(9) and w11201;
w11203 <= not w11200 and not w11202;
w11204 <= w854 and w7505;
w11205 <= w856 and w10711;
w11206 <= w858 and w7239;
w11207 <= not w11205 and not w11206;
w11208 <= not w11204 and not w11207;
w11209 <= w8043 and not w11208;
w11210 <= not w11204 and not w11208;
w11211 <= a(16) and a(54);
w11212 <= not w8917 and not w11211;
w11213 <= w11210 and not w11212;
w11214 <= not w11209 and not w11213;
w11215 <= not w11203 and not w11214;
w11216 <= not w11203 and not w11215;
w11217 <= not w11214 and not w11215;
w11218 <= not w11216 and not w11217;
w11219 <= w7973 and w10107;
w11220 <= w554 and w8242;
w11221 <= a(24) and a(58);
w11222 <= w7879 and w11221;
w11223 <= not w11220 and not w11222;
w11224 <= not w11219 and not w11223;
w11225 <= a(58) and not w11224;
w11226 <= a(12) and w11225;
w11227 <= not w11219 and not w11224;
w11228 <= a(13) and a(57);
w11229 <= not w5037 and not w11228;
w11230 <= w11227 and not w11229;
w11231 <= not w11226 and not w11230;
w11232 <= not w11218 and not w11231;
w11233 <= not w11218 and not w11232;
w11234 <= not w11231 and not w11232;
w11235 <= not w11233 and not w11234;
w11236 <= w10795 and w10856;
w11237 <= not w10795 and not w10856;
w11238 <= not w11236 and not w11237;
w11239 <= w3493 and w3956;
w11240 <= w2949 and w4371;
w11241 <= a(34) and a(38);
w11242 <= w10683 and w11241;
w11243 <= not w11240 and not w11242;
w11244 <= not w11239 and not w11243;
w11245 <= a(38) and not w11244;
w11246 <= a(32) and w11245;
w11247 <= not w11239 and not w11244;
w11248 <= a(33) and a(37);
w11249 <= not w4401 and not w11248;
w11250 <= w11247 and not w11249;
w11251 <= not w11246 and not w11250;
w11252 <= w11238 and not w11251;
w11253 <= w11238 and not w11252;
w11254 <= not w11251 and not w11252;
w11255 <= not w11253 and not w11254;
w11256 <= not w10983 and not w10985;
w11257 <= not w11255 and not w11256;
w11258 <= w11255 and w11256;
w11259 <= not w11257 and not w11258;
w11260 <= not w11235 and w11259;
w11261 <= w11235 and not w11259;
w11262 <= not w11260 and not w11261;
w11263 <= not w11190 and w11262;
w11264 <= w11190 and not w11262;
w11265 <= not w11263 and not w11264;
w11266 <= not w11189 and w11265;
w11267 <= not w11189 and not w11266;
w11268 <= w11265 and not w11266;
w11269 <= not w11267 and not w11268;
w11270 <= not w11101 and not w11269;
w11271 <= not w11101 and not w11270;
w11272 <= not w11269 and not w11270;
w11273 <= not w11271 and not w11272;
w11274 <= not w11026 and not w11030;
w11275 <= not w10925 and not w10959;
w11276 <= not w11001 and not w11005;
w11277 <= w10882 and w10934;
w11278 <= not w10882 and not w10934;
w11279 <= not w11277 and not w11278;
w11280 <= w10953 and not w11279;
w11281 <= not w10953 and w11279;
w11282 <= not w11280 and not w11281;
w11283 <= not w11008 and not w11011;
w11284 <= not w10975 and not w10978;
w11285 <= w11283 and w11284;
w11286 <= not w11283 and not w11284;
w11287 <= not w11285 and not w11286;
w11288 <= w11282 and w11287;
w11289 <= not w11282 and not w11287;
w11290 <= not w11288 and not w11289;
w11291 <= not w11276 and w11290;
w11292 <= not w11276 and not w11291;
w11293 <= w11290 and not w11291;
w11294 <= not w11292 and not w11293;
w11295 <= not w11275 and not w11294;
w11296 <= not w11275 and not w11295;
w11297 <= not w11294 and not w11295;
w11298 <= not w11296 and not w11297;
w11299 <= not w11274 and not w11298;
w11300 <= not w11274 and not w11299;
w11301 <= not w11298 and not w11299;
w11302 <= not w11300 and not w11301;
w11303 <= not w10873 and not w10962;
w11304 <= w11302 and w11303;
w11305 <= not w11302 and not w11303;
w11306 <= not w11304 and not w11305;
w11307 <= not w10787 and not w10967;
w11308 <= w11306 and not w11307;
w11309 <= w11306 and not w11308;
w11310 <= not w11307 and not w11308;
w11311 <= not w11309 and not w11310;
w11312 <= not w11273 and not w11311;
w11313 <= w11273 and not w11310;
w11314 <= not w11309 and w11313;
w11315 <= not w11312 and not w11314;
w11316 <= w11056 and not w11315;
w11317 <= not w11056 and w11315;
w11318 <= not w11316 and not w11317;
w11319 <= w11055 and not w11318;
w11320 <= not w11055 and not w11316;
w11321 <= not w11317 and w11320;
w11322 <= not w11319 and not w11321;
w11323 <= not w11317 and not w11320;
w11324 <= not w11308 and not w11312;
w11325 <= not w11263 and not w11266;
w11326 <= not w11237 and not w11252;
w11327 <= w11070 and w11326;
w11328 <= not w11070 and not w11326;
w11329 <= not w11327 and not w11328;
w11330 <= not w11059 and not w11062;
w11331 <= not w11329 and w11330;
w11332 <= w11329 and not w11330;
w11333 <= not w11331 and not w11332;
w11334 <= not w11073 and not w11079;
w11335 <= not w11333 and w11334;
w11336 <= w11333 and not w11334;
w11337 <= not w11335 and not w11336;
w11338 <= not w11257 and not w11260;
w11339 <= not w11337 and w11338;
w11340 <= w11337 and not w11338;
w11341 <= not w11339 and not w11340;
w11342 <= not w11091 and not w11095;
w11343 <= w11341 and not w11342;
w11344 <= not w11341 and w11342;
w11345 <= not w11343 and not w11344;
w11346 <= w11325 and not w11345;
w11347 <= not w11325 and w11345;
w11348 <= not w11346 and not w11347;
w11349 <= not w11097 and not w11270;
w11350 <= not w11348 and w11349;
w11351 <= w11348 and not w11349;
w11352 <= not w11350 and not w11351;
w11353 <= not w11299 and not w11305;
w11354 <= not w11215 and not w11232;
w11355 <= not w11278 and not w11281;
w11356 <= w11354 and w11355;
w11357 <= not w11354 and not w11355;
w11358 <= not w11356 and not w11357;
w11359 <= not w11161 and not w11178;
w11360 <= not w11358 and w11359;
w11361 <= w11358 and not w11359;
w11362 <= not w11360 and not w11361;
w11363 <= not w11187 and w11362;
w11364 <= w11187 and not w11362;
w11365 <= not w11363 and not w11364;
w11366 <= not w11128 and not w11134;
w11367 <= w11196 and w11227;
w11368 <= not w11196 and not w11227;
w11369 <= not w11367 and not w11368;
w11370 <= w11158 and not w11369;
w11371 <= not w11158 and w11369;
w11372 <= not w11370 and not w11371;
w11373 <= w11122 and w11143;
w11374 <= not w11122 and not w11143;
w11375 <= not w11373 and not w11374;
w11376 <= w11110 and not w11375;
w11377 <= not w11110 and w11375;
w11378 <= not w11376 and not w11377;
w11379 <= not w11372 and not w11378;
w11380 <= w11372 and w11378;
w11381 <= not w11379 and not w11380;
w11382 <= not w11366 and w11381;
w11383 <= w11366 and not w11381;
w11384 <= not w11382 and not w11383;
w11385 <= w11365 and w11384;
w11386 <= not w11365 and not w11384;
w11387 <= not w11385 and not w11386;
w11388 <= not w11353 and w11387;
w11389 <= w11353 and not w11387;
w11390 <= not w11388 and not w11389;
w11391 <= not w11291 and not w11295;
w11392 <= a(9) and a(62);
w11393 <= not a(36) and not w11392;
w11394 <= a(36) and a(62);
w11395 <= a(9) and w11394;
w11396 <= a(49) and not w11395;
w11397 <= a(22) and w11396;
w11398 <= not w11393 and w11397;
w11399 <= not w11395 and not w11398;
w11400 <= not w11393 and w11399;
w11401 <= a(49) and not w11398;
w11402 <= a(22) and w11401;
w11403 <= not w11400 and not w11402;
w11404 <= w1296 and w6774;
w11405 <= w1298 and w6772;
w11406 <= w1300 and w6370;
w11407 <= not w11405 and not w11406;
w11408 <= not w11404 and not w11407;
w11409 <= a(50) and not w11408;
w11410 <= a(21) and w11409;
w11411 <= a(19) and a(52);
w11412 <= a(20) and a(51);
w11413 <= not w11411 and not w11412;
w11414 <= not w11404 and not w11408;
w11415 <= not w11413 and w11414;
w11416 <= not w11410 and not w11415;
w11417 <= not w11403 and not w11416;
w11418 <= not w11403 and not w11417;
w11419 <= not w11416 and not w11417;
w11420 <= not w11418 and not w11419;
w11421 <= a(34) and a(37);
w11422 <= w3634 and w11421;
w11423 <= w3634 and w4369;
w11424 <= w3956 and w4371;
w11425 <= not w11423 and not w11424;
w11426 <= not w11422 and not w11425;
w11427 <= w4369 and not w11426;
w11428 <= not w11422 and not w11426;
w11429 <= not w3634 and not w11421;
w11430 <= w11428 and not w11429;
w11431 <= not w11427 and not w11430;
w11432 <= not w11420 and not w11431;
w11433 <= not w11420 and not w11432;
w11434 <= not w11431 and not w11432;
w11435 <= not w11433 and not w11434;
w11436 <= w11210 and w11247;
w11437 <= not w11210 and not w11247;
w11438 <= not w11436 and not w11437;
w11439 <= w184 and w9715;
w11440 <= a(60) and a(63);
w11441 <= w767 and w11440;
w11442 <= w529 and w9318;
w11443 <= not w11441 and not w11442;
w11444 <= not w11439 and not w11443;
w11445 <= a(60) and not w11444;
w11446 <= a(11) and w11445;
w11447 <= a(8) and a(63);
w11448 <= a(10) and a(61);
w11449 <= not w11447 and not w11448;
w11450 <= not w11439 and not w11444;
w11451 <= not w11449 and w11450;
w11452 <= not w11446 and not w11451;
w11453 <= w11438 and not w11452;
w11454 <= w11438 and not w11453;
w11455 <= not w11452 and not w11453;
w11456 <= not w11454 and not w11455;
w11457 <= not w11286 and not w11288;
w11458 <= not w11456 and not w11457;
w11459 <= w11456 and w11457;
w11460 <= not w11458 and not w11459;
w11461 <= not w11435 and w11460;
w11462 <= w11435 and not w11460;
w11463 <= not w11461 and not w11462;
w11464 <= not w11391 and w11463;
w11465 <= w11391 and not w11463;
w11466 <= not w11464 and not w11465;
w11467 <= not w11085 and not w11089;
w11468 <= w2140 and w4824;
w11469 <= w1847 and w4445;
w11470 <= w2137 and w5102;
w11471 <= not w11469 and not w11470;
w11472 <= not w11468 and not w11471;
w11473 <= not w11468 and not w11472;
w11474 <= a(28) and a(43);
w11475 <= a(29) and a(42);
w11476 <= not w11474 and not w11475;
w11477 <= w11473 and not w11476;
w11478 <= a(44) and not w11472;
w11479 <= a(27) and w11478;
w11480 <= not w11477 and not w11479;
w11481 <= w3618 and w3977;
w11482 <= w2294 and w3790;
w11483 <= w2671 and w5219;
w11484 <= not w11482 and not w11483;
w11485 <= not w11481 and not w11484;
w11486 <= a(41) and not w11485;
w11487 <= a(30) and w11486;
w11488 <= a(31) and a(40);
w11489 <= a(32) and a(39);
w11490 <= not w11488 and not w11489;
w11491 <= not w11481 and not w11485;
w11492 <= not w11490 and w11491;
w11493 <= not w11487 and not w11492;
w11494 <= not w11480 and not w11493;
w11495 <= not w11480 and not w11494;
w11496 <= not w11493 and not w11494;
w11497 <= not w11495 and not w11496;
w11498 <= a(17) and a(54);
w11499 <= not w8370 and not w11498;
w11500 <= w858 and w7505;
w11501 <= a(48) and not w11500;
w11502 <= a(23) and w11501;
w11503 <= not w11499 and w11502;
w11504 <= a(48) and not w11503;
w11505 <= a(23) and w11504;
w11506 <= not w11500 and not w11503;
w11507 <= not w11499 and w11506;
w11508 <= not w11505 and not w11507;
w11509 <= not w11497 and not w11508;
w11510 <= not w11497 and not w11509;
w11511 <= not w11508 and not w11509;
w11512 <= not w11510 and not w11511;
w11513 <= w554 and w8793;
w11514 <= a(58) and not w11513;
w11515 <= a(13) and w11514;
w11516 <= a(59) and not w11513;
w11517 <= a(12) and w11516;
w11518 <= not w11515 and not w11517;
w11519 <= not w11172 and not w11518;
w11520 <= not w11172 and not w11519;
w11521 <= not w11518 and not w11519;
w11522 <= not w11520 and not w11521;
w11523 <= w697 and w8967;
w11524 <= a(55) and a(57);
w11525 <= w699 and w11524;
w11526 <= w701 and w8006;
w11527 <= not w11525 and not w11526;
w11528 <= not w11523 and not w11527;
w11529 <= not w11523 and not w11528;
w11530 <= a(15) and a(56);
w11531 <= a(16) and a(55);
w11532 <= not w11530 and not w11531;
w11533 <= w11529 and not w11532;
w11534 <= a(57) and not w11528;
w11535 <= a(14) and w11534;
w11536 <= not w11533 and not w11535;
w11537 <= w2269 and w5366;
w11538 <= w2107 and w5056;
w11539 <= w1710 and w5472;
w11540 <= not w11538 and not w11539;
w11541 <= not w11537 and not w11540;
w11542 <= a(47) and not w11541;
w11543 <= a(24) and w11542;
w11544 <= not w11537 and not w11541;
w11545 <= a(26) and a(45);
w11546 <= not w10260 and not w11545;
w11547 <= w11544 and not w11546;
w11548 <= not w11543 and not w11547;
w11549 <= not w11536 and not w11548;
w11550 <= not w11536 and not w11549;
w11551 <= not w11548 and not w11549;
w11552 <= not w11550 and not w11551;
w11553 <= not w11522 and w11552;
w11554 <= w11522 and not w11552;
w11555 <= not w11553 and not w11554;
w11556 <= not w11512 and not w11555;
w11557 <= w11512 and w11555;
w11558 <= not w11556 and not w11557;
w11559 <= not w11467 and w11558;
w11560 <= w11467 and not w11558;
w11561 <= not w11559 and not w11560;
w11562 <= w11466 and w11561;
w11563 <= not w11466 and not w11561;
w11564 <= not w11562 and not w11563;
w11565 <= w11390 and w11564;
w11566 <= not w11390 and not w11564;
w11567 <= not w11565 and not w11566;
w11568 <= not w11352 and not w11567;
w11569 <= w11352 and w11567;
w11570 <= not w11568 and not w11569;
w11571 <= w11324 and not w11570;
w11572 <= not w11324 and w11570;
w11573 <= not w11571 and not w11572;
w11574 <= not w11323 and not w11573;
w11575 <= w11323 and w11573;
w11576 <= not w11574 and not w11575;
w11577 <= not w11323 and not w11571;
w11578 <= not w11572 and not w11577;
w11579 <= not w11464 and not w11562;
w11580 <= not w11380 and not w11382;
w11581 <= not w11437 and not w11453;
w11582 <= w2671 and w5150;
w11583 <= w3258 and w4613;
w11584 <= w2423 and w4824;
w11585 <= not w11583 and not w11584;
w11586 <= not w11582 and not w11585;
w11587 <= a(43) and not w11586;
w11588 <= a(29) and w11587;
w11589 <= a(30) and a(42);
w11590 <= not w4765 and not w11589;
w11591 <= not w11582 and not w11586;
w11592 <= not w11590 and w11591;
w11593 <= not w11588 and not w11592;
w11594 <= not w11581 and not w11593;
w11595 <= not w11581 and not w11594;
w11596 <= not w11593 and not w11594;
w11597 <= not w11595 and not w11596;
w11598 <= not w11374 and not w11377;
w11599 <= w11597 and w11598;
w11600 <= not w11597 and not w11598;
w11601 <= not w11599 and not w11600;
w11602 <= not w11580 and w11601;
w11603 <= w11580 and not w11601;
w11604 <= not w11602 and not w11603;
w11605 <= not w11458 and not w11461;
w11606 <= not w11604 and w11605;
w11607 <= w11604 and not w11605;
w11608 <= not w11606 and not w11607;
w11609 <= not w11363 and not w11385;
w11610 <= w11608 and not w11609;
w11611 <= not w11608 and w11609;
w11612 <= not w11610 and not w11611;
w11613 <= w11579 and not w11612;
w11614 <= not w11579 and w11612;
w11615 <= not w11613 and not w11614;
w11616 <= not w11388 and not w11565;
w11617 <= not w11615 and w11616;
w11618 <= w11615 and not w11616;
w11619 <= not w11617 and not w11618;
w11620 <= not w11343 and not w11347;
w11621 <= not w11494 and not w11509;
w11622 <= not w11368 and not w11371;
w11623 <= w11621 and w11622;
w11624 <= not w11621 and not w11622;
w11625 <= not w11623 and not w11624;
w11626 <= not w11417 and not w11432;
w11627 <= not w11625 and w11626;
w11628 <= w11625 and not w11626;
w11629 <= not w11627 and not w11628;
w11630 <= not w11556 and not w11559;
w11631 <= not w11629 and w11630;
w11632 <= w11629 and not w11630;
w11633 <= not w11631 and not w11632;
w11634 <= not w11522 and not w11552;
w11635 <= not w11549 and not w11634;
w11636 <= w11473 and w11506;
w11637 <= not w11473 and not w11506;
w11638 <= not w11636 and not w11637;
w11639 <= w11491 and not w11638;
w11640 <= not w11491 and w11638;
w11641 <= not w11639 and not w11640;
w11642 <= w11399 and w11428;
w11643 <= not w11399 and not w11428;
w11644 <= not w11642 and not w11643;
w11645 <= w11414 and not w11644;
w11646 <= not w11414 and w11644;
w11647 <= not w11645 and not w11646;
w11648 <= w11641 and w11647;
w11649 <= not w11641 and not w11647;
w11650 <= not w11648 and not w11649;
w11651 <= not w11635 and w11650;
w11652 <= w11635 and not w11650;
w11653 <= not w11651 and not w11652;
w11654 <= w11633 and w11653;
w11655 <= not w11633 and not w11653;
w11656 <= not w11654 and not w11655;
w11657 <= w11620 and not w11656;
w11658 <= not w11620 and w11656;
w11659 <= not w11657 and not w11658;
w11660 <= not w11357 and not w11361;
w11661 <= a(16) and a(56);
w11662 <= a(23) and a(49);
w11663 <= not w11661 and not w11662;
w11664 <= w11661 and w11662;
w11665 <= a(32) and not w11664;
w11666 <= a(40) and w11665;
w11667 <= not w11663 and w11666;
w11668 <= not w11664 and not w11667;
w11669 <= not w11663 and w11668;
w11670 <= a(40) and not w11667;
w11671 <= a(32) and w11670;
w11672 <= not w11669 and not w11671;
w11673 <= a(21) and a(51);
w11674 <= a(22) and a(50);
w11675 <= not w11673 and not w11674;
w11676 <= w1380 and w6370;
w11677 <= w4837 and not w11676;
w11678 <= not w11675 and w11677;
w11679 <= w4837 and not w11678;
w11680 <= not w11676 and not w11678;
w11681 <= not w11675 and w11680;
w11682 <= not w11679 and not w11681;
w11683 <= not w11672 and not w11682;
w11684 <= not w11672 and not w11683;
w11685 <= not w11682 and not w11683;
w11686 <= not w11684 and not w11685;
w11687 <= a(17) and a(55);
w11688 <= w1137 and w10711;
w11689 <= w858 and w7507;
w11690 <= a(20) and a(52);
w11691 <= w11687 and w11690;
w11692 <= not w11689 and not w11691;
w11693 <= not w11688 and not w11692;
w11694 <= w11687 and not w11693;
w11695 <= not w8842 and not w11690;
w11696 <= not w11688 and not w11693;
w11697 <= not w11695 and w11696;
w11698 <= not w11694 and not w11697;
w11699 <= not w11686 and not w11698;
w11700 <= not w11686 and not w11699;
w11701 <= not w11698 and not w11699;
w11702 <= not w11700 and not w11701;
w11703 <= w529 and w9527;
w11704 <= w882 and w9715;
w11705 <= w290 and w9598;
w11706 <= not w11704 and not w11705;
w11707 <= not w11703 and not w11706;
w11708 <= not w11703 and not w11707;
w11709 <= a(10) and a(62);
w11710 <= a(11) and a(61);
w11711 <= not w11709 and not w11710;
w11712 <= w11708 and not w11711;
w11713 <= a(63) and not w11707;
w11714 <= a(9) and w11713;
w11715 <= not w11712 and not w11714;
w11716 <= not w11513 and not w11519;
w11717 <= a(24) and a(48);
w11718 <= a(25) and a(47);
w11719 <= not w11717 and not w11718;
w11720 <= w1710 and w6058;
w11721 <= a(60) and not w11720;
w11722 <= a(12) and w11721;
w11723 <= not w11719 and w11722;
w11724 <= a(60) and not w11723;
w11725 <= a(12) and w11724;
w11726 <= not w11720 and not w11723;
w11727 <= not w11719 and w11726;
w11728 <= not w11725 and not w11727;
w11729 <= not w11716 and not w11728;
w11730 <= not w11716 and not w11729;
w11731 <= not w11728 and not w11729;
w11732 <= not w11730 and not w11731;
w11733 <= not w11715 and not w11732;
w11734 <= w11715 and not w11731;
w11735 <= not w11730 and w11734;
w11736 <= not w11733 and not w11735;
w11737 <= not w11702 and w11736;
w11738 <= w11702 and not w11736;
w11739 <= not w11737 and not w11738;
w11740 <= not w11660 and w11739;
w11741 <= w11660 and not w11739;
w11742 <= not w11740 and not w11741;
w11743 <= not w11336 and not w11340;
w11744 <= w11529 and w11544;
w11745 <= not w11529 and not w11544;
w11746 <= not w11744 and not w11745;
w11747 <= w11450 and not w11746;
w11748 <= not w11450 and w11746;
w11749 <= not w11747 and not w11748;
w11750 <= not w11328 and not w11332;
w11751 <= not w11749 and w11750;
w11752 <= w11749 and not w11750;
w11753 <= not w11751 and not w11752;
w11754 <= w701 and w8242;
w11755 <= w627 and w8791;
w11756 <= w551 and w8793;
w11757 <= not w11755 and not w11756;
w11758 <= not w11754 and not w11757;
w11759 <= not w11754 and not w11758;
w11760 <= a(14) and a(58);
w11761 <= a(15) and a(57);
w11762 <= not w11760 and not w11761;
w11763 <= w11759 and not w11762;
w11764 <= a(59) and not w11758;
w11765 <= a(13) and w11764;
w11766 <= not w11763 and not w11765;
w11767 <= w2137 and w5519;
w11768 <= w2606 and w7553;
w11769 <= w2033 and w5366;
w11770 <= not w11768 and not w11769;
w11771 <= not w11767 and not w11770;
w11772 <= a(46) and not w11771;
w11773 <= a(26) and w11772;
w11774 <= not w11767 and not w11771;
w11775 <= a(27) and a(45);
w11776 <= a(28) and a(44);
w11777 <= not w11775 and not w11776;
w11778 <= w11774 and not w11777;
w11779 <= not w11773 and not w11778;
w11780 <= not w11766 and not w11779;
w11781 <= not w11766 and not w11780;
w11782 <= not w11779 and not w11780;
w11783 <= not w11781 and not w11782;
w11784 <= a(19) and a(53);
w11785 <= a(33) and a(39);
w11786 <= not w11241 and not w11785;
w11787 <= w3956 and w4889;
w11788 <= w11784 and not w11787;
w11789 <= not w11786 and w11788;
w11790 <= w11784 and not w11789;
w11791 <= not w11787 and not w11789;
w11792 <= not w11786 and w11791;
w11793 <= not w11790 and not w11792;
w11794 <= not w11783 and not w11793;
w11795 <= not w11783 and not w11794;
w11796 <= not w11793 and not w11794;
w11797 <= not w11795 and not w11796;
w11798 <= not w11753 and w11797;
w11799 <= w11753 and not w11797;
w11800 <= not w11798 and not w11799;
w11801 <= not w11743 and w11800;
w11802 <= not w11743 and not w11801;
w11803 <= w11800 and not w11801;
w11804 <= not w11802 and not w11803;
w11805 <= w11742 and not w11804;
w11806 <= w11742 and not w11805;
w11807 <= not w11804 and not w11805;
w11808 <= not w11806 and not w11807;
w11809 <= w11659 and not w11808;
w11810 <= w11659 and not w11809;
w11811 <= not w11808 and not w11809;
w11812 <= not w11810 and not w11811;
w11813 <= not w11619 and w11812;
w11814 <= w11619 and not w11812;
w11815 <= not w11813 and not w11814;
w11816 <= not w11351 and not w11569;
w11817 <= not w11815 and w11816;
w11818 <= w11815 and not w11816;
w11819 <= not w11817 and not w11818;
w11820 <= w11578 and not w11819;
w11821 <= not w11578 and not w11817;
w11822 <= not w11818 and w11821;
w11823 <= not w11820 and not w11822;
w11824 <= not w11818 and not w11821;
w11825 <= not w11618 and not w11814;
w11826 <= not w11658 and not w11809;
w11827 <= not w11801 and not w11805;
w11828 <= not w11632 and not w11654;
w11829 <= not w11752 and not w11799;
w11830 <= not w11745 and not w11748;
w11831 <= w2949 and w5219;
w11832 <= w2404 and w6259;
w11833 <= w3618 and w5150;
w11834 <= not w11832 and not w11833;
w11835 <= not w11831 and not w11834;
w11836 <= a(42) and not w11835;
w11837 <= a(31) and w11836;
w11838 <= not w11831 and not w11835;
w11839 <= a(32) and a(41);
w11840 <= a(33) and a(40);
w11841 <= not w11839 and not w11840;
w11842 <= w11838 and not w11841;
w11843 <= not w11837 and not w11842;
w11844 <= not w11830 and not w11843;
w11845 <= not w11830 and not w11844;
w11846 <= not w11843 and not w11844;
w11847 <= not w11845 and not w11846;
w11848 <= not w11637 and not w11640;
w11849 <= w11847 and w11848;
w11850 <= not w11847 and not w11848;
w11851 <= not w11849 and not w11850;
w11852 <= not w11648 and not w11651;
w11853 <= w11851 and not w11852;
w11854 <= not w11851 and w11852;
w11855 <= not w11853 and not w11854;
w11856 <= not w11829 and w11855;
w11857 <= w11829 and not w11855;
w11858 <= not w11856 and not w11857;
w11859 <= not w11828 and w11858;
w11860 <= w11828 and not w11858;
w11861 <= not w11859 and not w11860;
w11862 <= not w11827 and w11861;
w11863 <= w11827 and not w11861;
w11864 <= not w11862 and not w11863;
w11865 <= w11826 and not w11864;
w11866 <= not w11826 and w11864;
w11867 <= not w11865 and not w11866;
w11868 <= not w11610 and not w11614;
w11869 <= not w11729 and not w11733;
w11870 <= not w11643 and not w11646;
w11871 <= w11869 and w11870;
w11872 <= not w11869 and not w11870;
w11873 <= not w11871 and not w11872;
w11874 <= not w11780 and not w11794;
w11875 <= not w11873 and w11874;
w11876 <= w11873 and not w11874;
w11877 <= not w11875 and not w11876;
w11878 <= not w11737 and not w11740;
w11879 <= not w11877 and w11878;
w11880 <= w11877 and not w11878;
w11881 <= not w11879 and not w11880;
w11882 <= not w11683 and not w11699;
w11883 <= a(13) and a(60);
w11884 <= not w11680 and w11883;
w11885 <= w11680 and not w11883;
w11886 <= not w11884 and not w11885;
w11887 <= w11791 and not w11886;
w11888 <= not w11791 and w11886;
w11889 <= not w11887 and not w11888;
w11890 <= w11708 and w11726;
w11891 <= not w11708 and not w11726;
w11892 <= not w11890 and not w11891;
w11893 <= w11696 and not w11892;
w11894 <= not w11696 and w11892;
w11895 <= not w11893 and not w11894;
w11896 <= w11889 and w11895;
w11897 <= not w11889 and not w11895;
w11898 <= not w11896 and not w11897;
w11899 <= not w11882 and w11898;
w11900 <= w11882 and not w11898;
w11901 <= not w11899 and not w11900;
w11902 <= w11881 and w11901;
w11903 <= not w11881 and not w11901;
w11904 <= not w11902 and not w11903;
w11905 <= w11868 and not w11904;
w11906 <= not w11868 and w11904;
w11907 <= not w11905 and not w11906;
w11908 <= a(11) and a(62);
w11909 <= not a(37) and not w11908;
w11910 <= a(62) and w4367;
w11911 <= a(50) and not w11910;
w11912 <= a(23) and w11911;
w11913 <= not w11909 and w11912;
w11914 <= not w11910 and not w11913;
w11915 <= not w11909 and w11914;
w11916 <= a(50) and not w11913;
w11917 <= a(23) and w11916;
w11918 <= not w11915 and not w11917;
w11919 <= a(49) and a(54);
w11920 <= w1470 and w11919;
w11921 <= w955 and w7507;
w11922 <= w3997 and w9607;
w11923 <= not w11921 and not w11922;
w11924 <= not w11920 and not w11923;
w11925 <= a(55) and not w11924;
w11926 <= a(18) and w11925;
w11927 <= not w11920 and not w11924;
w11928 <= a(24) and a(49);
w11929 <= not w8845 and not w11928;
w11930 <= w11927 and not w11929;
w11931 <= not w11926 and not w11930;
w11932 <= not w11918 and not w11931;
w11933 <= not w11918 and not w11932;
w11934 <= not w11931 and not w11932;
w11935 <= not w11933 and not w11934;
w11936 <= w1300 and w7239;
w11937 <= w1499 and w7038;
w11938 <= w1380 and w6774;
w11939 <= not w11937 and not w11938;
w11940 <= not w11936 and not w11939;
w11941 <= a(51) and not w11940;
w11942 <= a(22) and w11941;
w11943 <= not w11936 and not w11940;
w11944 <= a(20) and a(53);
w11945 <= a(21) and a(52);
w11946 <= not w11944 and not w11945;
w11947 <= w11943 and not w11946;
w11948 <= not w11942 and not w11947;
w11949 <= not w11935 and not w11948;
w11950 <= not w11935 and not w11949;
w11951 <= not w11948 and not w11949;
w11952 <= not w11950 and not w11951;
w11953 <= a(15) and a(58);
w11954 <= a(16) and a(57);
w11955 <= not w11953 and not w11954;
w11956 <= w697 and w8242;
w11957 <= w699 and w8791;
w11958 <= w701 and w8793;
w11959 <= not w11957 and not w11958;
w11960 <= not w11956 and not w11959;
w11961 <= not w11956 and not w11960;
w11962 <= not w11955 and w11961;
w11963 <= a(59) and not w11960;
w11964 <= a(14) and w11963;
w11965 <= not w11962 and not w11964;
w11966 <= a(26) and a(47);
w11967 <= a(27) and a(46);
w11968 <= not w11966 and not w11967;
w11969 <= w2033 and w5472;
w11970 <= a(56) and not w11969;
w11971 <= a(17) and w11970;
w11972 <= not w11968 and w11971;
w11973 <= a(56) and not w11972;
w11974 <= a(17) and w11973;
w11975 <= not w11969 and not w11972;
w11976 <= not w11968 and w11975;
w11977 <= not w11974 and not w11976;
w11978 <= not w11668 and not w11977;
w11979 <= w11668 and w11977;
w11980 <= not w11978 and not w11979;
w11981 <= not w11965 and w11980;
w11982 <= not w11965 and not w11981;
w11983 <= w11980 and not w11981;
w11984 <= not w11982 and not w11983;
w11985 <= not w11952 and not w11984;
w11986 <= not w11952 and not w11985;
w11987 <= not w11984 and not w11985;
w11988 <= not w11986 and not w11987;
w11989 <= not w11624 and not w11628;
w11990 <= w11988 and w11989;
w11991 <= not w11988 and not w11989;
w11992 <= not w11990 and not w11991;
w11993 <= not w11602 and not w11607;
w11994 <= w11759 and w11774;
w11995 <= not w11759 and not w11774;
w11996 <= not w11994 and not w11995;
w11997 <= w11591 and not w11996;
w11998 <= not w11591 and w11996;
w11999 <= not w11997 and not w11998;
w12000 <= not w11594 and not w11600;
w12001 <= not w11999 and w12000;
w12002 <= w11999 and not w12000;
w12003 <= not w12001 and not w12002;
w12004 <= a(10) and a(63);
w12005 <= a(12) and a(61);
w12006 <= not w12004 and not w12005;
w12007 <= w286 and w9715;
w12008 <= a(48) and not w12007;
w12009 <= a(25) and w12008;
w12010 <= not w12006 and w12009;
w12011 <= not w12007 and not w12010;
w12012 <= not w12006 and w12011;
w12013 <= a(48) and not w12010;
w12014 <= a(25) and w12013;
w12015 <= not w12012 and not w12014;
w12016 <= w2423 and w5102;
w12017 <= w2916 and w4617;
w12018 <= w2140 and w5519;
w12019 <= not w12017 and not w12018;
w12020 <= not w12016 and not w12019;
w12021 <= a(45) and not w12020;
w12022 <= a(28) and w12021;
w12023 <= not w12016 and not w12020;
w12024 <= a(29) and a(44);
w12025 <= a(30) and a(43);
w12026 <= not w12024 and not w12025;
w12027 <= w12023 and not w12026;
w12028 <= not w12022 and not w12027;
w12029 <= not w12015 and not w12028;
w12030 <= not w12015 and not w12029;
w12031 <= not w12028 and not w12029;
w12032 <= not w12030 and not w12031;
w12033 <= w3634 and w4371;
w12034 <= w3493 and w4554;
w12035 <= w3125 and w4889;
w12036 <= not w12034 and not w12035;
w12037 <= not w12033 and not w12036;
w12038 <= w4554 and not w12037;
w12039 <= not w12033 and not w12037;
w12040 <= a(35) and a(38);
w12041 <= not w3493 and not w12040;
w12042 <= w12039 and not w12041;
w12043 <= not w12038 and not w12042;
w12044 <= not w12032 and not w12043;
w12045 <= not w12032 and not w12044;
w12046 <= not w12043 and not w12044;
w12047 <= not w12045 and not w12046;
w12048 <= not w12003 and w12047;
w12049 <= w12003 and not w12047;
w12050 <= not w12048 and not w12049;
w12051 <= not w11993 and w12050;
w12052 <= not w11993 and not w12051;
w12053 <= w12050 and not w12051;
w12054 <= not w12052 and not w12053;
w12055 <= w11992 and not w12054;
w12056 <= w11992 and not w12055;
w12057 <= not w12054 and not w12055;
w12058 <= not w12056 and not w12057;
w12059 <= w11907 and not w12058;
w12060 <= w11907 and not w12059;
w12061 <= not w12058 and not w12059;
w12062 <= not w12060 and not w12061;
w12063 <= not w11867 and w12062;
w12064 <= w11867 and not w12062;
w12065 <= not w12063 and not w12064;
w12066 <= w11825 and not w12065;
w12067 <= not w11825 and w12065;
w12068 <= not w12066 and not w12067;
w12069 <= not w11824 and not w12068;
w12070 <= w11824 and w12068;
w12071 <= not w12069 and not w12070;
w12072 <= not w11866 and not w12064;
w12073 <= not w11859 and not w11862;
w12074 <= w11838 and w12039;
w12075 <= not w11838 and not w12039;
w12076 <= not w12074 and not w12075;
w12077 <= w697 and w8793;
w12078 <= w699 and w9895;
w12079 <= w701 and w9315;
w12080 <= not w12078 and not w12079;
w12081 <= not w12077 and not w12080;
w12082 <= a(60) and not w12081;
w12083 <= a(14) and w12082;
w12084 <= a(15) and a(59);
w12085 <= a(16) and a(58);
w12086 <= not w12084 and not w12085;
w12087 <= not w12077 and not w12081;
w12088 <= not w12086 and w12087;
w12089 <= not w12083 and not w12088;
w12090 <= w12076 and not w12089;
w12091 <= w12076 and not w12090;
w12092 <= not w12089 and not w12090;
w12093 <= not w12091 and not w12092;
w12094 <= not w11932 and not w11949;
w12095 <= w12093 and w12094;
w12096 <= not w12093 and not w12094;
w12097 <= not w12095 and not w12096;
w12098 <= not w11844 and not w11850;
w12099 <= not w12097 and w12098;
w12100 <= w12097 and not w12098;
w12101 <= not w12099 and not w12100;
w12102 <= not w11985 and not w11991;
w12103 <= not w12002 and not w12049;
w12104 <= not w12102 and not w12103;
w12105 <= not w12102 and not w12104;
w12106 <= not w12103 and not w12104;
w12107 <= not w12105 and not w12106;
w12108 <= w12101 and not w12107;
w12109 <= not w12101 and w12107;
w12110 <= not w12073 and not w12109;
w12111 <= not w12108 and w12110;
w12112 <= not w12073 and not w12111;
w12113 <= not w12109 and not w12111;
w12114 <= not w12108 and w12113;
w12115 <= not w12112 and not w12114;
w12116 <= w554 and w9527;
w12117 <= a(61) and not w12116;
w12118 <= a(13) and w12117;
w12119 <= a(62) and not w12116;
w12120 <= a(12) and w12119;
w12121 <= not w12118 and not w12120;
w12122 <= not w11914 and not w12121;
w12123 <= not w11914 and not w12122;
w12124 <= not w12121 and not w12122;
w12125 <= not w12123 and not w12124;
w12126 <= a(30) and a(44);
w12127 <= w9424 and w12126;
w12128 <= w2423 and w5519;
w12129 <= a(29) and a(57);
w12130 <= w8925 and w12129;
w12131 <= not w12128 and not w12130;
w12132 <= not w12127 and not w12131;
w12133 <= a(45) and not w12132;
w12134 <= a(29) and w12133;
w12135 <= not w12127 and not w12132;
w12136 <= not w9424 and not w12126;
w12137 <= w12135 and not w12136;
w12138 <= not w12134 and not w12137;
w12139 <= not w12125 and not w12138;
w12140 <= not w12125 and not w12139;
w12141 <= not w12138 and not w12139;
w12142 <= not w12140 and not w12141;
w12143 <= not w11995 and not w11998;
w12144 <= w12142 and w12143;
w12145 <= not w12142 and not w12143;
w12146 <= not w12144 and not w12145;
w12147 <= a(31) and a(43);
w12148 <= a(32) and a(42);
w12149 <= not w12147 and not w12148;
w12150 <= w3618 and w4824;
w12151 <= a(63) and not w12150;
w12152 <= not w12149 and w12151;
w12153 <= a(11) and w12152;
w12154 <= not w12150 and not w12153;
w12155 <= not w12149 and w12154;
w12156 <= a(63) and not w12153;
w12157 <= a(11) and w12156;
w12158 <= not w12155 and not w12157;
w12159 <= a(18) and a(56);
w12160 <= a(25) and a(49);
w12161 <= not w12159 and not w12160;
w12162 <= a(25) and a(56);
w12163 <= w10296 and w12162;
w12164 <= w5148 and not w12163;
w12165 <= not w12161 and w12164;
w12166 <= w5148 and not w12165;
w12167 <= not w12163 and not w12165;
w12168 <= not w12161 and w12167;
w12169 <= not w12166 and not w12168;
w12170 <= not w12158 and not w12169;
w12171 <= not w12158 and not w12170;
w12172 <= not w12169 and not w12170;
w12173 <= not w12171 and not w12172;
w12174 <= w2137 and w5472;
w12175 <= w2606 and w8384;
w12176 <= w2033 and w6058;
w12177 <= not w12175 and not w12176;
w12178 <= not w12174 and not w12177;
w12179 <= a(48) and not w12178;
w12180 <= a(26) and w12179;
w12181 <= not w12174 and not w12178;
w12182 <= a(27) and a(47);
w12183 <= a(28) and a(46);
w12184 <= not w12182 and not w12183;
w12185 <= w12181 and not w12184;
w12186 <= not w12180 and not w12185;
w12187 <= not w12173 and not w12186;
w12188 <= not w12173 and not w12187;
w12189 <= not w12186 and not w12187;
w12190 <= not w12188 and not w12189;
w12191 <= a(21) and a(53);
w12192 <= not w8018 and not w12191;
w12193 <= w1298 and w7503;
w12194 <= a(52) and a(55);
w12195 <= w3842 and w12194;
w12196 <= w1380 and w7239;
w12197 <= not w12195 and not w12196;
w12198 <= not w12193 and not w12197;
w12199 <= not w12193 and not w12198;
w12200 <= not w12192 and w12199;
w12201 <= a(52) and not w12198;
w12202 <= a(22) and w12201;
w12203 <= not w12200 and not w12202;
w12204 <= a(35) and a(39);
w12205 <= not w5001 and not w12204;
w12206 <= w3125 and w3977;
w12207 <= w10849 and not w12206;
w12208 <= not w12205 and w12207;
w12209 <= w10849 and not w12208;
w12210 <= not w12206 and not w12208;
w12211 <= not w12205 and w12210;
w12212 <= not w12209 and not w12211;
w12213 <= not w12203 and not w12212;
w12214 <= not w12203 and not w12213;
w12215 <= not w12212 and not w12213;
w12216 <= not w12214 and not w12215;
w12217 <= a(23) and a(51);
w12218 <= a(24) and a(50);
w12219 <= not w12217 and not w12218;
w12220 <= w1472 and w6370;
w12221 <= w3336 and not w12220;
w12222 <= not w12219 and w12221;
w12223 <= w3336 and not w12222;
w12224 <= not w12220 and not w12222;
w12225 <= not w12219 and w12224;
w12226 <= not w12223 and not w12225;
w12227 <= not w12216 and not w12226;
w12228 <= not w12216 and not w12227;
w12229 <= not w12226 and not w12227;
w12230 <= not w12228 and not w12229;
w12231 <= not w12190 and w12230;
w12232 <= w12190 and not w12230;
w12233 <= not w12231 and not w12232;
w12234 <= w12146 and not w12233;
w12235 <= w12146 and not w12234;
w12236 <= not w12233 and not w12234;
w12237 <= not w12235 and not w12236;
w12238 <= not w11853 and not w11856;
w12239 <= w11975 and w12023;
w12240 <= not w11975 and not w12023;
w12241 <= not w12239 and not w12240;
w12242 <= w11961 and not w12241;
w12243 <= not w11961 and w12241;
w12244 <= not w12242 and not w12243;
w12245 <= w11927 and w11943;
w12246 <= not w11927 and not w11943;
w12247 <= not w12245 and not w12246;
w12248 <= w12011 and not w12247;
w12249 <= not w12011 and w12247;
w12250 <= not w12248 and not w12249;
w12251 <= not w12029 and not w12044;
w12252 <= not w12250 and w12251;
w12253 <= w12250 and not w12251;
w12254 <= not w12252 and not w12253;
w12255 <= w12244 and w12254;
w12256 <= not w12244 and not w12254;
w12257 <= not w12255 and not w12256;
w12258 <= not w12238 and w12257;
w12259 <= w12238 and not w12257;
w12260 <= not w12258 and not w12259;
w12261 <= not w12237 and w12260;
w12262 <= w12260 and not w12261;
w12263 <= not w12237 and not w12261;
w12264 <= not w12262 and not w12263;
w12265 <= not w12115 and w12264;
w12266 <= w12115 and not w12264;
w12267 <= not w12265 and not w12266;
w12268 <= not w11906 and not w12059;
w12269 <= not w12051 and not w12055;
w12270 <= not w11880 and not w11902;
w12271 <= not w11891 and not w11894;
w12272 <= not w11884 and not w11888;
w12273 <= w12271 and w12272;
w12274 <= not w12271 and not w12272;
w12275 <= not w12273 and not w12274;
w12276 <= not w11978 and not w11981;
w12277 <= not w12275 and w12276;
w12278 <= w12275 and not w12276;
w12279 <= not w12277 and not w12278;
w12280 <= not w11896 and not w11899;
w12281 <= not w11872 and not w11876;
w12282 <= w12280 and w12281;
w12283 <= not w12280 and not w12281;
w12284 <= not w12282 and not w12283;
w12285 <= w12279 and w12284;
w12286 <= not w12279 and not w12284;
w12287 <= not w12285 and not w12286;
w12288 <= not w12270 and w12287;
w12289 <= w12270 and not w12287;
w12290 <= not w12288 and not w12289;
w12291 <= not w12269 and w12290;
w12292 <= w12269 and not w12290;
w12293 <= not w12291 and not w12292;
w12294 <= not w12268 and w12293;
w12295 <= w12268 and not w12293;
w12296 <= not w12294 and not w12295;
w12297 <= not w12267 and w12296;
w12298 <= w12267 and not w12296;
w12299 <= not w12297 and not w12298;
w12300 <= w12072 and not w12299;
w12301 <= not w12072 and w12299;
w12302 <= not w12300 and not w12301;
w12303 <= not w11824 and not w12066;
w12304 <= not w12067 and not w12303;
w12305 <= not w12302 and w12304;
w12306 <= w12302 and not w12304;
w12307 <= not w12305 and not w12306;
w12308 <= not w12294 and not w12297;
w12309 <= not w12288 and not w12291;
w12310 <= not w12075 and not w12090;
w12311 <= not w12246 and not w12249;
w12312 <= w12310 and w12311;
w12313 <= not w12310 and not w12311;
w12314 <= not w12312 and not w12313;
w12315 <= not w12240 and not w12243;
w12316 <= not w12314 and w12315;
w12317 <= w12314 and not w12315;
w12318 <= not w12316 and not w12317;
w12319 <= not w12190 and not w12230;
w12320 <= not w12234 and not w12319;
w12321 <= w12318 and not w12320;
w12322 <= not w12318 and w12320;
w12323 <= not w12321 and not w12322;
w12324 <= not w12139 and not w12145;
w12325 <= w12210 and w12224;
w12326 <= not w12210 and not w12224;
w12327 <= not w12325 and not w12326;
w12328 <= w12199 and not w12327;
w12329 <= not w12199 and w12327;
w12330 <= not w12328 and not w12329;
w12331 <= w12154 and w12167;
w12332 <= not w12154 and not w12167;
w12333 <= not w12331 and not w12332;
w12334 <= not w12116 and not w12122;
w12335 <= not w12333 and w12334;
w12336 <= w12333 and not w12334;
w12337 <= not w12335 and not w12336;
w12338 <= w12330 and w12337;
w12339 <= not w12330 and not w12337;
w12340 <= not w12338 and not w12339;
w12341 <= not w12324 and w12340;
w12342 <= w12324 and not w12340;
w12343 <= not w12341 and not w12342;
w12344 <= w12323 and w12343;
w12345 <= not w12323 and not w12343;
w12346 <= not w12344 and not w12345;
w12347 <= w12309 and not w12346;
w12348 <= not w12309 and w12346;
w12349 <= not w12347 and not w12348;
w12350 <= a(12) and a(63);
w12351 <= a(19) and a(56);
w12352 <= not w12350 and not w12351;
w12353 <= a(19) and a(63);
w12354 <= w10691 and w12353;
w12355 <= a(45) and not w12354;
w12356 <= a(30) and w12355;
w12357 <= not w12352 and w12356;
w12358 <= not w12354 and not w12357;
w12359 <= not w12352 and w12358;
w12360 <= a(45) and not w12357;
w12361 <= a(30) and w12360;
w12362 <= not w12359 and not w12361;
w12363 <= a(23) and a(52);
w12364 <= a(35) and a(40);
w12365 <= not w8742 and not w12364;
w12366 <= w3634 and w3977;
w12367 <= w12363 and not w12366;
w12368 <= not w12365 and w12367;
w12369 <= w12363 and not w12368;
w12370 <= not w12366 and not w12368;
w12371 <= not w12365 and w12370;
w12372 <= not w12369 and not w12371;
w12373 <= not w12362 and not w12372;
w12374 <= not w12362 and not w12373;
w12375 <= not w12372 and not w12373;
w12376 <= not w12374 and not w12375;
w12377 <= a(38) and a(62);
w12378 <= a(13) and w12377;
w12379 <= w4371 and not w12378;
w12380 <= w4371 and not w12379;
w12381 <= not w12378 and not w12379;
w12382 <= a(13) and a(62);
w12383 <= not a(38) and not w12382;
w12384 <= w12381 and not w12383;
w12385 <= not w12380 and not w12384;
w12386 <= not w12376 and not w12385;
w12387 <= not w12376 and not w12386;
w12388 <= not w12385 and not w12386;
w12389 <= not w12387 and not w12388;
w12390 <= not w12274 and not w12278;
w12391 <= w12389 and w12390;
w12392 <= not w12389 and not w12390;
w12393 <= not w12391 and not w12392;
w12394 <= w697 and w9315;
w12395 <= w699 and w8711;
w12396 <= w701 and w9318;
w12397 <= not w12395 and not w12396;
w12398 <= not w12394 and not w12397;
w12399 <= not w12394 and not w12398;
w12400 <= a(15) and a(60);
w12401 <= a(16) and a(59);
w12402 <= not w12400 and not w12401;
w12403 <= w12399 and not w12402;
w12404 <= a(61) and not w12398;
w12405 <= a(14) and w12404;
w12406 <= not w12403 and not w12405;
w12407 <= a(49) and a(57);
w12408 <= w4349 and w12407;
w12409 <= a(26) and a(58);
w12410 <= w6869 and w12409;
w12411 <= w858 and w8242;
w12412 <= not w12410 and not w12411;
w12413 <= not w12408 and not w12412;
w12414 <= a(58) and not w12413;
w12415 <= a(17) and w12414;
w12416 <= not w12408 and not w12413;
w12417 <= a(18) and a(57);
w12418 <= a(26) and a(49);
w12419 <= not w12417 and not w12418;
w12420 <= w12416 and not w12419;
w12421 <= not w12415 and not w12420;
w12422 <= not w12406 and not w12421;
w12423 <= not w12406 and not w12422;
w12424 <= not w12421 and not w12422;
w12425 <= not w12423 and not w12424;
w12426 <= w2140 and w5472;
w12427 <= w1847 and w8384;
w12428 <= w2137 and w6058;
w12429 <= not w12427 and not w12428;
w12430 <= not w12426 and not w12429;
w12431 <= a(48) and not w12430;
w12432 <= a(27) and w12431;
w12433 <= not w12426 and not w12430;
w12434 <= a(28) and a(47);
w12435 <= a(29) and a(46);
w12436 <= not w12434 and not w12435;
w12437 <= w12433 and not w12436;
w12438 <= not w12432 and not w12437;
w12439 <= not w12425 and not w12438;
w12440 <= not w12425 and not w12439;
w12441 <= not w12438 and not w12439;
w12442 <= not w12440 and not w12441;
w12443 <= w12393 and not w12442;
w12444 <= not w12393 and w12442;
w12445 <= not w12283 and not w12285;
w12446 <= w12135 and w12181;
w12447 <= not w12135 and not w12181;
w12448 <= not w12446 and not w12447;
w12449 <= w12087 and not w12448;
w12450 <= not w12087 and w12448;
w12451 <= not w12449 and not w12450;
w12452 <= not w12213 and not w12227;
w12453 <= not w12170 and not w12187;
w12454 <= w12452 and w12453;
w12455 <= not w12452 and not w12453;
w12456 <= not w12454 and not w12455;
w12457 <= w12451 and w12456;
w12458 <= not w12451 and not w12456;
w12459 <= not w12457 and not w12458;
w12460 <= not w12445 and w12459;
w12461 <= w12445 and not w12459;
w12462 <= not w12460 and not w12461;
w12463 <= not w12444 and w12462;
w12464 <= not w12443 and w12463;
w12465 <= w12462 and not w12464;
w12466 <= not w12444 and not w12464;
w12467 <= not w12443 and w12466;
w12468 <= not w12465 and not w12467;
w12469 <= not w12349 and w12468;
w12470 <= w12349 and not w12468;
w12471 <= not w12469 and not w12470;
w12472 <= not w12096 and not w12100;
w12473 <= a(20) and a(55);
w12474 <= a(25) and a(50);
w12475 <= not w12473 and not w12474;
w12476 <= w12473 and w12474;
w12477 <= a(34) and not w12476;
w12478 <= a(41) and w12477;
w12479 <= not w12475 and w12478;
w12480 <= not w12476 and not w12479;
w12481 <= not w12475 and w12480;
w12482 <= a(41) and not w12479;
w12483 <= a(34) and w12482;
w12484 <= not w12481 and not w12483;
w12485 <= w2949 and w4824;
w12486 <= w2404 and w4445;
w12487 <= w3618 and w5102;
w12488 <= not w12486 and not w12487;
w12489 <= not w12485 and not w12488;
w12490 <= a(44) and not w12489;
w12491 <= a(31) and w12490;
w12492 <= a(33) and a(42);
w12493 <= not w5100 and not w12492;
w12494 <= not w12485 and not w12489;
w12495 <= not w12493 and w12494;
w12496 <= not w12491 and not w12495;
w12497 <= not w12484 and not w12496;
w12498 <= not w12484 and not w12497;
w12499 <= not w12496 and not w12497;
w12500 <= not w12498 and not w12499;
w12501 <= w1921 and w7038;
w12502 <= w1380 and w7505;
w12503 <= a(24) and a(54);
w12504 <= w11673 and w12503;
w12505 <= not w12502 and not w12504;
w12506 <= not w12501 and not w12505;
w12507 <= a(54) and not w12506;
w12508 <= a(21) and w12507;
w12509 <= not w12501 and not w12506;
w12510 <= a(22) and a(53);
w12511 <= a(24) and a(51);
w12512 <= not w12510 and not w12511;
w12513 <= w12509 and not w12512;
w12514 <= not w12508 and not w12513;
w12515 <= not w12500 and not w12514;
w12516 <= not w12500 and not w12515;
w12517 <= not w12514 and not w12515;
w12518 <= not w12516 and not w12517;
w12519 <= not w12253 and not w12255;
w12520 <= not w12518 and not w12519;
w12521 <= not w12518 and not w12520;
w12522 <= not w12519 and not w12520;
w12523 <= not w12521 and not w12522;
w12524 <= not w12472 and not w12523;
w12525 <= not w12472 and not w12524;
w12526 <= not w12523 and not w12524;
w12527 <= not w12525 and not w12526;
w12528 <= not w12104 and not w12108;
w12529 <= not w12527 and not w12528;
w12530 <= not w12527 and not w12529;
w12531 <= not w12528 and not w12529;
w12532 <= not w12530 and not w12531;
w12533 <= not w12258 and not w12261;
w12534 <= w12532 and w12533;
w12535 <= not w12532 and not w12533;
w12536 <= not w12534 and not w12535;
w12537 <= not w12115 and not w12264;
w12538 <= not w12111 and not w12537;
w12539 <= w12536 and not w12538;
w12540 <= not w12536 and w12538;
w12541 <= not w12539 and not w12540;
w12542 <= w12471 and w12541;
w12543 <= not w12471 and not w12541;
w12544 <= not w12542 and not w12543;
w12545 <= not w12308 and w12544;
w12546 <= w12308 and not w12544;
w12547 <= not w12545 and not w12546;
w12548 <= not w12300 and not w12304;
w12549 <= not w12301 and not w12548;
w12550 <= not w12547 and w12549;
w12551 <= w12547 and not w12549;
w12552 <= not w12550 and not w12551;
w12553 <= not w12546 and not w12549;
w12554 <= not w12545 and not w12553;
w12555 <= not w12539 and not w12542;
w12556 <= not w12332 and not w12336;
w12557 <= not w12447 and not w12450;
w12558 <= w12556 and w12557;
w12559 <= not w12556 and not w12557;
w12560 <= not w12558 and not w12559;
w12561 <= not w12326 and not w12329;
w12562 <= not w12560 and w12561;
w12563 <= w12560 and not w12561;
w12564 <= not w12562 and not w12563;
w12565 <= not w12392 and not w12443;
w12566 <= w12564 and not w12565;
w12567 <= not w12564 and w12565;
w12568 <= not w12566 and not w12567;
w12569 <= w12433 and w12480;
w12570 <= not w12433 and not w12480;
w12571 <= not w12569 and not w12570;
w12572 <= w12358 and not w12571;
w12573 <= not w12358 and w12571;
w12574 <= not w12572 and not w12573;
w12575 <= not w12497 and not w12515;
w12576 <= a(14) and a(62);
w12577 <= w12381 and not w12576;
w12578 <= not w12381 and w12576;
w12579 <= not w12370 and not w12578;
w12580 <= not w12577 and w12579;
w12581 <= not w12578 and not w12580;
w12582 <= not w12577 and w12581;
w12583 <= not w12370 and not w12580;
w12584 <= not w12582 and not w12583;
w12585 <= not w12575 and not w12584;
w12586 <= not w12575 and not w12585;
w12587 <= not w12584 and not w12585;
w12588 <= not w12586 and not w12587;
w12589 <= w12574 and not w12588;
w12590 <= w12574 and not w12589;
w12591 <= not w12588 and not w12589;
w12592 <= not w12590 and not w12591;
w12593 <= w12568 and not w12592;
w12594 <= w12568 and not w12593;
w12595 <= not w12592 and not w12593;
w12596 <= not w12594 and not w12595;
w12597 <= not w12529 and not w12535;
w12598 <= w12596 and w12597;
w12599 <= not w12596 and not w12597;
w12600 <= not w12598 and not w12599;
w12601 <= not w12520 and not w12524;
w12602 <= w12399 and w12416;
w12603 <= not w12399 and not w12416;
w12604 <= not w12602 and not w12603;
w12605 <= w12494 and not w12604;
w12606 <= not w12494 and w12604;
w12607 <= not w12605 and not w12606;
w12608 <= not w12422 and not w12439;
w12609 <= not w12373 and not w12386;
w12610 <= w12608 and w12609;
w12611 <= not w12608 and not w12609;
w12612 <= not w12610 and not w12611;
w12613 <= w12607 and w12612;
w12614 <= not w12607 and not w12612;
w12615 <= not w12613 and not w12614;
w12616 <= w12601 and not w12615;
w12617 <= not w12601 and w12615;
w12618 <= not w12616 and not w12617;
w12619 <= w2423 and w5472;
w12620 <= w2916 and w8384;
w12621 <= w2140 and w6058;
w12622 <= not w12620 and not w12621;
w12623 <= not w12619 and not w12622;
w12624 <= not w12619 and not w12623;
w12625 <= a(29) and a(47);
w12626 <= a(30) and a(46);
w12627 <= not w12625 and not w12626;
w12628 <= w12624 and not w12627;
w12629 <= a(48) and not w12623;
w12630 <= a(28) and w12629;
w12631 <= not w12628 and not w12630;
w12632 <= w3634 and w5219;
w12633 <= w4401 and w6259;
w12634 <= w3125 and w5150;
w12635 <= not w12633 and not w12634;
w12636 <= not w12632 and not w12635;
w12637 <= a(42) and not w12636;
w12638 <= a(34) and w12637;
w12639 <= not w12632 and not w12636;
w12640 <= a(35) and a(41);
w12641 <= a(36) and a(40);
w12642 <= not w12640 and not w12641;
w12643 <= w12639 and not w12642;
w12644 <= not w12638 and not w12643;
w12645 <= not w12631 and not w12644;
w12646 <= not w12631 and not w12645;
w12647 <= not w12644 and not w12645;
w12648 <= not w12646 and not w12647;
w12649 <= a(24) and a(52);
w12650 <= a(25) and a(51);
w12651 <= not w12649 and not w12650;
w12652 <= w1710 and w6774;
w12653 <= w5236 and not w12652;
w12654 <= not w12651 and w12653;
w12655 <= w5236 and not w12654;
w12656 <= not w12652 and not w12654;
w12657 <= not w12651 and w12656;
w12658 <= not w12655 and not w12657;
w12659 <= not w12648 and not w12658;
w12660 <= not w12648 and not w12659;
w12661 <= not w12658 and not w12659;
w12662 <= not w12660 and not w12661;
w12663 <= not w12313 and not w12317;
w12664 <= w12662 and w12663;
w12665 <= not w12662 and not w12663;
w12666 <= not w12664 and not w12665;
w12667 <= w854 and w9315;
w12668 <= w799 and w8711;
w12669 <= w697 and w9318;
w12670 <= not w12668 and not w12669;
w12671 <= not w12667 and not w12670;
w12672 <= a(61) and not w12671;
w12673 <= a(15) and w12672;
w12674 <= not w12667 and not w12671;
w12675 <= a(16) and a(60);
w12676 <= a(17) and a(59);
w12677 <= not w12675 and not w12676;
w12678 <= w12674 and not w12677;
w12679 <= not w12673 and not w12678;
w12680 <= w12509 and not w12679;
w12681 <= not w12509 and w12679;
w12682 <= not w12680 and not w12681;
w12683 <= a(26) and a(50);
w12684 <= a(27) and a(49);
w12685 <= not w12683 and not w12684;
w12686 <= w2033 and w6131;
w12687 <= a(58) and not w12686;
w12688 <= a(18) and w12687;
w12689 <= not w12685 and w12688;
w12690 <= a(58) and not w12689;
w12691 <= a(18) and w12690;
w12692 <= not w12686 and not w12689;
w12693 <= not w12685 and w12692;
w12694 <= not w12691 and not w12693;
w12695 <= not w12682 and not w12694;
w12696 <= w12682 and w12694;
w12697 <= not w12695 and not w12696;
w12698 <= w12666 and w12697;
w12699 <= not w12666 and not w12697;
w12700 <= w12618 and not w12699;
w12701 <= not w12698 and w12700;
w12702 <= w12618 and not w12701;
w12703 <= not w12699 and not w12701;
w12704 <= not w12698 and w12703;
w12705 <= not w12702 and not w12704;
w12706 <= w12600 and not w12705;
w12707 <= not w12600 and w12705;
w12708 <= not w12348 and not w12470;
w12709 <= not w12460 and not w12464;
w12710 <= not w12321 and not w12344;
w12711 <= not w12338 and not w12341;
w12712 <= a(31) and a(45);
w12713 <= a(32) and a(44);
w12714 <= not w12712 and not w12713;
w12715 <= w3618 and w5519;
w12716 <= a(63) and not w12715;
w12717 <= not w12714 and w12716;
w12718 <= a(13) and w12717;
w12719 <= not w12715 and not w12718;
w12720 <= not w12714 and w12719;
w12721 <= a(63) and not w12718;
w12722 <= a(13) and w12721;
w12723 <= not w12720 and not w12722;
w12724 <= a(19) and a(57);
w12725 <= a(23) and a(53);
w12726 <= not w12724 and not w12725;
w12727 <= w12724 and w12725;
w12728 <= w5255 and not w12727;
w12729 <= not w12726 and w12728;
w12730 <= w5255 and not w12729;
w12731 <= not w12727 and not w12729;
w12732 <= not w12726 and w12731;
w12733 <= not w12730 and not w12732;
w12734 <= not w12723 and not w12733;
w12735 <= not w12723 and not w12734;
w12736 <= not w12733 and not w12734;
w12737 <= not w12735 and not w12736;
w12738 <= w1380 and w7507;
w12739 <= w1499 and w7227;
w12740 <= w1300 and w8967;
w12741 <= not w12739 and not w12740;
w12742 <= not w12738 and not w12741;
w12743 <= w9791 and not w12742;
w12744 <= not w12738 and not w12742;
w12745 <= a(21) and a(55);
w12746 <= a(22) and a(54);
w12747 <= not w12745 and not w12746;
w12748 <= w12744 and not w12747;
w12749 <= not w12743 and not w12748;
w12750 <= not w12737 and not w12749;
w12751 <= not w12737 and not w12750;
w12752 <= not w12749 and not w12750;
w12753 <= not w12751 and not w12752;
w12754 <= not w12455 and not w12457;
w12755 <= not w12753 and not w12754;
w12756 <= w12753 and w12754;
w12757 <= not w12755 and not w12756;
w12758 <= not w12711 and w12757;
w12759 <= w12711 and not w12757;
w12760 <= not w12758 and not w12759;
w12761 <= not w12710 and w12760;
w12762 <= w12710 and not w12760;
w12763 <= not w12761 and not w12762;
w12764 <= not w12709 and w12763;
w12765 <= w12709 and not w12763;
w12766 <= not w12764 and not w12765;
w12767 <= not w12708 and w12766;
w12768 <= w12708 and not w12766;
w12769 <= not w12767 and not w12768;
w12770 <= not w12707 and w12769;
w12771 <= not w12706 and w12770;
w12772 <= w12769 and not w12771;
w12773 <= not w12707 and not w12771;
w12774 <= not w12706 and w12773;
w12775 <= not w12772 and not w12774;
w12776 <= not w12555 and not w12775;
w12777 <= w12555 and w12775;
w12778 <= not w12776 and not w12777;
w12779 <= not w12554 and w12778;
w12780 <= w12554 and not w12778;
w12781 <= not w12779 and not w12780;
w12782 <= not w12767 and not w12771;
w12783 <= not w12761 and not w12764;
w12784 <= w858 and w9315;
w12785 <= a(59) and not w12784;
w12786 <= a(18) and w12785;
w12787 <= a(60) and not w12784;
w12788 <= a(17) and w12787;
w12789 <= not w12786 and not w12788;
w12790 <= not w12656 and not w12789;
w12791 <= not w12656 and not w12790;
w12792 <= not w12789 and not w12790;
w12793 <= not w12791 and not w12792;
w12794 <= not w12603 and not w12606;
w12795 <= w12793 and w12794;
w12796 <= not w12793 and not w12794;
w12797 <= not w12795 and not w12796;
w12798 <= not w12570 and not w12573;
w12799 <= not w12797 and w12798;
w12800 <= w12797 and not w12798;
w12801 <= not w12799 and not w12800;
w12802 <= not w12665 and not w12698;
w12803 <= w12801 and not w12802;
w12804 <= not w12801 and w12802;
w12805 <= not w12803 and not w12804;
w12806 <= w12624 and w12744;
w12807 <= not w12624 and not w12744;
w12808 <= not w12806 and not w12807;
w12809 <= w12719 and not w12808;
w12810 <= not w12719 and w12808;
w12811 <= not w12809 and not w12810;
w12812 <= w12674 and w12692;
w12813 <= not w12674 and not w12692;
w12814 <= not w12812 and not w12813;
w12815 <= w12731 and not w12814;
w12816 <= not w12731 and w12814;
w12817 <= not w12815 and not w12816;
w12818 <= not w12734 and not w12750;
w12819 <= not w12817 and w12818;
w12820 <= w12817 and not w12818;
w12821 <= not w12819 and not w12820;
w12822 <= w12811 and w12821;
w12823 <= not w12811 and not w12821;
w12824 <= not w12822 and not w12823;
w12825 <= w12805 and w12824;
w12826 <= not w12805 and not w12824;
w12827 <= not w12825 and not w12826;
w12828 <= w12783 and not w12827;
w12829 <= not w12783 and w12827;
w12830 <= not w12828 and not w12829;
w12831 <= not w12509 and not w12679;
w12832 <= not w12695 and not w12831;
w12833 <= w12581 and w12832;
w12834 <= not w12581 and not w12832;
w12835 <= not w12833 and not w12834;
w12836 <= not w12645 and not w12659;
w12837 <= not w12835 and w12836;
w12838 <= w12835 and not w12836;
w12839 <= not w12837 and not w12838;
w12840 <= not w12755 and not w12758;
w12841 <= not w12839 and w12840;
w12842 <= w12839 and not w12840;
w12843 <= not w12841 and not w12842;
w12844 <= a(31) and a(63);
w12845 <= w7206 and w12844;
w12846 <= w2671 and w5472;
w12847 <= a(14) and a(63);
w12848 <= a(30) and a(47);
w12849 <= w12847 and w12848;
w12850 <= not w12846 and not w12849;
w12851 <= not w12845 and not w12850;
w12852 <= not w12845 and not w12851;
w12853 <= a(31) and a(46);
w12854 <= not w12847 and not w12853;
w12855 <= w12852 and not w12854;
w12856 <= w12848 and not w12851;
w12857 <= not w12855 and not w12856;
w12858 <= a(35) and a(42);
w12859 <= w3493 and w5219;
w12860 <= w4837 and w6259;
w12861 <= w3634 and w5150;
w12862 <= not w12860 and not w12861;
w12863 <= not w12859 and not w12862;
w12864 <= w12858 and not w12863;
w12865 <= not w12859 and not w12863;
w12866 <= a(36) and a(41);
w12867 <= not w5501 and not w12866;
w12868 <= w12865 and not w12867;
w12869 <= not w12864 and not w12868;
w12870 <= not w12857 and not w12869;
w12871 <= not w12857 and not w12870;
w12872 <= not w12869 and not w12870;
w12873 <= not w12871 and not w12872;
w12874 <= a(62) and w6787;
w12875 <= w4889 and not w12874;
w12876 <= w4889 and not w12875;
w12877 <= not w12874 and not w12875;
w12878 <= a(15) and a(62);
w12879 <= not a(39) and not w12878;
w12880 <= w12877 and not w12879;
w12881 <= not w12876 and not w12880;
w12882 <= not w12873 and not w12881;
w12883 <= not w12873 and not w12882;
w12884 <= not w12881 and not w12882;
w12885 <= not w12883 and not w12884;
w12886 <= not w12559 and not w12563;
w12887 <= w12885 and w12886;
w12888 <= not w12885 and not w12886;
w12889 <= not w12887 and not w12888;
w12890 <= w1300 and w8006;
w12891 <= w1298 and w7748;
w12892 <= w1296 and w8242;
w12893 <= not w12891 and not w12892;
w12894 <= not w12890 and not w12893;
w12895 <= a(58) and not w12894;
w12896 <= a(19) and w12895;
w12897 <= not w12890 and not w12894;
w12898 <= a(21) and a(56);
w12899 <= not w10464 and not w12898;
w12900 <= w12897 and not w12899;
w12901 <= not w12896 and not w12900;
w12902 <= w12639 and not w12901;
w12903 <= not w12639 and w12901;
w12904 <= not w12902 and not w12903;
w12905 <= w2140 and w6062;
w12906 <= w1847 and w5694;
w12907 <= w2137 and w6131;
w12908 <= not w12906 and not w12907;
w12909 <= not w12905 and not w12908;
w12910 <= a(50) and not w12909;
w12911 <= a(27) and w12910;
w12912 <= not w12905 and not w12909;
w12913 <= a(28) and a(49);
w12914 <= a(29) and a(48);
w12915 <= not w12913 and not w12914;
w12916 <= w12912 and not w12915;
w12917 <= not w12911 and not w12916;
w12918 <= not w12904 and not w12917;
w12919 <= w12904 and w12917;
w12920 <= not w12918 and not w12919;
w12921 <= w12889 and w12920;
w12922 <= not w12889 and not w12920;
w12923 <= w12843 and not w12922;
w12924 <= not w12921 and w12923;
w12925 <= w12843 and not w12924;
w12926 <= not w12922 and not w12924;
w12927 <= not w12921 and w12926;
w12928 <= not w12925 and not w12927;
w12929 <= w12830 and not w12928;
w12930 <= not w12830 and w12928;
w12931 <= not w12599 and not w12706;
w12932 <= not w12617 and not w12701;
w12933 <= not w12566 and not w12593;
w12934 <= not w12585 and not w12589;
w12935 <= a(22) and a(55);
w12936 <= a(26) and a(51);
w12937 <= not w12935 and not w12936;
w12938 <= w12935 and w12936;
w12939 <= a(43) and not w12938;
w12940 <= a(34) and w12939;
w12941 <= not w12937 and w12940;
w12942 <= not w12938 and not w12941;
w12943 <= not w12937 and w12942;
w12944 <= a(43) and not w12941;
w12945 <= a(34) and w12944;
w12946 <= not w12943 and not w12945;
w12947 <= w1472 and w7505;
w12948 <= w1353 and w10711;
w12949 <= w1710 and w7239;
w12950 <= not w12948 and not w12949;
w12951 <= not w12947 and not w12950;
w12952 <= a(52) and not w12951;
w12953 <= a(25) and w12952;
w12954 <= a(23) and a(54);
w12955 <= a(24) and a(53);
w12956 <= not w12954 and not w12955;
w12957 <= not w12947 and not w12951;
w12958 <= not w12956 and w12957;
w12959 <= not w12953 and not w12958;
w12960 <= not w12946 and not w12959;
w12961 <= not w12946 and not w12960;
w12962 <= not w12959 and not w12960;
w12963 <= not w12961 and not w12962;
w12964 <= a(32) and a(45);
w12965 <= not w5257 and not w12964;
w12966 <= w2949 and w5519;
w12967 <= a(61) and not w12966;
w12968 <= a(16) and w12967;
w12969 <= not w12965 and w12968;
w12970 <= a(61) and not w12969;
w12971 <= a(16) and w12970;
w12972 <= not w12966 and not w12969;
w12973 <= not w12965 and w12972;
w12974 <= not w12971 and not w12973;
w12975 <= not w12963 and not w12974;
w12976 <= not w12963 and not w12975;
w12977 <= not w12974 and not w12975;
w12978 <= not w12976 and not w12977;
w12979 <= not w12611 and not w12613;
w12980 <= not w12978 and not w12979;
w12981 <= not w12978 and not w12980;
w12982 <= not w12979 and not w12980;
w12983 <= not w12981 and not w12982;
w12984 <= not w12934 and not w12983;
w12985 <= w12934 and not w12982;
w12986 <= not w12981 and w12985;
w12987 <= not w12984 and not w12986;
w12988 <= not w12933 and w12987;
w12989 <= w12933 and not w12987;
w12990 <= not w12988 and not w12989;
w12991 <= not w12932 and w12990;
w12992 <= w12932 and not w12990;
w12993 <= not w12991 and not w12992;
w12994 <= not w12931 and w12993;
w12995 <= w12931 and not w12993;
w12996 <= not w12994 and not w12995;
w12997 <= not w12930 and w12996;
w12998 <= not w12929 and w12997;
w12999 <= w12996 and not w12998;
w13000 <= not w12930 and not w12998;
w13001 <= not w12929 and w13000;
w13002 <= not w12999 and not w13001;
w13003 <= not w12782 and not w13002;
w13004 <= w12782 and w13002;
w13005 <= not w13003 and not w13004;
w13006 <= not w12554 and not w12777;
w13007 <= not w12776 and not w13006;
w13008 <= not w13005 and w13007;
w13009 <= w13005 and not w13007;
w13010 <= not w13008 and not w13009;
w13011 <= not w13004 and not w13007;
w13012 <= not w13003 and not w13011;
w13013 <= not w12994 and not w12998;
w13014 <= not w12842 and not w12924;
w13015 <= not w12803 and not w12825;
w13016 <= not w12834 and not w12838;
w13017 <= w1298 and w8791;
w13018 <= a(57) and a(60);
w13019 <= w3454 and w13018;
w13020 <= w955 and w9315;
w13021 <= not w13019 and not w13020;
w13022 <= not w13017 and not w13021;
w13023 <= not w13017 and not w13022;
w13024 <= a(19) and a(59);
w13025 <= a(21) and a(57);
w13026 <= not w13024 and not w13025;
w13027 <= w13023 and not w13026;
w13028 <= a(60) and not w13022;
w13029 <= a(18) and w13028;
w13030 <= not w13027 and not w13029;
w13031 <= w2140 and w6131;
w13032 <= w1847 and w9740;
w13033 <= w2137 and w6370;
w13034 <= not w13032 and not w13033;
w13035 <= not w13031 and not w13034;
w13036 <= a(51) and not w13035;
w13037 <= a(27) and w13036;
w13038 <= not w13031 and not w13035;
w13039 <= a(28) and a(50);
w13040 <= a(29) and a(49);
w13041 <= not w13039 and not w13040;
w13042 <= w13038 and not w13041;
w13043 <= not w13037 and not w13042;
w13044 <= not w13030 and not w13043;
w13045 <= not w13030 and not w13044;
w13046 <= not w13043 and not w13044;
w13047 <= not w13045 and not w13046;
w13048 <= w854 and w9527;
w13049 <= w799 and w9715;
w13050 <= w697 and w9598;
w13051 <= not w13049 and not w13050;
w13052 <= not w13048 and not w13051;
w13053 <= a(63) and not w13052;
w13054 <= a(15) and w13053;
w13055 <= not w13048 and not w13052;
w13056 <= a(16) and a(62);
w13057 <= a(17) and a(61);
w13058 <= not w13056 and not w13057;
w13059 <= w13055 and not w13058;
w13060 <= not w13054 and not w13059;
w13061 <= not w13047 and not w13060;
w13062 <= not w13047 and not w13061;
w13063 <= not w13060 and not w13061;
w13064 <= not w13062 and not w13063;
w13065 <= a(30) and a(48);
w13066 <= a(31) and a(47);
w13067 <= not w13065 and not w13066;
w13068 <= w2671 and w6058;
w13069 <= a(58) and not w13068;
w13070 <= a(20) and w13069;
w13071 <= not w13067 and w13070;
w13072 <= not w13068 and not w13071;
w13073 <= not w13067 and w13072;
w13074 <= a(58) and not w13071;
w13075 <= a(20) and w13074;
w13076 <= not w13073 and not w13075;
w13077 <= a(33) and a(45);
w13078 <= a(34) and a(44);
w13079 <= not w13077 and not w13078;
w13080 <= w3956 and w5519;
w13081 <= w3896 and w7553;
w13082 <= w2949 and w5366;
w13083 <= not w13081 and not w13082;
w13084 <= not w13080 and not w13083;
w13085 <= not w13080 and not w13084;
w13086 <= not w13079 and w13085;
w13087 <= w5364 and not w13084;
w13088 <= not w13086 and not w13087;
w13089 <= not w13076 and not w13088;
w13090 <= not w13076 and not w13089;
w13091 <= not w13088 and not w13089;
w13092 <= not w13090 and not w13091;
w13093 <= w1921 and w7227;
w13094 <= a(53) and a(56);
w13095 <= w5133 and w13094;
w13096 <= w1710 and w7505;
w13097 <= not w13095 and not w13096;
w13098 <= not w13093 and not w13097;
w13099 <= a(53) and not w13098;
w13100 <= a(25) and w13099;
w13101 <= a(22) and a(56);
w13102 <= not w12503 and not w13101;
w13103 <= not w13093 and not w13098;
w13104 <= not w13102 and w13103;
w13105 <= not w13100 and not w13104;
w13106 <= not w13092 and not w13105;
w13107 <= not w13092 and not w13106;
w13108 <= not w13105 and not w13106;
w13109 <= not w13107 and not w13108;
w13110 <= not w13064 and w13109;
w13111 <= w13064 and not w13109;
w13112 <= not w13110 and not w13111;
w13113 <= not w13016 and not w13112;
w13114 <= w13016 and w13112;
w13115 <= not w13113 and not w13114;
w13116 <= not w13015 and w13115;
w13117 <= w13015 and not w13115;
w13118 <= not w13116 and not w13117;
w13119 <= w13014 and not w13118;
w13120 <= not w13014 and w13118;
w13121 <= not w13119 and not w13120;
w13122 <= not w12829 and not w12929;
w13123 <= w13121 and not w13122;
w13124 <= not w13121 and w13122;
w13125 <= not w13123 and not w13124;
w13126 <= not w12988 and not w12991;
w13127 <= not w12639 and not w12901;
w13128 <= not w12918 and not w13127;
w13129 <= not w12870 and not w12882;
w13130 <= w13128 and w13129;
w13131 <= not w13128 and not w13129;
w13132 <= not w13130 and not w13131;
w13133 <= not w12960 and not w12975;
w13134 <= not w13132 and w13133;
w13135 <= w13132 and not w13133;
w13136 <= not w13134 and not w13135;
w13137 <= not w12820 and not w12822;
w13138 <= w13136 and not w13137;
w13139 <= not w13136 and w13137;
w13140 <= not w13138 and not w13139;
w13141 <= w12865 and w12877;
w13142 <= not w12865 and not w12877;
w13143 <= not w13141 and not w13142;
w13144 <= w12957 and not w13143;
w13145 <= not w12957 and w13143;
w13146 <= not w13144 and not w13145;
w13147 <= w12852 and w12912;
w13148 <= not w12852 and not w12912;
w13149 <= not w13147 and not w13148;
w13150 <= w12972 and not w13149;
w13151 <= not w12972 and w13149;
w13152 <= not w13150 and not w13151;
w13153 <= not w12813 and not w12816;
w13154 <= not w13152 and w13153;
w13155 <= w13152 and not w13153;
w13156 <= not w13154 and not w13155;
w13157 <= w13146 and w13156;
w13158 <= not w13146 and not w13156;
w13159 <= not w13157 and not w13158;
w13160 <= w13140 and w13159;
w13161 <= not w13140 and not w13159;
w13162 <= not w13160 and not w13161;
w13163 <= w13126 and not w13162;
w13164 <= not w13126 and w13162;
w13165 <= not w13163 and not w13164;
w13166 <= not w12980 and not w12984;
w13167 <= not w12888 and not w12921;
w13168 <= not w13166 and not w13167;
w13169 <= not w13166 and not w13168;
w13170 <= not w13167 and not w13168;
w13171 <= not w13169 and not w13170;
w13172 <= a(36) and a(42);
w13173 <= not w5451 and not w13172;
w13174 <= w3634 and w4824;
w13175 <= a(55) and not w13174;
w13176 <= a(23) and w13175;
w13177 <= not w13173 and w13176;
w13178 <= not w13174 and not w13177;
w13179 <= not w13173 and w13178;
w13180 <= a(55) and not w13177;
w13181 <= a(23) and w13180;
w13182 <= not w13179 and not w13181;
w13183 <= a(26) and a(52);
w13184 <= w3609 and w13183;
w13185 <= w5752 and w13183;
w13186 <= w4371 and w5219;
w13187 <= not w13185 and not w13186;
w13188 <= not w13184 and not w13187;
w13189 <= w5752 and not w13188;
w13190 <= not w13184 and not w13188;
w13191 <= not w3609 and not w13183;
w13192 <= w13190 and not w13191;
w13193 <= not w13189 and not w13192;
w13194 <= not w13182 and not w13193;
w13195 <= not w13182 and not w13194;
w13196 <= not w13193 and not w13194;
w13197 <= not w13195 and not w13196;
w13198 <= not w12807 and not w12810;
w13199 <= w13197 and w13198;
w13200 <= not w13197 and not w13198;
w13201 <= not w13199 and not w13200;
w13202 <= w12897 and w12942;
w13203 <= not w12897 and not w12942;
w13204 <= not w13202 and not w13203;
w13205 <= not w12784 and not w12790;
w13206 <= not w13204 and w13205;
w13207 <= w13204 and not w13205;
w13208 <= not w13206 and not w13207;
w13209 <= not w12796 and not w12800;
w13210 <= not w13208 and w13209;
w13211 <= w13208 and not w13209;
w13212 <= not w13210 and not w13211;
w13213 <= w13201 and w13212;
w13214 <= not w13201 and not w13212;
w13215 <= not w13213 and not w13214;
w13216 <= not w13171 and w13215;
w13217 <= not w13171 and not w13216;
w13218 <= w13215 and not w13216;
w13219 <= not w13217 and not w13218;
w13220 <= w13165 and not w13219;
w13221 <= not w13165 and w13219;
w13222 <= w13125 and not w13221;
w13223 <= not w13220 and w13222;
w13224 <= w13125 and not w13223;
w13225 <= not w13221 and not w13223;
w13226 <= not w13220 and w13225;
w13227 <= not w13224 and not w13226;
w13228 <= not w13013 and not w13227;
w13229 <= w13013 and w13227;
w13230 <= not w13228 and not w13229;
w13231 <= not w13012 and w13230;
w13232 <= w13012 and not w13230;
w13233 <= not w13231 and not w13232;
w13234 <= not w13123 and not w13223;
w13235 <= not w13168 and not w13216;
w13236 <= not w13064 and not w13109;
w13237 <= not w13113 and not w13236;
w13238 <= w13023 and w13038;
w13239 <= not w13023 and not w13038;
w13240 <= not w13238 and not w13239;
w13241 <= w13103 and not w13240;
w13242 <= not w13103 and w13240;
w13243 <= not w13241 and not w13242;
w13244 <= not w13194 and not w13200;
w13245 <= not w13243 and w13244;
w13246 <= w13243 and not w13244;
w13247 <= not w13245 and not w13246;
w13248 <= a(34) and a(45);
w13249 <= a(35) and a(44);
w13250 <= not w13248 and not w13249;
w13251 <= w3125 and w5519;
w13252 <= a(63) and not w13251;
w13253 <= a(16) and w13252;
w13254 <= not w13250 and w13253;
w13255 <= not w13251 and not w13254;
w13256 <= not w13250 and w13255;
w13257 <= a(63) and not w13254;
w13258 <= a(16) and w13257;
w13259 <= not w13256 and not w13258;
w13260 <= a(36) and a(43);
w13261 <= a(23) and a(56);
w13262 <= a(27) and a(52);
w13263 <= not w13261 and not w13262;
w13264 <= a(27) and a(56);
w13265 <= w12363 and w13264;
w13266 <= w13260 and not w13265;
w13267 <= not w13263 and w13266;
w13268 <= w13260 and not w13267;
w13269 <= not w13265 and not w13267;
w13270 <= not w13263 and w13269;
w13271 <= not w13268 and not w13270;
w13272 <= not w13259 and not w13271;
w13273 <= not w13259 and not w13272;
w13274 <= not w13271 and not w13272;
w13275 <= not w13273 and not w13274;
w13276 <= not w13203 and not w13207;
w13277 <= w13275 and w13276;
w13278 <= not w13275 and not w13276;
w13279 <= not w13277 and not w13278;
w13280 <= w13247 and w13279;
w13281 <= not w13247 and not w13279;
w13282 <= not w13280 and not w13281;
w13283 <= w13237 and not w13282;
w13284 <= not w13237 and w13282;
w13285 <= not w13283 and not w13284;
w13286 <= not w13089 and not w13106;
w13287 <= a(18) and a(61);
w13288 <= not w13190 and w13287;
w13289 <= w13190 and not w13287;
w13290 <= not w13288 and not w13289;
w13291 <= w13178 and not w13290;
w13292 <= not w13178 and w13290;
w13293 <= not w13291 and not w13292;
w13294 <= w13055 and w13072;
w13295 <= not w13055 and not w13072;
w13296 <= not w13294 and not w13295;
w13297 <= w13085 and not w13296;
w13298 <= not w13085 and w13296;
w13299 <= not w13297 and not w13298;
w13300 <= w13293 and w13299;
w13301 <= not w13293 and not w13299;
w13302 <= not w13300 and not w13301;
w13303 <= not w13286 and w13302;
w13304 <= w13286 and not w13302;
w13305 <= not w13303 and not w13304;
w13306 <= w13285 and w13305;
w13307 <= not w13285 and not w13305;
w13308 <= not w13306 and not w13307;
w13309 <= w13235 and not w13308;
w13310 <= not w13235 and w13308;
w13311 <= not w13309 and not w13310;
w13312 <= not w13116 and not w13120;
w13313 <= not w13311 and w13312;
w13314 <= w13311 and not w13312;
w13315 <= not w13313 and not w13314;
w13316 <= not w13164 and not w13220;
w13317 <= not w13138 and not w13160;
w13318 <= not w13155 and not w13157;
w13319 <= w2269 and w7505;
w13320 <= w2107 and w7503;
w13321 <= w1710 and w7507;
w13322 <= not w13320 and not w13321;
w13323 <= not w13319 and not w13322;
w13324 <= not w13319 and not w13323;
w13325 <= a(25) and a(54);
w13326 <= a(26) and a(53);
w13327 <= not w13325 and not w13326;
w13328 <= w13324 and not w13327;
w13329 <= a(55) and not w13323;
w13330 <= a(24) and w13329;
w13331 <= not w13328 and not w13330;
w13332 <= a(37) and a(42);
w13333 <= w4889 and w5219;
w13334 <= w3977 and w13332;
w13335 <= w4371 and w5150;
w13336 <= not w13334 and not w13335;
w13337 <= not w13333 and not w13336;
w13338 <= w13332 and not w13337;
w13339 <= not w13333 and not w13337;
w13340 <= a(38) and a(41);
w13341 <= not w3977 and not w13340;
w13342 <= w13339 and not w13341;
w13343 <= not w13338 and not w13342;
w13344 <= not w13331 and not w13343;
w13345 <= not w13331 and not w13344;
w13346 <= not w13343 and not w13344;
w13347 <= not w13345 and not w13346;
w13348 <= a(17) and a(62);
w13349 <= not a(40) and not w13348;
w13350 <= a(40) and a(62);
w13351 <= a(17) and w13350;
w13352 <= a(51) and not w13351;
w13353 <= a(28) and w13352;
w13354 <= not w13349 and w13353;
w13355 <= a(51) and not w13354;
w13356 <= a(28) and w13355;
w13357 <= not w13351 and not w13354;
w13358 <= not w13349 and w13357;
w13359 <= not w13356 and not w13358;
w13360 <= not w13347 and not w13359;
w13361 <= not w13347 and not w13360;
w13362 <= not w13359 and not w13360;
w13363 <= not w13361 and not w13362;
w13364 <= w1300 and w8793;
w13365 <= w1298 and w9895;
w13366 <= w1296 and w9315;
w13367 <= not w13365 and not w13366;
w13368 <= not w13364 and not w13367;
w13369 <= not w13364 and not w13368;
w13370 <= a(20) and a(59);
w13371 <= a(21) and a(58);
w13372 <= not w13370 and not w13371;
w13373 <= w13369 and not w13372;
w13374 <= a(60) and not w13368;
w13375 <= a(19) and w13374;
w13376 <= not w13373 and not w13375;
w13377 <= a(22) and a(57);
w13378 <= a(29) and a(50);
w13379 <= a(30) and a(49);
w13380 <= not w13378 and not w13379;
w13381 <= w2423 and w6131;
w13382 <= w13377 and not w13381;
w13383 <= not w13380 and w13382;
w13384 <= w13377 and not w13383;
w13385 <= not w13381 and not w13383;
w13386 <= not w13380 and w13385;
w13387 <= not w13384 and not w13386;
w13388 <= not w13376 and not w13387;
w13389 <= not w13376 and not w13388;
w13390 <= not w13387 and not w13388;
w13391 <= not w13389 and not w13390;
w13392 <= w2949 and w5472;
w13393 <= w2404 and w8384;
w13394 <= w3618 and w6058;
w13395 <= not w13393 and not w13394;
w13396 <= not w13392 and not w13395;
w13397 <= a(48) and not w13396;
w13398 <= a(31) and w13397;
w13399 <= a(32) and a(47);
w13400 <= not w5702 and not w13399;
w13401 <= not w13392 and not w13396;
w13402 <= not w13400 and w13401;
w13403 <= not w13398 and not w13402;
w13404 <= not w13391 and not w13403;
w13405 <= not w13391 and not w13404;
w13406 <= not w13403 and not w13404;
w13407 <= not w13405 and not w13406;
w13408 <= w13363 and w13407;
w13409 <= not w13363 and not w13407;
w13410 <= not w13408 and not w13409;
w13411 <= not w13318 and w13410;
w13412 <= w13318 and not w13410;
w13413 <= not w13411 and not w13412;
w13414 <= w13317 and not w13413;
w13415 <= not w13317 and w13413;
w13416 <= not w13414 and not w13415;
w13417 <= not w13148 and not w13151;
w13418 <= not w13142 and not w13145;
w13419 <= w13417 and w13418;
w13420 <= not w13417 and not w13418;
w13421 <= not w13419 and not w13420;
w13422 <= not w13044 and not w13061;
w13423 <= not w13421 and w13422;
w13424 <= w13421 and not w13422;
w13425 <= not w13423 and not w13424;
w13426 <= not w13131 and not w13135;
w13427 <= not w13425 and w13426;
w13428 <= w13425 and not w13426;
w13429 <= not w13427 and not w13428;
w13430 <= not w13211 and not w13213;
w13431 <= w13429 and not w13430;
w13432 <= not w13429 and w13430;
w13433 <= not w13431 and not w13432;
w13434 <= w13416 and w13433;
w13435 <= not w13416 and not w13433;
w13436 <= not w13434 and not w13435;
w13437 <= not w13316 and w13436;
w13438 <= w13436 and not w13437;
w13439 <= not w13316 and not w13437;
w13440 <= not w13438 and not w13439;
w13441 <= w13315 and not w13440;
w13442 <= not w13315 and not w13439;
w13443 <= not w13438 and w13442;
w13444 <= not w13441 and not w13443;
w13445 <= not w13234 and w13444;
w13446 <= w13234 and not w13444;
w13447 <= not w13445 and not w13446;
w13448 <= not w13012 and not w13229;
w13449 <= not w13228 and not w13448;
w13450 <= not w13447 and w13449;
w13451 <= w13447 and not w13449;
w13452 <= not w13450 and not w13451;
w13453 <= not w13446 and not w13449;
w13454 <= not w13445 and not w13453;
w13455 <= not w13437 and not w13441;
w13456 <= not w13310 and not w13314;
w13457 <= not w13284 and not w13306;
w13458 <= not w13428 and not w13431;
w13459 <= a(17) and a(63);
w13460 <= a(29) and a(51);
w13461 <= not w13459 and not w13460;
w13462 <= a(29) and a(63);
w13463 <= w7578 and w13462;
w13464 <= a(33) and not w13463;
w13465 <= a(47) and w13464;
w13466 <= not w13461 and w13465;
w13467 <= not w13463 and not w13466;
w13468 <= not w13461 and w13467;
w13469 <= a(47) and not w13466;
w13470 <= a(33) and w13469;
w13471 <= not w13468 and not w13470;
w13472 <= w3634 and w5519;
w13473 <= w4401 and w7553;
w13474 <= w3125 and w5366;
w13475 <= not w13473 and not w13474;
w13476 <= not w13472 and not w13475;
w13477 <= a(46) and not w13476;
w13478 <= a(34) and w13477;
w13479 <= not w13472 and not w13476;
w13480 <= not w5654 and not w5739;
w13481 <= w13479 and not w13480;
w13482 <= not w13478 and not w13481;
w13483 <= not w13471 and not w13482;
w13484 <= not w13471 and not w13483;
w13485 <= not w13482 and not w13483;
w13486 <= not w13484 and not w13485;
w13487 <= w955 and w9527;
w13488 <= a(61) and not w13487;
w13489 <= a(19) and w13488;
w13490 <= a(62) and not w13487;
w13491 <= a(18) and w13490;
w13492 <= not w13489 and not w13491;
w13493 <= not w13357 and not w13492;
w13494 <= not w13357 and not w13493;
w13495 <= not w13492 and not w13493;
w13496 <= not w13494 and not w13495;
w13497 <= not w13486 and w13496;
w13498 <= w13486 and not w13496;
w13499 <= not w13497 and not w13498;
w13500 <= w1380 and w8793;
w13501 <= w1499 and w9895;
w13502 <= w1300 and w9315;
w13503 <= not w13501 and not w13502;
w13504 <= not w13500 and not w13503;
w13505 <= a(21) and a(59);
w13506 <= a(22) and a(58);
w13507 <= not w13505 and not w13506;
w13508 <= not w13500 and not w13507;
w13509 <= a(20) and a(60);
w13510 <= not w13508 and not w13509;
w13511 <= not w13504 and not w13510;
w13512 <= not w13339 and w13511;
w13513 <= w13339 and not w13511;
w13514 <= not w13512 and not w13513;
w13515 <= w3618 and w6062;
w13516 <= w2294 and w5694;
w13517 <= w2671 and w6131;
w13518 <= not w13516 and not w13517;
w13519 <= not w13515 and not w13518;
w13520 <= a(50) and not w13519;
w13521 <= a(30) and w13520;
w13522 <= not w13515 and not w13519;
w13523 <= a(31) and a(49);
w13524 <= a(32) and a(48);
w13525 <= not w13523 and not w13524;
w13526 <= w13522 and not w13525;
w13527 <= not w13521 and not w13526;
w13528 <= w13514 and not w13527;
w13529 <= w13514 and not w13528;
w13530 <= not w13527 and not w13528;
w13531 <= not w13529 and not w13530;
w13532 <= a(24) and a(56);
w13533 <= a(26) and a(54);
w13534 <= not w13532 and not w13533;
w13535 <= w2107 and w7227;
w13536 <= a(54) and a(57);
w13537 <= w2109 and w13536;
w13538 <= w1472 and w8006;
w13539 <= not w13537 and not w13538;
w13540 <= not w13535 and not w13539;
w13541 <= not w13535 and not w13540;
w13542 <= not w13534 and w13541;
w13543 <= a(57) and not w13540;
w13544 <= a(23) and w13543;
w13545 <= not w13542 and not w13544;
w13546 <= a(25) and a(55);
w13547 <= a(37) and a(43);
w13548 <= a(38) and a(42);
w13549 <= not w13547 and not w13548;
w13550 <= w4371 and w4824;
w13551 <= w13546 and not w13550;
w13552 <= not w13549 and w13551;
w13553 <= w13546 and not w13552;
w13554 <= not w13550 and not w13552;
w13555 <= not w13549 and w13554;
w13556 <= not w13553 and not w13555;
w13557 <= not w13545 and not w13556;
w13558 <= not w13545 and not w13557;
w13559 <= not w13556 and not w13557;
w13560 <= not w13558 and not w13559;
w13561 <= a(27) and a(53);
w13562 <= a(28) and a(52);
w13563 <= not w13561 and not w13562;
w13564 <= w2137 and w7239;
w13565 <= w3790 and not w13564;
w13566 <= not w13563 and w13565;
w13567 <= w3790 and not w13566;
w13568 <= not w13564 and not w13566;
w13569 <= not w13563 and w13568;
w13570 <= not w13567 and not w13569;
w13571 <= not w13560 and not w13570;
w13572 <= not w13560 and not w13571;
w13573 <= not w13570 and not w13571;
w13574 <= not w13572 and not w13573;
w13575 <= not w13531 and w13574;
w13576 <= w13531 and not w13574;
w13577 <= not w13575 and not w13576;
w13578 <= not w13499 and not w13577;
w13579 <= w13499 and w13577;
w13580 <= not w13578 and not w13579;
w13581 <= not w13458 and w13580;
w13582 <= w13458 and not w13580;
w13583 <= not w13581 and not w13582;
w13584 <= not w13457 and w13583;
w13585 <= w13457 and not w13583;
w13586 <= not w13584 and not w13585;
w13587 <= w13456 and not w13586;
w13588 <= not w13456 and w13586;
w13589 <= not w13587 and not w13588;
w13590 <= not w13415 and not w13434;
w13591 <= not w13239 and not w13242;
w13592 <= not w13295 and not w13298;
w13593 <= w13591 and w13592;
w13594 <= not w13591 and not w13592;
w13595 <= not w13593 and not w13594;
w13596 <= not w13288 and not w13292;
w13597 <= not w13595 and w13596;
w13598 <= w13595 and not w13596;
w13599 <= not w13597 and not w13598;
w13600 <= not w13246 and not w13280;
w13601 <= not w13300 and not w13303;
w13602 <= not w13600 and not w13601;
w13603 <= not w13600 and not w13602;
w13604 <= not w13601 and not w13602;
w13605 <= not w13603 and not w13604;
w13606 <= not w13599 and w13605;
w13607 <= w13599 and not w13605;
w13608 <= not w13606 and not w13607;
w13609 <= not w13409 and not w13411;
w13610 <= w13255 and w13324;
w13611 <= not w13255 and not w13324;
w13612 <= not w13610 and not w13611;
w13613 <= w13269 and not w13612;
w13614 <= not w13269 and w13612;
w13615 <= not w13613 and not w13614;
w13616 <= not w13272 and not w13278;
w13617 <= not w13615 and w13616;
w13618 <= w13615 and not w13616;
w13619 <= not w13617 and not w13618;
w13620 <= not w13420 and not w13424;
w13621 <= not w13619 and w13620;
w13622 <= w13619 and not w13620;
w13623 <= not w13621 and not w13622;
w13624 <= not w13609 and w13623;
w13625 <= w13609 and not w13623;
w13626 <= not w13624 and not w13625;
w13627 <= w13369 and w13385;
w13628 <= not w13369 and not w13385;
w13629 <= not w13627 and not w13628;
w13630 <= w13401 and not w13629;
w13631 <= not w13401 and w13629;
w13632 <= not w13630 and not w13631;
w13633 <= not w13344 and not w13360;
w13634 <= not w13388 and not w13404;
w13635 <= w13633 and w13634;
w13636 <= not w13633 and not w13634;
w13637 <= not w13635 and not w13636;
w13638 <= w13632 and w13637;
w13639 <= not w13632 and not w13637;
w13640 <= not w13638 and not w13639;
w13641 <= w13626 and w13640;
w13642 <= not w13626 and not w13640;
w13643 <= not w13641 and not w13642;
w13644 <= w13608 and w13643;
w13645 <= w13643 and not w13644;
w13646 <= w13608 and not w13644;
w13647 <= not w13645 and not w13646;
w13648 <= not w13590 and not w13647;
w13649 <= w13590 and not w13646;
w13650 <= not w13645 and w13649;
w13651 <= not w13648 and not w13650;
w13652 <= w13589 and w13651;
w13653 <= not w13589 and not w13651;
w13654 <= not w13652 and not w13653;
w13655 <= w13455 and not w13654;
w13656 <= not w13455 and w13654;
w13657 <= not w13655 and not w13656;
w13658 <= w13454 and not w13657;
w13659 <= not w13454 and not w13655;
w13660 <= not w13656 and w13659;
w13661 <= not w13658 and not w13660;
w13662 <= not w13656 and not w13659;
w13663 <= not w13644 and not w13648;
w13664 <= not w13624 and not w13641;
w13665 <= not w13602 and not w13607;
w13666 <= a(41) and a(62);
w13667 <= a(19) and w13666;
w13668 <= w5219 and not w13667;
w13669 <= not w13667 and not w13668;
w13670 <= a(19) and a(62);
w13671 <= not a(41) and not w13670;
w13672 <= w13669 and not w13671;
w13673 <= w5219 and not w13668;
w13674 <= not w13672 and not w13673;
w13675 <= w1353 and w7748;
w13676 <= a(56) and a(59);
w13677 <= w5133 and w13676;
w13678 <= w1725 and w8793;
w13679 <= not w13677 and not w13678;
w13680 <= not w13675 and not w13679;
w13681 <= a(59) and not w13680;
w13682 <= a(22) and w13681;
w13683 <= not w13675 and not w13680;
w13684 <= a(23) and a(58);
w13685 <= not w12162 and not w13684;
w13686 <= w13683 and not w13685;
w13687 <= not w13682 and not w13686;
w13688 <= not w13674 and not w13687;
w13689 <= not w13674 and not w13688;
w13690 <= not w13687 and not w13688;
w13691 <= not w13689 and not w13690;
w13692 <= a(33) and a(48);
w13693 <= a(34) and a(47);
w13694 <= not w13692 and not w13693;
w13695 <= w3956 and w6058;
w13696 <= w10107 and not w13695;
w13697 <= not w13694 and w13696;
w13698 <= w10107 and not w13697;
w13699 <= not w13695 and not w13697;
w13700 <= not w13694 and w13699;
w13701 <= not w13698 and not w13700;
w13702 <= not w13691 and not w13701;
w13703 <= not w13691 and not w13702;
w13704 <= not w13701 and not w13702;
w13705 <= not w13703 and not w13704;
w13706 <= not w13594 and not w13598;
w13707 <= w13705 and w13706;
w13708 <= not w13705 and not w13706;
w13709 <= not w13707 and not w13708;
w13710 <= w1300 and w9318;
w13711 <= w3454 and w11440;
w13712 <= w1137 and w9715;
w13713 <= not w13711 and not w13712;
w13714 <= not w13710 and not w13713;
w13715 <= not w13710 and not w13714;
w13716 <= a(20) and a(61);
w13717 <= a(21) and a(60);
w13718 <= not w13716 and not w13717;
w13719 <= w13715 and not w13718;
w13720 <= a(63) and not w13714;
w13721 <= a(18) and w13720;
w13722 <= not w13719 and not w13721;
w13723 <= a(35) and a(46);
w13724 <= w3493 and w5519;
w13725 <= w3634 and w5366;
w13726 <= a(37) and a(44);
w13727 <= w13723 and w13726;
w13728 <= not w13725 and not w13727;
w13729 <= not w13724 and not w13728;
w13730 <= w13723 and not w13729;
w13731 <= a(36) and a(45);
w13732 <= not w13726 and not w13731;
w13733 <= not w13724 and not w13729;
w13734 <= not w13732 and w13733;
w13735 <= not w13730 and not w13734;
w13736 <= not w13722 and not w13735;
w13737 <= not w13722 and not w13736;
w13738 <= not w13735 and not w13736;
w13739 <= not w13737 and not w13738;
w13740 <= a(29) and w13183;
w13741 <= a(53) and w2606;
w13742 <= not w13740 and not w13741;
w13743 <= w2140 and w7239;
w13744 <= a(55) and not w13743;
w13745 <= not w13742 and w13744;
w13746 <= a(55) and not w13745;
w13747 <= a(26) and w13746;
w13748 <= a(28) and a(53);
w13749 <= a(29) and a(52);
w13750 <= not w13748 and not w13749;
w13751 <= not w13743 and not w13745;
w13752 <= not w13750 and w13751;
w13753 <= not w13747 and not w13752;
w13754 <= not w13739 and not w13753;
w13755 <= not w13739 and not w13754;
w13756 <= not w13753 and not w13754;
w13757 <= not w13755 and not w13756;
w13758 <= not w13709 and w13757;
w13759 <= w13709 and not w13757;
w13760 <= not w13758 and not w13759;
w13761 <= not w13665 and w13760;
w13762 <= not w13665 and not w13761;
w13763 <= w13760 and not w13761;
w13764 <= not w13762 and not w13763;
w13765 <= not w13664 and not w13764;
w13766 <= not w13664 and not w13765;
w13767 <= not w13764 and not w13765;
w13768 <= not w13766 and not w13767;
w13769 <= not w13663 and not w13768;
w13770 <= not w13663 and not w13769;
w13771 <= not w13768 and not w13769;
w13772 <= not w13770 and not w13771;
w13773 <= not w13581 and not w13584;
w13774 <= not w13628 and not w13631;
w13775 <= a(27) and a(54);
w13776 <= a(38) and a(43);
w13777 <= a(39) and a(42);
w13778 <= not w13776 and not w13777;
w13779 <= w4824 and w4889;
w13780 <= w13775 and not w13779;
w13781 <= not w13778 and w13780;
w13782 <= w13775 and not w13781;
w13783 <= not w13779 and not w13781;
w13784 <= not w13778 and w13783;
w13785 <= not w13782 and not w13784;
w13786 <= not w13774 and not w13785;
w13787 <= not w13774 and not w13786;
w13788 <= not w13785 and not w13786;
w13789 <= not w13787 and not w13788;
w13790 <= not w13611 and not w13614;
w13791 <= w13789 and w13790;
w13792 <= not w13789 and not w13790;
w13793 <= not w13791 and not w13792;
w13794 <= not w13618 and not w13622;
w13795 <= not w13636 and not w13638;
w13796 <= not w13794 and not w13795;
w13797 <= not w13794 and not w13796;
w13798 <= not w13795 and not w13796;
w13799 <= not w13797 and not w13798;
w13800 <= w13793 and not w13799;
w13801 <= not w13793 and w13799;
w13802 <= not w13773 and not w13801;
w13803 <= not w13800 and w13802;
w13804 <= not w13773 and not w13803;
w13805 <= not w13801 and not w13803;
w13806 <= not w13800 and w13805;
w13807 <= not w13804 and not w13806;
w13808 <= not w13487 and not w13493;
w13809 <= w13479 and w13808;
w13810 <= not w13479 and not w13808;
w13811 <= not w13809 and not w13810;
w13812 <= w3618 and w6131;
w13813 <= w2294 and w9740;
w13814 <= w2671 and w6370;
w13815 <= not w13813 and not w13814;
w13816 <= not w13812 and not w13815;
w13817 <= a(51) and not w13816;
w13818 <= a(30) and w13817;
w13819 <= not w13812 and not w13816;
w13820 <= a(31) and a(50);
w13821 <= a(32) and a(49);
w13822 <= not w13820 and not w13821;
w13823 <= w13819 and not w13822;
w13824 <= not w13818 and not w13823;
w13825 <= w13811 and not w13824;
w13826 <= w13811 and not w13825;
w13827 <= not w13824 and not w13825;
w13828 <= not w13826 and not w13827;
w13829 <= w13467 and w13522;
w13830 <= not w13467 and not w13522;
w13831 <= not w13829 and not w13830;
w13832 <= not w13500 and not w13504;
w13833 <= not w13831 and w13832;
w13834 <= w13831 and not w13832;
w13835 <= not w13833 and not w13834;
w13836 <= not w13486 and not w13496;
w13837 <= not w13483 and not w13836;
w13838 <= w13835 and not w13837;
w13839 <= not w13835 and w13837;
w13840 <= not w13838 and not w13839;
w13841 <= w13828 and w13840;
w13842 <= not w13828 and not w13840;
w13843 <= not w13841 and not w13842;
w13844 <= not w13531 and not w13574;
w13845 <= not w13578 and not w13844;
w13846 <= w13843 and w13845;
w13847 <= not w13843 and not w13845;
w13848 <= not w13846 and not w13847;
w13849 <= w13554 and w13568;
w13850 <= not w13554 and not w13568;
w13851 <= not w13849 and not w13850;
w13852 <= w13541 and not w13851;
w13853 <= not w13541 and w13851;
w13854 <= not w13852 and not w13853;
w13855 <= not w13557 and not w13571;
w13856 <= not w13512 and not w13528;
w13857 <= w13855 and w13856;
w13858 <= not w13855 and not w13856;
w13859 <= not w13857 and not w13858;
w13860 <= w13854 and w13859;
w13861 <= not w13854 and not w13859;
w13862 <= not w13860 and not w13861;
w13863 <= w13848 and w13862;
w13864 <= not w13848 and not w13862;
w13865 <= not w13863 and not w13864;
w13866 <= not w13807 and not w13865;
w13867 <= w13807 and w13865;
w13868 <= not w13866 and not w13867;
w13869 <= not w13772 and not w13868;
w13870 <= not w13772 and not w13869;
w13871 <= not w13868 and not w13869;
w13872 <= not w13870 and not w13871;
w13873 <= not w13588 and not w13652;
w13874 <= not w13872 and not w13873;
w13875 <= w13872 and w13873;
w13876 <= not w13874 and not w13875;
w13877 <= not w13662 and not w13876;
w13878 <= w13662 and w13876;
w13879 <= not w13877 and not w13878;
w13880 <= not w13662 and not w13875;
w13881 <= not w13874 and not w13880;
w13882 <= not w13769 and not w13869;
w13883 <= not w13807 and w13865;
w13884 <= not w13803 and not w13883;
w13885 <= not w13847 and not w13863;
w13886 <= not w13796 and not w13800;
w13887 <= a(51) and a(62);
w13888 <= w5904 and w13887;
w13889 <= w1300 and w9527;
w13890 <= not w13888 and not w13889;
w13891 <= a(31) and a(51);
w13892 <= a(21) and a(61);
w13893 <= w13891 and w13892;
w13894 <= not w13890 and not w13893;
w13895 <= not w13893 and not w13894;
w13896 <= not w13891 and not w13892;
w13897 <= w13895 and not w13896;
w13898 <= a(62) and not w13894;
w13899 <= a(20) and w13898;
w13900 <= not w13897 and not w13899;
w13901 <= w3956 and w6062;
w13902 <= w3896 and w5694;
w13903 <= w2949 and w6131;
w13904 <= not w13902 and not w13903;
w13905 <= not w13901 and not w13904;
w13906 <= a(50) and not w13905;
w13907 <= a(32) and w13906;
w13908 <= not w13901 and not w13905;
w13909 <= a(33) and a(49);
w13910 <= a(34) and a(48);
w13911 <= not w13909 and not w13910;
w13912 <= w13908 and not w13911;
w13913 <= not w13907 and not w13912;
w13914 <= not w13900 and not w13913;
w13915 <= not w13900 and not w13914;
w13916 <= not w13913 and not w13914;
w13917 <= not w13915 and not w13916;
w13918 <= w1472 and w8793;
w13919 <= w1921 and w9895;
w13920 <= w1725 and w9315;
w13921 <= not w13919 and not w13920;
w13922 <= not w13918 and not w13921;
w13923 <= a(60) and not w13922;
w13924 <= a(22) and w13923;
w13925 <= not w13918 and not w13922;
w13926 <= a(23) and a(59);
w13927 <= not w11221 and not w13926;
w13928 <= w13925 and not w13927;
w13929 <= not w13924 and not w13928;
w13930 <= not w13917 and not w13929;
w13931 <= not w13917 and not w13930;
w13932 <= not w13929 and not w13930;
w13933 <= not w13931 and not w13932;
w13934 <= not w13786 and not w13792;
w13935 <= w13933 and w13934;
w13936 <= not w13933 and not w13934;
w13937 <= not w13935 and not w13936;
w13938 <= a(38) and a(44);
w13939 <= a(39) and a(43);
w13940 <= not w13938 and not w13939;
w13941 <= w4889 and w5102;
w13942 <= a(56) and not w13941;
w13943 <= a(26) and w13942;
w13944 <= not w13940 and w13943;
w13945 <= not w13941 and not w13944;
w13946 <= not w13940 and w13945;
w13947 <= a(56) and not w13944;
w13948 <= a(26) and w13947;
w13949 <= not w13946 and not w13948;
w13950 <= a(29) and a(53);
w13951 <= a(30) and a(52);
w13952 <= not w13950 and not w13951;
w13953 <= w2423 and w7239;
w13954 <= w6259 and not w13953;
w13955 <= not w13952 and w13954;
w13956 <= w6259 and not w13955;
w13957 <= not w13953 and not w13955;
w13958 <= not w13952 and w13957;
w13959 <= not w13956 and not w13958;
w13960 <= not w13949 and not w13959;
w13961 <= not w13949 and not w13960;
w13962 <= not w13959 and not w13960;
w13963 <= not w13961 and not w13962;
w13964 <= w3493 and w5366;
w13965 <= a(37) and a(47);
w13966 <= w5654 and w13965;
w13967 <= w3634 and w5472;
w13968 <= not w13966 and not w13967;
w13969 <= not w13964 and not w13968;
w13970 <= a(47) and not w13969;
w13971 <= a(35) and w13970;
w13972 <= not w13964 and not w13969;
w13973 <= not w5952 and not w6243;
w13974 <= w13972 and not w13973;
w13975 <= not w13971 and not w13974;
w13976 <= not w13963 and not w13975;
w13977 <= not w13963 and not w13976;
w13978 <= not w13975 and not w13976;
w13979 <= not w13977 and not w13978;
w13980 <= not w13937 and w13979;
w13981 <= w13937 and not w13979;
w13982 <= not w13980 and not w13981;
w13983 <= not w13886 and w13982;
w13984 <= not w13886 and not w13983;
w13985 <= w13982 and not w13983;
w13986 <= not w13984 and not w13985;
w13987 <= not w13885 and not w13986;
w13988 <= not w13885 and not w13987;
w13989 <= not w13986 and not w13987;
w13990 <= not w13988 and not w13989;
w13991 <= not w13884 and not w13990;
w13992 <= not w13884 and not w13991;
w13993 <= not w13990 and not w13991;
w13994 <= not w13992 and not w13993;
w13995 <= not w13761 and not w13765;
w13996 <= not w13830 and not w13834;
w13997 <= w2439 and w11524;
w13998 <= w2137 and w7507;
w13999 <= a(25) and a(57);
w14000 <= w6925 and w13999;
w14001 <= not w13998 and not w14000;
w14002 <= not w13997 and not w14001;
w14003 <= w6925 and not w14002;
w14004 <= a(27) and a(55);
w14005 <= not w13999 and not w14004;
w14006 <= not w13997 and not w14002;
w14007 <= not w14005 and w14006;
w14008 <= not w14003 and not w14007;
w14009 <= not w13996 and not w14008;
w14010 <= not w13996 and not w14009;
w14011 <= not w14008 and not w14009;
w14012 <= not w14010 and not w14011;
w14013 <= not w13850 and not w13853;
w14014 <= w14012 and w14013;
w14015 <= not w14012 and not w14013;
w14016 <= not w14014 and not w14015;
w14017 <= not w13828 and w13840;
w14018 <= not w13838 and not w14017;
w14019 <= not w13858 and not w13860;
w14020 <= not w14018 and not w14019;
w14021 <= not w14018 and not w14020;
w14022 <= not w14019 and not w14020;
w14023 <= not w14021 and not w14022;
w14024 <= w14016 and not w14023;
w14025 <= not w14016 and w14023;
w14026 <= not w13995 and not w14025;
w14027 <= not w14024 and w14026;
w14028 <= not w13995 and not w14027;
w14029 <= not w14025 and not w14027;
w14030 <= not w14024 and w14029;
w14031 <= not w14028 and not w14030;
w14032 <= not w13708 and not w13759;
w14033 <= w13699 and w13819;
w14034 <= not w13699 and not w13819;
w14035 <= not w14033 and not w14034;
w14036 <= w13751 and not w14035;
w14037 <= not w13751 and w14035;
w14038 <= not w14036 and not w14037;
w14039 <= w13683 and w13715;
w14040 <= not w13683 and not w13715;
w14041 <= not w14039 and not w14040;
w14042 <= w13733 and not w14041;
w14043 <= not w13733 and w14041;
w14044 <= not w14042 and not w14043;
w14045 <= not w13736 and not w13754;
w14046 <= not w14044 and w14045;
w14047 <= w14044 and not w14045;
w14048 <= not w14046 and not w14047;
w14049 <= w14038 and w14048;
w14050 <= not w14038 and not w14048;
w14051 <= not w14049 and not w14050;
w14052 <= w14032 and not w14051;
w14053 <= not w14032 and w14051;
w14054 <= not w14052 and not w14053;
w14055 <= not w13810 and not w13825;
w14056 <= not w13688 and not w13702;
w14057 <= w14055 and w14056;
w14058 <= not w14055 and not w14056;
w14059 <= not w14057 and not w14058;
w14060 <= w12353 and not w13669;
w14061 <= not w12353 and w13669;
w14062 <= not w14060 and not w14061;
w14063 <= w13783 and not w14062;
w14064 <= not w13783 and w14062;
w14065 <= not w14063 and not w14064;
w14066 <= w14059 and w14065;
w14067 <= not w14059 and not w14065;
w14068 <= not w14066 and not w14067;
w14069 <= w14054 and w14068;
w14070 <= not w14054 and not w14068;
w14071 <= not w14069 and not w14070;
w14072 <= not w14031 and not w14071;
w14073 <= w14031 and w14071;
w14074 <= not w14072 and not w14073;
w14075 <= not w13994 and not w14074;
w14076 <= not w13994 and not w14075;
w14077 <= not w14074 and not w14075;
w14078 <= not w14076 and not w14077;
w14079 <= not w13882 and not w14078;
w14080 <= w13882 and w14078;
w14081 <= not w14079 and not w14080;
w14082 <= not w13881 and w14081;
w14083 <= w13881 and not w14081;
w14084 <= not w14082 and not w14083;
w14085 <= not w13991 and not w14075;
w14086 <= not w13936 and not w13981;
w14087 <= not w14047 and not w14049;
w14088 <= not w14086 and not w14087;
w14089 <= not w14086 and not w14088;
w14090 <= not w14087 and not w14088;
w14091 <= not w14089 and not w14090;
w14092 <= w13925 and w13972;
w14093 <= not w13925 and not w13972;
w14094 <= not w14092 and not w14093;
w14095 <= w13945 and not w14094;
w14096 <= not w13945 and w14094;
w14097 <= not w14095 and not w14096;
w14098 <= w13895 and w13908;
w14099 <= not w13895 and not w13908;
w14100 <= not w14098 and not w14099;
w14101 <= w14006 and not w14100;
w14102 <= not w14006 and w14100;
w14103 <= not w14101 and not w14102;
w14104 <= not w13960 and not w13976;
w14105 <= not w14103 and w14104;
w14106 <= w14103 and not w14104;
w14107 <= not w14105 and not w14106;
w14108 <= w14097 and w14107;
w14109 <= not w14097 and not w14107;
w14110 <= not w14108 and not w14109;
w14111 <= not w14091 and w14110;
w14112 <= not w14091 and not w14111;
w14113 <= w14110 and not w14111;
w14114 <= not w14112 and not w14113;
w14115 <= not w13983 and not w13987;
w14116 <= not w14034 and not w14037;
w14117 <= not w14040 and not w14043;
w14118 <= w14116 and w14117;
w14119 <= not w14116 and not w14117;
w14120 <= not w14118 and not w14119;
w14121 <= not w13914 and not w13930;
w14122 <= not w14120 and w14121;
w14123 <= w14120 and not w14121;
w14124 <= not w14122 and not w14123;
w14125 <= w1472 and w9315;
w14126 <= a(59) and not w14125;
w14127 <= a(24) and w14126;
w14128 <= a(60) and not w14125;
w14129 <= a(23) and w14128;
w14130 <= not w14127 and not w14129;
w14131 <= not w13957 and not w14130;
w14132 <= not w13957 and not w14131;
w14133 <= not w14130 and not w14131;
w14134 <= not w14132 and not w14133;
w14135 <= w2916 and w7503;
w14136 <= w2671 and w7239;
w14137 <= a(31) and a(55);
w14138 <= w13562 and w14137;
w14139 <= not w14136 and not w14138;
w14140 <= not w14135 and not w14139;
w14141 <= a(52) and not w14140;
w14142 <= a(31) and w14141;
w14143 <= a(28) and a(55);
w14144 <= a(30) and a(53);
w14145 <= not w14143 and not w14144;
w14146 <= not w14135 and not w14140;
w14147 <= not w14145 and w14146;
w14148 <= not w14142 and not w14147;
w14149 <= not w14134 and not w14148;
w14150 <= not w14134 and not w14149;
w14151 <= not w14148 and not w14149;
w14152 <= not w14150 and not w14151;
w14153 <= not w14060 and not w14064;
w14154 <= w14152 and w14153;
w14155 <= not w14152 and not w14153;
w14156 <= not w14154 and not w14155;
w14157 <= not w14058 and not w14066;
w14158 <= w14156 and not w14157;
w14159 <= not w14156 and w14157;
w14160 <= not w14158 and not w14159;
w14161 <= w14124 and w14160;
w14162 <= not w14124 and not w14160;
w14163 <= not w14161 and not w14162;
w14164 <= not w14115 and w14163;
w14165 <= w14115 and not w14163;
w14166 <= not w14164 and not w14165;
w14167 <= w14114 and w14166;
w14168 <= not w14114 and not w14166;
w14169 <= not w14167 and not w14168;
w14170 <= not w14031 and w14071;
w14171 <= not w14027 and not w14170;
w14172 <= not w14053 and not w14069;
w14173 <= not w14020 and not w14024;
w14174 <= a(42) and a(62);
w14175 <= a(21) and w14174;
w14176 <= w5150 and not w14175;
w14177 <= not w14175 and not w14176;
w14178 <= a(21) and a(62);
w14179 <= not a(42) and not w14178;
w14180 <= w14177 and not w14179;
w14181 <= w5150 and not w14176;
w14182 <= not w14180 and not w14181;
w14183 <= a(39) and a(44);
w14184 <= a(40) and a(43);
w14185 <= not w14183 and not w14184;
w14186 <= w3977 and w5102;
w14187 <= a(54) and not w14186;
w14188 <= a(29) and w14187;
w14189 <= not w14185 and w14188;
w14190 <= a(54) and not w14189;
w14191 <= a(29) and w14190;
w14192 <= not w14186 and not w14189;
w14193 <= not w14185 and w14192;
w14194 <= not w14191 and not w14193;
w14195 <= not w14182 and not w14194;
w14196 <= not w14182 and not w14195;
w14197 <= not w14194 and not w14195;
w14198 <= not w14196 and not w14197;
w14199 <= w3125 and w6062;
w14200 <= w2778 and w5694;
w14201 <= w3956 and w6131;
w14202 <= not w14200 and not w14201;
w14203 <= not w14199 and not w14202;
w14204 <= a(50) and not w14203;
w14205 <= a(33) and w14204;
w14206 <= not w14199 and not w14203;
w14207 <= a(34) and a(49);
w14208 <= a(35) and a(48);
w14209 <= not w14207 and not w14208;
w14210 <= w14206 and not w14209;
w14211 <= not w14205 and not w14210;
w14212 <= not w14198 and not w14211;
w14213 <= not w14198 and not w14212;
w14214 <= not w14211 and not w14212;
w14215 <= not w14213 and not w14214;
w14216 <= not w14009 and not w14015;
w14217 <= w14215 and w14216;
w14218 <= not w14215 and not w14216;
w14219 <= not w14217 and not w14218;
w14220 <= a(26) and a(57);
w14221 <= a(32) and a(51);
w14222 <= not w14220 and not w14221;
w14223 <= a(51) and a(57);
w14224 <= w3072 and w14223;
w14225 <= w2269 and w8242;
w14226 <= a(32) and a(58);
w14227 <= w12650 and w14226;
w14228 <= not w14225 and not w14227;
w14229 <= not w14224 and not w14228;
w14230 <= not w14224 and not w14229;
w14231 <= not w14222 and w14230;
w14232 <= a(58) and not w14229;
w14233 <= a(25) and w14232;
w14234 <= not w14231 and not w14233;
w14235 <= w4371 and w5366;
w14236 <= w3336 and w5056;
w14237 <= w3493 and w5472;
w14238 <= not w14236 and not w14237;
w14239 <= not w14235 and not w14238;
w14240 <= a(47) and not w14239;
w14241 <= a(36) and w14240;
w14242 <= not w14235 and not w14239;
w14243 <= a(37) and a(46);
w14244 <= a(38) and a(45);
w14245 <= not w14243 and not w14244;
w14246 <= w14242 and not w14245;
w14247 <= not w14241 and not w14246;
w14248 <= not w14234 and not w14247;
w14249 <= not w14234 and not w14248;
w14250 <= not w14247 and not w14248;
w14251 <= not w14249 and not w14250;
w14252 <= a(20) and a(63);
w14253 <= a(22) and a(61);
w14254 <= not w14252 and not w14253;
w14255 <= w1499 and w9715;
w14256 <= w13264 and not w14255;
w14257 <= not w14254 and w14256;
w14258 <= w13264 and not w14257;
w14259 <= not w14255 and not w14257;
w14260 <= not w14254 and w14259;
w14261 <= not w14258 and not w14260;
w14262 <= not w14251 and not w14261;
w14263 <= not w14251 and not w14262;
w14264 <= not w14261 and not w14262;
w14265 <= not w14263 and not w14264;
w14266 <= not w14219 and w14265;
w14267 <= w14219 and not w14265;
w14268 <= not w14266 and not w14267;
w14269 <= not w14173 and w14268;
w14270 <= w14173 and not w14268;
w14271 <= not w14269 and not w14270;
w14272 <= not w14172 and w14271;
w14273 <= w14172 and not w14271;
w14274 <= not w14272 and not w14273;
w14275 <= not w14171 and w14274;
w14276 <= w14171 and not w14274;
w14277 <= not w14275 and not w14276;
w14278 <= not w14169 and w14277;
w14279 <= w14277 and not w14278;
w14280 <= not w14169 and not w14278;
w14281 <= not w14279 and not w14280;
w14282 <= not w14085 and not w14281;
w14283 <= w14085 and w14281;
w14284 <= not w14282 and not w14283;
w14285 <= not w13881 and not w14080;
w14286 <= not w14079 and not w14285;
w14287 <= not w14284 and w14286;
w14288 <= w14284 and not w14286;
w14289 <= not w14287 and not w14288;
w14290 <= not w14283 and not w14286;
w14291 <= not w14282 and not w14290;
w14292 <= not w14275 and not w14278;
w14293 <= not w14114 and w14166;
w14294 <= not w14164 and not w14293;
w14295 <= not w14125 and not w14131;
w14296 <= w14259 and w14295;
w14297 <= not w14259 and not w14295;
w14298 <= not w14296 and not w14297;
w14299 <= a(31) and a(53);
w14300 <= a(32) and a(52);
w14301 <= not w14299 and not w14300;
w14302 <= w3618 and w7239;
w14303 <= w12409 and not w14302;
w14304 <= not w14301 and w14303;
w14305 <= w12409 and not w14304;
w14306 <= not w14302 and not w14304;
w14307 <= not w14301 and w14306;
w14308 <= not w14305 and not w14307;
w14309 <= w14298 and not w14308;
w14310 <= w14298 and not w14309;
w14311 <= not w14308 and not w14309;
w14312 <= not w14310 and not w14311;
w14313 <= not w14149 and not w14155;
w14314 <= w14312 and w14313;
w14315 <= not w14312 and not w14313;
w14316 <= not w14314 and not w14315;
w14317 <= not w14119 and not w14123;
w14318 <= not w14316 and w14317;
w14319 <= w14316 and not w14317;
w14320 <= not w14318 and not w14319;
w14321 <= not w14158 and not w14161;
w14322 <= not w14320 and w14321;
w14323 <= w14320 and not w14321;
w14324 <= not w14322 and not w14323;
w14325 <= w1725 and w9527;
w14326 <= w1173 and w9715;
w14327 <= w1380 and w9598;
w14328 <= not w14326 and not w14327;
w14329 <= not w14325 and not w14328;
w14330 <= not w14325 and not w14329;
w14331 <= a(22) and a(62);
w14332 <= a(23) and a(61);
w14333 <= not w14331 and not w14332;
w14334 <= w14330 and not w14333;
w14335 <= a(63) and not w14329;
w14336 <= a(21) and w14335;
w14337 <= not w14334 and not w14336;
w14338 <= a(24) and a(60);
w14339 <= a(25) and a(59);
w14340 <= not w14338 and not w14339;
w14341 <= w1710 and w9315;
w14342 <= a(33) and not w14341;
w14343 <= a(51) and w14342;
w14344 <= not w14340 and w14343;
w14345 <= a(51) and not w14344;
w14346 <= a(33) and w14345;
w14347 <= not w14341 and not w14344;
w14348 <= not w14340 and w14347;
w14349 <= not w14346 and not w14348;
w14350 <= not w14337 and not w14349;
w14351 <= not w14337 and not w14350;
w14352 <= not w14349 and not w14350;
w14353 <= not w14351 and not w14352;
w14354 <= w3634 and w6062;
w14355 <= w4401 and w5694;
w14356 <= w3125 and w6131;
w14357 <= not w14355 and not w14356;
w14358 <= not w14354 and not w14357;
w14359 <= a(50) and not w14358;
w14360 <= a(34) and w14359;
w14361 <= not w14354 and not w14358;
w14362 <= a(35) and a(49);
w14363 <= a(36) and a(48);
w14364 <= not w14362 and not w14363;
w14365 <= w14361 and not w14364;
w14366 <= not w14360 and not w14365;
w14367 <= not w14353 and not w14366;
w14368 <= not w14353 and not w14367;
w14369 <= not w14366 and not w14367;
w14370 <= not w14368 and not w14369;
w14371 <= a(29) and a(55);
w14372 <= a(38) and a(46);
w14373 <= not w14371 and not w14372;
w14374 <= w2140 and w8967;
w14375 <= a(38) and a(56);
w14376 <= w12183 and w14375;
w14377 <= not w14374 and not w14376;
w14378 <= w14371 and w14372;
w14379 <= not w14377 and not w14378;
w14380 <= not w14378 and not w14379;
w14381 <= not w14373 and w14380;
w14382 <= a(56) and not w14379;
w14383 <= a(28) and w14382;
w14384 <= not w14381 and not w14383;
w14385 <= w5102 and w5219;
w14386 <= w3790 and w4617;
w14387 <= w3977 and w5519;
w14388 <= not w14386 and not w14387;
w14389 <= not w14385 and not w14388;
w14390 <= a(45) and not w14389;
w14391 <= a(39) and w14390;
w14392 <= not w14385 and not w14389;
w14393 <= a(40) and a(44);
w14394 <= not w4613 and not w14393;
w14395 <= w14392 and not w14394;
w14396 <= not w14391 and not w14395;
w14397 <= not w14384 and not w14396;
w14398 <= not w14384 and not w14397;
w14399 <= not w14396 and not w14397;
w14400 <= not w14398 and not w14399;
w14401 <= a(27) and a(57);
w14402 <= a(30) and a(54);
w14403 <= not w14401 and not w14402;
w14404 <= a(30) and a(57);
w14405 <= w13775 and w14404;
w14406 <= w13965 and not w14405;
w14407 <= not w14403 and w14406;
w14408 <= w13965 and not w14407;
w14409 <= not w14405 and not w14407;
w14410 <= not w14403 and w14409;
w14411 <= not w14408 and not w14410;
w14412 <= not w14400 and not w14411;
w14413 <= not w14400 and not w14412;
w14414 <= not w14411 and not w14412;
w14415 <= not w14413 and not w14414;
w14416 <= not w14370 and w14415;
w14417 <= w14370 and not w14415;
w14418 <= not w14416 and not w14417;
w14419 <= w14206 and w14242;
w14420 <= not w14206 and not w14242;
w14421 <= not w14419 and not w14420;
w14422 <= w14230 and not w14421;
w14423 <= not w14230 and w14421;
w14424 <= not w14422 and not w14423;
w14425 <= not w14093 and not w14096;
w14426 <= not w14099 and not w14102;
w14427 <= w14425 and w14426;
w14428 <= not w14425 and not w14426;
w14429 <= not w14427 and not w14428;
w14430 <= w14424 and w14429;
w14431 <= not w14424 and not w14429;
w14432 <= not w14430 and not w14431;
w14433 <= not w14418 and w14432;
w14434 <= not w14418 and not w14433;
w14435 <= w14432 and not w14433;
w14436 <= not w14434 and not w14435;
w14437 <= w14324 and not w14436;
w14438 <= not w14324 and w14436;
w14439 <= not w14294 and not w14438;
w14440 <= not w14437 and w14439;
w14441 <= not w14294 and not w14440;
w14442 <= not w14438 and not w14440;
w14443 <= not w14437 and w14442;
w14444 <= not w14441 and not w14443;
w14445 <= not w14269 and not w14272;
w14446 <= not w14088 and not w14111;
w14447 <= w14445 and w14446;
w14448 <= not w14445 and not w14446;
w14449 <= not w14447 and not w14448;
w14450 <= not w14218 and not w14267;
w14451 <= not w14106 and not w14108;
w14452 <= not w14450 and not w14451;
w14453 <= not w14450 and not w14452;
w14454 <= not w14451 and not w14452;
w14455 <= not w14453 and not w14454;
w14456 <= w14177 and w14192;
w14457 <= not w14177 and not w14192;
w14458 <= not w14456 and not w14457;
w14459 <= w14146 and not w14458;
w14460 <= not w14146 and w14458;
w14461 <= not w14459 and not w14460;
w14462 <= not w14248 and not w14262;
w14463 <= not w14195 and not w14212;
w14464 <= w14462 and w14463;
w14465 <= not w14462 and not w14463;
w14466 <= not w14464 and not w14465;
w14467 <= w14461 and w14466;
w14468 <= not w14461 and not w14466;
w14469 <= not w14467 and not w14468;
w14470 <= not w14455 and w14469;
w14471 <= not w14455 and not w14470;
w14472 <= w14469 and not w14470;
w14473 <= not w14471 and not w14472;
w14474 <= w14449 and not w14473;
w14475 <= not w14449 and w14473;
w14476 <= not w14444 and not w14475;
w14477 <= not w14474 and w14476;
w14478 <= not w14444 and not w14477;
w14479 <= not w14475 and not w14477;
w14480 <= not w14474 and w14479;
w14481 <= not w14478 and not w14480;
w14482 <= not w14292 and not w14481;
w14483 <= w14292 and w14481;
w14484 <= not w14482 and not w14483;
w14485 <= not w14291 and w14484;
w14486 <= w14291 and not w14484;
w14487 <= not w14485 and not w14486;
w14488 <= not w14291 and not w14483;
w14489 <= not w14482 and not w14488;
w14490 <= not w14440 and not w14477;
w14491 <= not w14448 and not w14474;
w14492 <= a(22) and a(63);
w14493 <= a(28) and a(57);
w14494 <= not w14492 and not w14493;
w14495 <= w14492 and w14493;
w14496 <= a(50) and not w14495;
w14497 <= a(35) and w14496;
w14498 <= not w14494 and w14497;
w14499 <= not w14495 and not w14498;
w14500 <= not w14494 and w14499;
w14501 <= a(50) and not w14498;
w14502 <= a(35) and w14501;
w14503 <= not w14500 and not w14502;
w14504 <= w3956 and w6774;
w14505 <= w3896 and w7038;
w14506 <= w2949 and w7239;
w14507 <= not w14505 and not w14506;
w14508 <= not w14504 and not w14507;
w14509 <= a(53) and not w14508;
w14510 <= a(32) and w14509;
w14511 <= not w14504 and not w14508;
w14512 <= a(33) and a(52);
w14513 <= a(34) and a(51);
w14514 <= not w14512 and not w14513;
w14515 <= w14511 and not w14514;
w14516 <= not w14510 and not w14515;
w14517 <= not w14503 and not w14516;
w14518 <= not w14503 and not w14517;
w14519 <= not w14516 and not w14517;
w14520 <= not w14518 and not w14519;
w14521 <= w5219 and w5519;
w14522 <= w3790 and w7553;
w14523 <= w3977 and w5366;
w14524 <= not w14522 and not w14523;
w14525 <= not w14521 and not w14524;
w14526 <= a(46) and not w14525;
w14527 <= a(39) and w14526;
w14528 <= not w14521 and not w14525;
w14529 <= a(40) and a(45);
w14530 <= a(41) and a(44);
w14531 <= not w14529 and not w14530;
w14532 <= w14528 and not w14531;
w14533 <= not w14527 and not w14532;
w14534 <= not w14520 and not w14533;
w14535 <= not w14520 and not w14534;
w14536 <= not w14533 and not w14534;
w14537 <= not w14535 and not w14536;
w14538 <= a(43) and a(62);
w14539 <= a(23) and w14538;
w14540 <= w4824 and not w14539;
w14541 <= not w14539 and not w14540;
w14542 <= a(23) and a(62);
w14543 <= not a(43) and not w14542;
w14544 <= w14541 and not w14543;
w14545 <= w4824 and not w14540;
w14546 <= not w14544 and not w14545;
w14547 <= w4371 and w6058;
w14548 <= w3336 and w6060;
w14549 <= w3493 and w6062;
w14550 <= not w14548 and not w14549;
w14551 <= not w14547 and not w14550;
w14552 <= a(49) and not w14551;
w14553 <= a(36) and w14552;
w14554 <= a(37) and a(48);
w14555 <= a(38) and a(47);
w14556 <= not w14554 and not w14555;
w14557 <= not w14547 and not w14551;
w14558 <= not w14556 and w14557;
w14559 <= not w14553 and not w14558;
w14560 <= not w14546 and not w14559;
w14561 <= not w14546 and not w14560;
w14562 <= not w14559 and not w14560;
w14563 <= not w14561 and not w14562;
w14564 <= w2671 and w7507;
w14565 <= w3258 and w7227;
w14566 <= w2423 and w8967;
w14567 <= not w14565 and not w14566;
w14568 <= not w14564 and not w14567;
w14569 <= a(56) and not w14568;
w14570 <= a(29) and w14569;
w14571 <= not w14564 and not w14568;
w14572 <= a(30) and a(55);
w14573 <= a(31) and a(54);
w14574 <= not w14572 and not w14573;
w14575 <= w14571 and not w14574;
w14576 <= not w14570 and not w14575;
w14577 <= not w14563 and not w14576;
w14578 <= not w14563 and not w14577;
w14579 <= not w14576 and not w14577;
w14580 <= not w14578 and not w14579;
w14581 <= not w14537 and w14580;
w14582 <= w14537 and not w14580;
w14583 <= not w14581 and not w14582;
w14584 <= not w14465 and not w14467;
w14585 <= w14583 and w14584;
w14586 <= not w14583 and not w14584;
w14587 <= not w14585 and not w14586;
w14588 <= not w14428 and not w14430;
w14589 <= a(24) and a(61);
w14590 <= not w14392 and w14589;
w14591 <= w14392 and not w14589;
w14592 <= not w14590 and not w14591;
w14593 <= w14380 and not w14592;
w14594 <= not w14380 and w14592;
w14595 <= not w14593 and not w14594;
w14596 <= w14306 and w14409;
w14597 <= not w14306 and not w14409;
w14598 <= not w14596 and not w14597;
w14599 <= w2033 and w8793;
w14600 <= w2439 and w9895;
w14601 <= w2269 and w9315;
w14602 <= not w14600 and not w14601;
w14603 <= not w14599 and not w14602;
w14604 <= a(60) and not w14603;
w14605 <= a(25) and w14604;
w14606 <= not w14599 and not w14603;
w14607 <= a(27) and a(58);
w14608 <= not w8117 and not w14607;
w14609 <= w14606 and not w14608;
w14610 <= not w14605 and not w14609;
w14611 <= w14598 and not w14610;
w14612 <= w14598 and not w14611;
w14613 <= not w14610 and not w14611;
w14614 <= not w14612 and not w14613;
w14615 <= w14595 and not w14614;
w14616 <= not w14595 and w14614;
w14617 <= not w14588 and not w14616;
w14618 <= not w14615 and w14617;
w14619 <= not w14588 and not w14618;
w14620 <= not w14615 and not w14618;
w14621 <= not w14616 and w14620;
w14622 <= not w14619 and not w14621;
w14623 <= w14330 and w14361;
w14624 <= not w14330 and not w14361;
w14625 <= not w14623 and not w14624;
w14626 <= w14347 and not w14625;
w14627 <= not w14347 and w14625;
w14628 <= not w14626 and not w14627;
w14629 <= not w14397 and not w14412;
w14630 <= not w14350 and not w14367;
w14631 <= w14629 and w14630;
w14632 <= not w14629 and not w14630;
w14633 <= not w14631 and not w14632;
w14634 <= w14628 and w14633;
w14635 <= not w14628 and not w14633;
w14636 <= not w14634 and not w14635;
w14637 <= not w14622 and w14636;
w14638 <= not w14622 and not w14637;
w14639 <= w14636 and not w14637;
w14640 <= not w14638 and not w14639;
w14641 <= w14587 and not w14640;
w14642 <= w14587 and not w14641;
w14643 <= not w14640 and not w14641;
w14644 <= not w14642 and not w14643;
w14645 <= not w14491 and not w14644;
w14646 <= not w14491 and not w14645;
w14647 <= not w14644 and not w14645;
w14648 <= not w14646 and not w14647;
w14649 <= not w14452 and not w14470;
w14650 <= not w14420 and not w14423;
w14651 <= not w14457 and not w14460;
w14652 <= w14650 and w14651;
w14653 <= not w14650 and not w14651;
w14654 <= not w14652 and not w14653;
w14655 <= not w14297 and not w14309;
w14656 <= not w14654 and w14655;
w14657 <= w14654 and not w14655;
w14658 <= not w14656 and not w14657;
w14659 <= not w14315 and not w14319;
w14660 <= not w14658 and w14659;
w14661 <= w14658 and not w14659;
w14662 <= not w14660 and not w14661;
w14663 <= not w14370 and not w14415;
w14664 <= not w14433 and not w14663;
w14665 <= w14662 and not w14664;
w14666 <= not w14662 and w14664;
w14667 <= not w14665 and not w14666;
w14668 <= w14649 and not w14667;
w14669 <= not w14649 and w14667;
w14670 <= not w14668 and not w14669;
w14671 <= not w14323 and not w14437;
w14672 <= w14670 and not w14671;
w14673 <= not w14670 and w14671;
w14674 <= not w14672 and not w14673;
w14675 <= not w14648 and not w14674;
w14676 <= w14648 and w14674;
w14677 <= not w14675 and not w14676;
w14678 <= not w14490 and not w14677;
w14679 <= w14490 and w14677;
w14680 <= not w14678 and not w14679;
w14681 <= not w14489 and not w14680;
w14682 <= w14489 and w14680;
w14683 <= not w14681 and not w14682;
w14684 <= not w14489 and not w14679;
w14685 <= not w14678 and not w14684;
w14686 <= not w14648 and w14674;
w14687 <= not w14645 and not w14686;
w14688 <= not w14669 and not w14672;
w14689 <= not w14597 and not w14611;
w14690 <= not w14517 and not w14534;
w14691 <= w14689 and w14690;
w14692 <= not w14689 and not w14690;
w14693 <= not w14691 and not w14692;
w14694 <= not w14560 and not w14577;
w14695 <= not w14693 and w14694;
w14696 <= w14693 and not w14694;
w14697 <= not w14695 and not w14696;
w14698 <= not w14653 and not w14657;
w14699 <= w14528 and w14571;
w14700 <= not w14528 and not w14571;
w14701 <= not w14699 and not w14700;
w14702 <= w14557 and not w14701;
w14703 <= not w14557 and w14701;
w14704 <= not w14702 and not w14703;
w14705 <= w14511 and w14606;
w14706 <= not w14511 and not w14606;
w14707 <= not w14705 and not w14706;
w14708 <= w14499 and not w14707;
w14709 <= not w14499 and w14707;
w14710 <= not w14708 and not w14709;
w14711 <= w14704 and w14710;
w14712 <= not w14704 and not w14710;
w14713 <= not w14711 and not w14712;
w14714 <= not w14698 and w14713;
w14715 <= w14698 and not w14713;
w14716 <= not w14714 and not w14715;
w14717 <= w14697 and w14716;
w14718 <= not w14697 and not w14716;
w14719 <= not w14717 and not w14718;
w14720 <= not w14632 and not w14634;
w14721 <= a(36) and a(50);
w14722 <= a(37) and a(49);
w14723 <= not w14721 and not w14722;
w14724 <= w3493 and w6131;
w14725 <= a(63) and not w14724;
w14726 <= not w14723 and w14725;
w14727 <= a(23) and w14726;
w14728 <= not w14724 and not w14727;
w14729 <= not w14723 and w14728;
w14730 <= a(63) and not w14727;
w14731 <= a(23) and w14730;
w14732 <= not w14729 and not w14731;
w14733 <= w3125 and w6774;
w14734 <= w2778 and w7038;
w14735 <= w3956 and w7239;
w14736 <= not w14734 and not w14735;
w14737 <= not w14733 and not w14736;
w14738 <= a(53) and not w14737;
w14739 <= a(33) and w14738;
w14740 <= not w14733 and not w14737;
w14741 <= a(34) and a(52);
w14742 <= a(35) and a(51);
w14743 <= not w14741 and not w14742;
w14744 <= w14740 and not w14743;
w14745 <= not w14739 and not w14744;
w14746 <= not w14732 and not w14745;
w14747 <= not w14732 and not w14746;
w14748 <= not w14745 and not w14746;
w14749 <= not w14747 and not w14748;
w14750 <= not w12129 and not w14137;
w14751 <= w3258 and w11524;
w14752 <= w6748 and not w14751;
w14753 <= not w14750 and w14752;
w14754 <= w6748 and not w14753;
w14755 <= not w14751 and not w14753;
w14756 <= not w14750 and w14755;
w14757 <= not w14754 and not w14756;
w14758 <= not w14749 and not w14757;
w14759 <= not w14749 and not w14758;
w14760 <= not w14757 and not w14758;
w14761 <= not w14759 and not w14760;
w14762 <= w2137 and w8793;
w14763 <= w2606 and w9895;
w14764 <= w2033 and w9315;
w14765 <= not w14763 and not w14764;
w14766 <= not w14762 and not w14765;
w14767 <= not w14762 and not w14766;
w14768 <= a(27) and a(59);
w14769 <= a(28) and a(58);
w14770 <= not w14768 and not w14769;
w14771 <= w14767 and not w14770;
w14772 <= a(60) and not w14766;
w14773 <= a(26) and w14772;
w14774 <= not w14771 and not w14773;
w14775 <= a(32) and a(54);
w14776 <= w4445 and w14775;
w14777 <= w4615 and w14775;
w14778 <= w5150 and w5519;
w14779 <= not w14777 and not w14778;
w14780 <= not w14776 and not w14779;
w14781 <= w4615 and not w14780;
w14782 <= not w14776 and not w14780;
w14783 <= not w4445 and not w14775;
w14784 <= w14782 and not w14783;
w14785 <= not w14781 and not w14784;
w14786 <= not w14774 and not w14785;
w14787 <= not w14774 and not w14786;
w14788 <= not w14785 and not w14786;
w14789 <= not w14787 and not w14788;
w14790 <= a(39) and a(47);
w14791 <= not w6879 and not w14790;
w14792 <= w3977 and w5472;
w14793 <= a(56) and not w14792;
w14794 <= a(30) and w14793;
w14795 <= not w14791 and w14794;
w14796 <= a(56) and not w14795;
w14797 <= a(30) and w14796;
w14798 <= not w14792 and not w14795;
w14799 <= not w14791 and w14798;
w14800 <= not w14797 and not w14799;
w14801 <= not w14789 and not w14800;
w14802 <= not w14789 and not w14801;
w14803 <= not w14800 and not w14801;
w14804 <= not w14802 and not w14803;
w14805 <= w14761 and w14804;
w14806 <= not w14761 and not w14804;
w14807 <= not w14805 and not w14806;
w14808 <= not w14720 and w14807;
w14809 <= w14720 and not w14807;
w14810 <= not w14808 and not w14809;
w14811 <= w14719 and w14810;
w14812 <= not w14719 and not w14810;
w14813 <= not w14811 and not w14812;
w14814 <= not w14688 and w14813;
w14815 <= not w14688 and not w14814;
w14816 <= w14813 and not w14814;
w14817 <= not w14815 and not w14816;
w14818 <= not w14637 and not w14641;
w14819 <= not w14661 and not w14665;
w14820 <= w14818 and w14819;
w14821 <= not w14818 and not w14819;
w14822 <= not w14820 and not w14821;
w14823 <= w1710 and w9527;
w14824 <= a(61) and not w14823;
w14825 <= a(25) and w14824;
w14826 <= a(62) and not w14823;
w14827 <= a(24) and w14826;
w14828 <= not w14825 and not w14827;
w14829 <= not w14541 and not w14828;
w14830 <= not w14541 and not w14829;
w14831 <= not w14828 and not w14829;
w14832 <= not w14830 and not w14831;
w14833 <= not w14590 and not w14594;
w14834 <= w14832 and w14833;
w14835 <= not w14832 and not w14833;
w14836 <= not w14834 and not w14835;
w14837 <= not w14624 and not w14627;
w14838 <= not w14836 and w14837;
w14839 <= w14836 and not w14837;
w14840 <= not w14838 and not w14839;
w14841 <= not w14620 and w14840;
w14842 <= w14620 and not w14840;
w14843 <= not w14841 and not w14842;
w14844 <= not w14537 and not w14580;
w14845 <= not w14586 and not w14844;
w14846 <= w14843 and not w14845;
w14847 <= not w14843 and w14845;
w14848 <= not w14846 and not w14847;
w14849 <= w14822 and w14848;
w14850 <= not w14822 and not w14848;
w14851 <= not w14849 and not w14850;
w14852 <= not w14817 and w14851;
w14853 <= not w14816 and not w14851;
w14854 <= not w14815 and w14853;
w14855 <= not w14852 and not w14854;
w14856 <= w14687 and not w14855;
w14857 <= not w14687 and w14855;
w14858 <= not w14856 and not w14857;
w14859 <= w14685 and not w14858;
w14860 <= not w14685 and not w14856;
w14861 <= not w14857 and w14860;
w14862 <= not w14859 and not w14861;
w14863 <= not w14857 and not w14860;
w14864 <= not w14814 and not w14852;
w14865 <= not w14806 and not w14808;
w14866 <= not w14700 and not w14703;
w14867 <= not w14746 and not w14758;
w14868 <= w14866 and w14867;
w14869 <= not w14866 and not w14867;
w14870 <= not w14868 and not w14869;
w14871 <= not w14786 and not w14801;
w14872 <= not w14870 and w14871;
w14873 <= w14870 and not w14871;
w14874 <= not w14872 and not w14873;
w14875 <= not w14865 and w14874;
w14876 <= w14865 and not w14874;
w14877 <= not w14875 and not w14876;
w14878 <= not w14841 and not w14846;
w14879 <= not w14877 and w14878;
w14880 <= w14877 and not w14878;
w14881 <= not w14879 and not w14880;
w14882 <= not w14821 and not w14849;
w14883 <= not w14881 and w14882;
w14884 <= w14881 and not w14882;
w14885 <= not w14883 and not w14884;
w14886 <= not w14711 and not w14714;
w14887 <= not w14692 and not w14696;
w14888 <= w14886 and w14887;
w14889 <= not w14886 and not w14887;
w14890 <= not w14888 and not w14889;
w14891 <= not w14835 and not w14839;
w14892 <= w14782 and w14798;
w14893 <= not w14782 and not w14798;
w14894 <= not w14892 and not w14893;
w14895 <= w14755 and not w14894;
w14896 <= not w14755 and w14894;
w14897 <= not w14895 and not w14896;
w14898 <= w14740 and w14767;
w14899 <= not w14740 and not w14767;
w14900 <= not w14898 and not w14899;
w14901 <= w14728 and not w14900;
w14902 <= not w14728 and w14900;
w14903 <= not w14901 and not w14902;
w14904 <= not w14897 and not w14903;
w14905 <= w14897 and w14903;
w14906 <= not w14904 and not w14905;
w14907 <= not w14891 and w14906;
w14908 <= w14891 and not w14906;
w14909 <= not w14907 and not w14908;
w14910 <= w14890 and w14909;
w14911 <= not w14890 and not w14909;
w14912 <= not w14717 and not w14811;
w14913 <= a(44) and a(62);
w14914 <= a(25) and w14913;
w14915 <= w5102 and not w14914;
w14916 <= not w14914 and not w14915;
w14917 <= a(25) and a(62);
w14918 <= not a(44) and not w14917;
w14919 <= w14916 and not w14918;
w14920 <= w5102 and not w14915;
w14921 <= not w14919 and not w14920;
w14922 <= a(31) and a(56);
w14923 <= a(33) and a(54);
w14924 <= not w14922 and not w14923;
w14925 <= w2404 and w7227;
w14926 <= a(47) and not w14925;
w14927 <= a(40) and w14926;
w14928 <= not w14924 and w14927;
w14929 <= a(47) and not w14928;
w14930 <= a(40) and w14929;
w14931 <= not w14925 and not w14928;
w14932 <= not w14924 and w14931;
w14933 <= not w14930 and not w14932;
w14934 <= not w14921 and not w14933;
w14935 <= not w14921 and not w14934;
w14936 <= not w14933 and not w14934;
w14937 <= not w14935 and not w14936;
w14938 <= not w14706 and not w14709;
w14939 <= w14937 and w14938;
w14940 <= not w14937 and not w14938;
w14941 <= not w14939 and not w14940;
w14942 <= w2033 and w9318;
w14943 <= w2107 and w9715;
w14944 <= w6002 and w11440;
w14945 <= not w14943 and not w14944;
w14946 <= not w14942 and not w14945;
w14947 <= not w14942 and not w14946;
w14948 <= a(26) and a(61);
w14949 <= a(27) and a(60);
w14950 <= not w14948 and not w14949;
w14951 <= w14947 and not w14950;
w14952 <= a(63) and not w14946;
w14953 <= a(24) and w14952;
w14954 <= not w14951 and not w14953;
w14955 <= w4889 and w6062;
w14956 <= w5236 and w5694;
w14957 <= w4371 and w6131;
w14958 <= not w14956 and not w14957;
w14959 <= not w14955 and not w14958;
w14960 <= a(50) and not w14959;
w14961 <= a(37) and w14960;
w14962 <= a(38) and a(49);
w14963 <= a(39) and a(48);
w14964 <= not w14962 and not w14963;
w14965 <= not w14955 and not w14959;
w14966 <= not w14964 and w14965;
w14967 <= not w14961 and not w14966;
w14968 <= not w14954 and not w14967;
w14969 <= not w14954 and not w14968;
w14970 <= not w14967 and not w14968;
w14971 <= not w14969 and not w14970;
w14972 <= a(41) and a(46);
w14973 <= a(42) and a(45);
w14974 <= not w14972 and not w14973;
w14975 <= w5150 and w5366;
w14976 <= a(55) and not w14975;
w14977 <= a(32) and w14976;
w14978 <= not w14974 and w14977;
w14979 <= a(55) and not w14978;
w14980 <= a(32) and w14979;
w14981 <= not w14975 and not w14978;
w14982 <= not w14974 and w14981;
w14983 <= not w14980 and not w14982;
w14984 <= not w14971 and not w14983;
w14985 <= not w14971 and not w14984;
w14986 <= not w14983 and not w14984;
w14987 <= not w14985 and not w14986;
w14988 <= not w14941 and w14987;
w14989 <= w14941 and not w14987;
w14990 <= not w14988 and not w14989;
w14991 <= a(34) and a(53);
w14992 <= w14404 and w14991;
w14993 <= w2916 and w8791;
w14994 <= a(34) and a(59);
w14995 <= w13748 and w14994;
w14996 <= not w14993 and not w14995;
w14997 <= not w14992 and not w14996;
w14998 <= a(59) and not w14997;
w14999 <= a(28) and w14998;
w15000 <= not w14992 and not w14997;
w15001 <= not w14404 and not w14991;
w15002 <= w15000 and not w15001;
w15003 <= not w14999 and not w15002;
w15004 <= not w14823 and not w14829;
w15005 <= not w15003 and w15004;
w15006 <= w15003 and not w15004;
w15007 <= not w15005 and not w15006;
w15008 <= w3634 and w6774;
w15009 <= a(35) and a(58);
w15010 <= w13749 and w15009;
w15011 <= not w15008 and not w15010;
w15012 <= a(29) and a(58);
w15013 <= a(36) and a(51);
w15014 <= w15012 and w15013;
w15015 <= not w15011 and not w15014;
w15016 <= a(52) and not w15015;
w15017 <= a(35) and w15016;
w15018 <= not w15014 and not w15015;
w15019 <= not w15012 and not w15013;
w15020 <= w15018 and not w15019;
w15021 <= not w15017 and not w15020;
w15022 <= not w15007 and not w15021;
w15023 <= w15007 and w15021;
w15024 <= not w15022 and not w15023;
w15025 <= w14990 and w15024;
w15026 <= not w14990 and not w15024;
w15027 <= not w15025 and not w15026;
w15028 <= not w14912 and w15027;
w15029 <= w14912 and not w15027;
w15030 <= not w15028 and not w15029;
w15031 <= not w14911 and w15030;
w15032 <= not w14910 and w15031;
w15033 <= w15030 and not w15032;
w15034 <= not w14911 and not w15032;
w15035 <= not w14910 and w15034;
w15036 <= not w15033 and not w15035;
w15037 <= not w14885 and w15036;
w15038 <= w14885 and not w15036;
w15039 <= not w15037 and not w15038;
w15040 <= w14864 and not w15039;
w15041 <= not w14864 and w15039;
w15042 <= not w15040 and not w15041;
w15043 <= not w14863 and not w15042;
w15044 <= w14863 and w15042;
w15045 <= not w15043 and not w15044;
w15046 <= not w14884 and not w15038;
w15047 <= not w14875 and not w14880;
w15048 <= w2137 and w9318;
w15049 <= w2606 and w8891;
w15050 <= w2033 and w9527;
w15051 <= not w15049 and not w15050;
w15052 <= not w15048 and not w15051;
w15053 <= not w15048 and not w15052;
w15054 <= a(27) and a(61);
w15055 <= a(28) and a(60);
w15056 <= not w15054 and not w15055;
w15057 <= w15053 and not w15056;
w15058 <= a(62) and not w15052;
w15059 <= a(26) and w15058;
w15060 <= not w15057 and not w15059;
w15061 <= a(42) and a(46);
w15062 <= a(41) and a(47);
w15063 <= not w15061 and not w15062;
w15064 <= w5150 and w5472;
w15065 <= a(31) and not w15064;
w15066 <= a(57) and w15065;
w15067 <= not w15063 and w15066;
w15068 <= a(57) and not w15067;
w15069 <= a(31) and w15068;
w15070 <= not w15064 and not w15067;
w15071 <= not w15063 and w15070;
w15072 <= not w15069 and not w15071;
w15073 <= not w15060 and not w15072;
w15074 <= not w15060 and not w15073;
w15075 <= not w15072 and not w15073;
w15076 <= not w15074 and not w15075;
w15077 <= w3493 and w6774;
w15078 <= w4837 and w7038;
w15079 <= w3634 and w7239;
w15080 <= not w15078 and not w15079;
w15081 <= not w15077 and not w15080;
w15082 <= a(53) and not w15081;
w15083 <= a(35) and w15082;
w15084 <= not w15077 and not w15081;
w15085 <= a(37) and a(51);
w15086 <= a(36) and a(52);
w15087 <= not w15085 and not w15086;
w15088 <= w15084 and not w15087;
w15089 <= not w15083 and not w15088;
w15090 <= not w15076 and not w15089;
w15091 <= not w15076 and not w15090;
w15092 <= not w15089 and not w15090;
w15093 <= not w15091 and not w15092;
w15094 <= a(38) and a(50);
w15095 <= a(39) and a(49);
w15096 <= not w15094 and not w15095;
w15097 <= w4889 and w6131;
w15098 <= a(29) and not w15097;
w15099 <= a(59) and w15098;
w15100 <= not w15096 and w15099;
w15101 <= not w15097 and not w15100;
w15102 <= not w15096 and w15101;
w15103 <= a(59) and not w15100;
w15104 <= a(29) and w15103;
w15105 <= not w15102 and not w15104;
w15106 <= a(30) and a(58);
w15107 <= a(32) and a(56);
w15108 <= not w15106 and not w15107;
w15109 <= w2294 and w7748;
w15110 <= w7159 and not w15109;
w15111 <= not w15108 and w15110;
w15112 <= w7159 and not w15111;
w15113 <= not w15109 and not w15111;
w15114 <= not w15108 and w15113;
w15115 <= not w15112 and not w15114;
w15116 <= not w15105 and not w15115;
w15117 <= not w15105 and not w15116;
w15118 <= not w15115 and not w15116;
w15119 <= not w15117 and not w15118;
w15120 <= not w14893 and not w14896;
w15121 <= w15119 and w15120;
w15122 <= not w15119 and not w15120;
w15123 <= not w15121 and not w15122;
w15124 <= a(25) and a(63);
w15125 <= not w14916 and w15124;
w15126 <= w14916 and not w15124;
w15127 <= not w15125 and not w15126;
w15128 <= w14981 and not w15127;
w15129 <= not w14981 and w15127;
w15130 <= not w15128 and not w15129;
w15131 <= w15123 and w15130;
w15132 <= not w15123 and not w15130;
w15133 <= not w15131 and not w15132;
w15134 <= not w15093 and w15133;
w15135 <= not w15093 and not w15134;
w15136 <= w15133 and not w15134;
w15137 <= not w15135 and not w15136;
w15138 <= not w15047 and not w15137;
w15139 <= not w15047 and not w15138;
w15140 <= not w15137 and not w15138;
w15141 <= not w15139 and not w15140;
w15142 <= not w14905 and not w14907;
w15143 <= not w14869 and not w14873;
w15144 <= w15142 and w15143;
w15145 <= not w15142 and not w15143;
w15146 <= not w15144 and not w15145;
w15147 <= w14947 and w15000;
w15148 <= not w14947 and not w15000;
w15149 <= not w15147 and not w15148;
w15150 <= w14965 and not w15149;
w15151 <= not w14965 and w15149;
w15152 <= not w15150 and not w15151;
w15153 <= w14931 and w15018;
w15154 <= not w14931 and not w15018;
w15155 <= not w15153 and not w15154;
w15156 <= a(33) and a(55);
w15157 <= a(34) and a(54);
w15158 <= not w15156 and not w15157;
w15159 <= w3956 and w7507;
w15160 <= w4617 and not w15159;
w15161 <= not w15158 and w15160;
w15162 <= w4617 and not w15161;
w15163 <= not w15159 and not w15161;
w15164 <= not w15158 and w15163;
w15165 <= not w15162 and not w15164;
w15166 <= w15155 and not w15165;
w15167 <= w15155 and not w15166;
w15168 <= not w15165 and not w15166;
w15169 <= not w15167 and not w15168;
w15170 <= not w14934 and not w14940;
w15171 <= w15169 and w15170;
w15172 <= not w15169 and not w15170;
w15173 <= not w15171 and not w15172;
w15174 <= w15152 and w15173;
w15175 <= not w15152 and not w15173;
w15176 <= not w15174 and not w15175;
w15177 <= w15146 and w15176;
w15178 <= not w15146 and not w15176;
w15179 <= not w15177 and not w15178;
w15180 <= not w15141 and not w15179;
w15181 <= w15141 and w15179;
w15182 <= not w15180 and not w15181;
w15183 <= not w15028 and not w15032;
w15184 <= not w14889 and not w14910;
w15185 <= not w14899 and not w14902;
w15186 <= not w15003 and not w15004;
w15187 <= not w15022 and not w15186;
w15188 <= w15185 and w15187;
w15189 <= not w15185 and not w15187;
w15190 <= not w15188 and not w15189;
w15191 <= not w14968 and not w14984;
w15192 <= not w15190 and w15191;
w15193 <= w15190 and not w15191;
w15194 <= not w15192 and not w15193;
w15195 <= not w14989 and not w15025;
w15196 <= w15194 and not w15195;
w15197 <= not w15194 and w15195;
w15198 <= not w15196 and not w15197;
w15199 <= not w15184 and w15198;
w15200 <= w15184 and not w15198;
w15201 <= not w15199 and not w15200;
w15202 <= not w15183 and w15201;
w15203 <= w15183 and not w15201;
w15204 <= not w15202 and not w15203;
w15205 <= not w15182 and w15204;
w15206 <= w15204 and not w15205;
w15207 <= not w15182 and not w15205;
w15208 <= not w15206 and not w15207;
w15209 <= w15046 and w15208;
w15210 <= not w15046 and not w15208;
w15211 <= not w15209 and not w15210;
w15212 <= not w14863 and not w15040;
w15213 <= not w15041 and not w15212;
w15214 <= not w15211 and w15213;
w15215 <= w15211 and not w15213;
w15216 <= not w15214 and not w15215;
w15217 <= not w15202 and not w15205;
w15218 <= not w15196 and not w15199;
w15219 <= a(33) and a(56);
w15220 <= a(35) and a(54);
w15221 <= not w15219 and not w15220;
w15222 <= w2778 and w7227;
w15223 <= a(48) and not w15222;
w15224 <= a(41) and w15223;
w15225 <= not w15221 and w15224;
w15226 <= not w15222 and not w15225;
w15227 <= not w15221 and w15226;
w15228 <= a(48) and not w15225;
w15229 <= a(41) and w15228;
w15230 <= not w15227 and not w15229;
w15231 <= w4371 and w6774;
w15232 <= w3336 and w7038;
w15233 <= w3493 and w7239;
w15234 <= not w15232 and not w15233;
w15235 <= not w15231 and not w15234;
w15236 <= a(53) and not w15235;
w15237 <= a(36) and w15236;
w15238 <= not w15231 and not w15235;
w15239 <= not w7342 and not w10362;
w15240 <= w15238 and not w15239;
w15241 <= not w15237 and not w15240;
w15242 <= not w15230 and not w15241;
w15243 <= not w15230 and not w15242;
w15244 <= not w15241 and not w15242;
w15245 <= not w15243 and not w15244;
w15246 <= w3618 and w8242;
w15247 <= w2294 and w8791;
w15248 <= w2671 and w8793;
w15249 <= not w15247 and not w15248;
w15250 <= not w15246 and not w15249;
w15251 <= a(59) and not w15250;
w15252 <= a(30) and w15251;
w15253 <= not w15246 and not w15250;
w15254 <= a(31) and a(58);
w15255 <= a(32) and a(57);
w15256 <= not w15254 and not w15255;
w15257 <= w15253 and not w15256;
w15258 <= not w15252 and not w15257;
w15259 <= not w15245 and not w15258;
w15260 <= not w15245 and not w15259;
w15261 <= not w15258 and not w15259;
w15262 <= not w15260 and not w15261;
w15263 <= w15053 and w15084;
w15264 <= not w15053 and not w15084;
w15265 <= not w15263 and not w15264;
w15266 <= w15113 and not w15265;
w15267 <= not w15113 and w15265;
w15268 <= not w15266 and not w15267;
w15269 <= a(45) and a(62);
w15270 <= a(27) and w15269;
w15271 <= w5519 and not w15270;
w15272 <= not w15270 and not w15271;
w15273 <= a(27) and a(62);
w15274 <= not a(45) and not w15273;
w15275 <= w15272 and not w15274;
w15276 <= w5519 and not w15271;
w15277 <= not w15275 and not w15276;
w15278 <= a(34) and a(55);
w15279 <= a(42) and a(47);
w15280 <= a(43) and a(46);
w15281 <= not w15279 and not w15280;
w15282 <= w4824 and w5472;
w15283 <= w15278 and not w15282;
w15284 <= not w15281 and w15283;
w15285 <= w15278 and not w15284;
w15286 <= not w15282 and not w15284;
w15287 <= not w15281 and w15286;
w15288 <= not w15285 and not w15287;
w15289 <= not w15277 and not w15288;
w15290 <= not w15277 and not w15289;
w15291 <= not w15288 and not w15289;
w15292 <= not w15290 and not w15291;
w15293 <= w2140 and w9318;
w15294 <= a(60) and not w15293;
w15295 <= a(29) and w15294;
w15296 <= a(61) and not w15293;
w15297 <= a(28) and w15296;
w15298 <= not w15295 and not w15297;
w15299 <= not w15163 and not w15298;
w15300 <= not w15163 and not w15299;
w15301 <= not w15298 and not w15299;
w15302 <= not w15300 and not w15301;
w15303 <= not w15292 and w15302;
w15304 <= w15292 and not w15302;
w15305 <= not w15303 and not w15304;
w15306 <= w15268 and not w15305;
w15307 <= w15268 and not w15306;
w15308 <= not w15305 and not w15306;
w15309 <= not w15307 and not w15308;
w15310 <= not w15262 and not w15309;
w15311 <= not w15262 and not w15310;
w15312 <= not w15309 and not w15310;
w15313 <= not w15311 and not w15312;
w15314 <= not w15218 and not w15313;
w15315 <= not w15218 and not w15314;
w15316 <= not w15313 and not w15314;
w15317 <= not w15315 and not w15316;
w15318 <= not w15148 and not w15151;
w15319 <= not w15125 and not w15129;
w15320 <= w15318 and w15319;
w15321 <= not w15318 and not w15319;
w15322 <= not w15320 and not w15321;
w15323 <= not w15154 and not w15166;
w15324 <= not w15322 and w15323;
w15325 <= w15322 and not w15323;
w15326 <= not w15324 and not w15325;
w15327 <= not w15189 and not w15193;
w15328 <= not w15326 and w15327;
w15329 <= w15326 and not w15327;
w15330 <= not w15328 and not w15329;
w15331 <= not w15172 and not w15174;
w15332 <= w15330 and not w15331;
w15333 <= not w15330 and w15331;
w15334 <= not w15332 and not w15333;
w15335 <= not w15317 and w15334;
w15336 <= not w15317 and not w15335;
w15337 <= w15334 and not w15335;
w15338 <= not w15336 and not w15337;
w15339 <= not w15141 and w15179;
w15340 <= not w15138 and not w15339;
w15341 <= not w15145 and not w15177;
w15342 <= not w15131 and not w15134;
w15343 <= not w15116 and not w15122;
w15344 <= not w15073 and not w15090;
w15345 <= w15343 and w15344;
w15346 <= not w15343 and not w15344;
w15347 <= not w15345 and not w15346;
w15348 <= w15070 and w15101;
w15349 <= not w15070 and not w15101;
w15350 <= not w15348 and not w15349;
w15351 <= a(39) and a(50);
w15352 <= a(40) and a(49);
w15353 <= not w15351 and not w15352;
w15354 <= w3977 and w6131;
w15355 <= a(63) and not w15354;
w15356 <= not w15353 and w15355;
w15357 <= a(26) and w15356;
w15358 <= a(63) and not w15357;
w15359 <= a(26) and w15358;
w15360 <= not w15354 and not w15357;
w15361 <= not w15353 and w15360;
w15362 <= not w15359 and not w15361;
w15363 <= w15350 and not w15362;
w15364 <= w15350 and not w15363;
w15365 <= not w15362 and not w15363;
w15366 <= not w15364 and not w15365;
w15367 <= not w15347 and w15366;
w15368 <= w15347 and not w15366;
w15369 <= not w15367 and not w15368;
w15370 <= not w15342 and w15369;
w15371 <= w15342 and not w15369;
w15372 <= not w15370 and not w15371;
w15373 <= not w15341 and w15372;
w15374 <= w15341 and not w15372;
w15375 <= not w15373 and not w15374;
w15376 <= not w15340 and w15375;
w15377 <= w15375 and not w15376;
w15378 <= not w15340 and not w15376;
w15379 <= not w15377 and not w15378;
w15380 <= not w15338 and not w15379;
w15381 <= w15338 and not w15378;
w15382 <= not w15377 and w15381;
w15383 <= not w15380 and not w15382;
w15384 <= not w15217 and w15383;
w15385 <= w15217 and not w15383;
w15386 <= not w15384 and not w15385;
w15387 <= not w15209 and not w15213;
w15388 <= not w15210 and not w15387;
w15389 <= not w15386 and w15388;
w15390 <= w15386 and not w15388;
w15391 <= not w15389 and not w15390;
w15392 <= not w15385 and not w15388;
w15393 <= not w15384 and not w15392;
w15394 <= not w15376 and not w15380;
w15395 <= not w15329 and not w15332;
w15396 <= not w15306 and not w15310;
w15397 <= w15272 and w15286;
w15398 <= not w15272 and not w15286;
w15399 <= not w15397 and not w15398;
w15400 <= w15226 and not w15399;
w15401 <= not w15226 and w15399;
w15402 <= not w15400 and not w15401;
w15403 <= not w15292 and not w15302;
w15404 <= not w15289 and not w15403;
w15405 <= not w15242 and not w15259;
w15406 <= w15404 and w15405;
w15407 <= not w15404 and not w15405;
w15408 <= not w15406 and not w15407;
w15409 <= w15402 and w15408;
w15410 <= not w15402 and not w15408;
w15411 <= not w15409 and not w15410;
w15412 <= not w15396 and w15411;
w15413 <= w15396 and not w15411;
w15414 <= not w15412 and not w15413;
w15415 <= w15395 and not w15414;
w15416 <= not w15395 and w15414;
w15417 <= not w15415 and not w15416;
w15418 <= not w15314 and not w15335;
w15419 <= not w15417 and w15418;
w15420 <= w15417 and not w15418;
w15421 <= not w15419 and not w15420;
w15422 <= not w15370 and not w15373;
w15423 <= w15238 and w15253;
w15424 <= not w15238 and not w15253;
w15425 <= not w15423 and not w15424;
w15426 <= w15360 and not w15425;
w15427 <= not w15360 and w15425;
w15428 <= not w15426 and not w15427;
w15429 <= not w15321 and not w15325;
w15430 <= not w15428 and w15429;
w15431 <= w15428 and not w15429;
w15432 <= not w15430 and not w15431;
w15433 <= a(33) and a(57);
w15434 <= a(34) and a(56);
w15435 <= not w15433 and not w15434;
w15436 <= w3956 and w8006;
w15437 <= w2778 and w11524;
w15438 <= w3125 and w8967;
w15439 <= not w15437 and not w15438;
w15440 <= not w15436 and not w15439;
w15441 <= not w15436 and not w15440;
w15442 <= not w15435 and w15441;
w15443 <= a(55) and not w15440;
w15444 <= a(35) and w15443;
w15445 <= not w15442 and not w15444;
w15446 <= w4371 and w7239;
w15447 <= w3336 and w10711;
w15448 <= w3493 and w7505;
w15449 <= not w15447 and not w15448;
w15450 <= not w15446 and not w15449;
w15451 <= a(54) and not w15450;
w15452 <= a(36) and w15451;
w15453 <= not w15446 and not w15450;
w15454 <= a(38) and a(52);
w15455 <= not w7241 and not w15454;
w15456 <= w15453 and not w15455;
w15457 <= not w15452 and not w15456;
w15458 <= not w15445 and not w15457;
w15459 <= not w15445 and not w15458;
w15460 <= not w15457 and not w15458;
w15461 <= not w15459 and not w15460;
w15462 <= w5102 and w5472;
w15463 <= w4445 and w8384;
w15464 <= w4824 and w6058;
w15465 <= not w15463 and not w15464;
w15466 <= not w15462 and not w15465;
w15467 <= a(48) and not w15466;
w15468 <= a(42) and w15467;
w15469 <= not w15462 and not w15466;
w15470 <= not w7553 and not w7859;
w15471 <= w15469 and not w15470;
w15472 <= not w15468 and not w15471;
w15473 <= not w15461 and not w15472;
w15474 <= not w15461 and not w15473;
w15475 <= not w15472 and not w15473;
w15476 <= not w15474 and not w15475;
w15477 <= w15432 and not w15476;
w15478 <= not w15432 and w15476;
w15479 <= not w15422 and not w15478;
w15480 <= not w15477 and w15479;
w15481 <= not w15422 and not w15480;
w15482 <= not w15478 and not w15480;
w15483 <= not w15477 and w15482;
w15484 <= not w15481 and not w15483;
w15485 <= not w15346 and not w15368;
w15486 <= not w15264 and not w15267;
w15487 <= w5219 and w6131;
w15488 <= w3790 and w9740;
w15489 <= w3977 and w6370;
w15490 <= not w15488 and not w15489;
w15491 <= not w15487 and not w15490;
w15492 <= w7580 and not w15491;
w15493 <= not w15487 and not w15491;
w15494 <= a(41) and a(49);
w15495 <= a(40) and a(50);
w15496 <= not w15494 and not w15495;
w15497 <= w15493 and not w15496;
w15498 <= not w15492 and not w15497;
w15499 <= not w15486 and not w15498;
w15500 <= not w15486 and not w15499;
w15501 <= not w15498 and not w15499;
w15502 <= not w15500 and not w15501;
w15503 <= not w15349 and not w15363;
w15504 <= w15502 and w15503;
w15505 <= not w15502 and not w15503;
w15506 <= not w15504 and not w15505;
w15507 <= w2140 and w9527;
w15508 <= w2137 and w9598;
w15509 <= w1847 and w9715;
w15510 <= not w15508 and not w15509;
w15511 <= not w15507 and not w15510;
w15512 <= not w15507 and not w15511;
w15513 <= a(28) and a(62);
w15514 <= a(29) and a(61);
w15515 <= not w15513 and not w15514;
w15516 <= w15512 and not w15515;
w15517 <= a(63) and not w15511;
w15518 <= a(27) and w15517;
w15519 <= not w15516 and not w15518;
w15520 <= not w15293 and not w15299;
w15521 <= w3618 and w8793;
w15522 <= w2294 and w9895;
w15523 <= w2671 and w9315;
w15524 <= not w15522 and not w15523;
w15525 <= not w15521 and not w15524;
w15526 <= a(31) and a(59);
w15527 <= not w14226 and not w15526;
w15528 <= not w15521 and not w15527;
w15529 <= a(30) and a(60);
w15530 <= not w15528 and not w15529;
w15531 <= not w15525 and not w15530;
w15532 <= not w15520 and w15531;
w15533 <= not w15520 and not w15532;
w15534 <= w15531 and not w15532;
w15535 <= not w15533 and not w15534;
w15536 <= not w15519 and not w15535;
w15537 <= w15519 and not w15534;
w15538 <= not w15533 and w15537;
w15539 <= not w15536 and not w15538;
w15540 <= w15506 and w15539;
w15541 <= w15506 and not w15540;
w15542 <= w15539 and not w15540;
w15543 <= not w15541 and not w15542;
w15544 <= not w15485 and not w15543;
w15545 <= not w15485 and not w15544;
w15546 <= not w15543 and not w15544;
w15547 <= not w15545 and not w15546;
w15548 <= not w15484 and not w15547;
w15549 <= not w15484 and not w15548;
w15550 <= not w15547 and not w15548;
w15551 <= not w15549 and not w15550;
w15552 <= not w15421 and w15551;
w15553 <= w15421 and not w15551;
w15554 <= not w15552 and not w15553;
w15555 <= w15394 and not w15554;
w15556 <= not w15394 and w15554;
w15557 <= not w15555 and not w15556;
w15558 <= w15393 and not w15557;
w15559 <= not w15393 and not w15555;
w15560 <= not w15556 and w15559;
w15561 <= not w15558 and not w15560;
w15562 <= not w15556 and not w15559;
w15563 <= not w15420 and not w15553;
w15564 <= not w15398 and not w15401;
w15565 <= a(34) and a(57);
w15566 <= a(36) and a(55);
w15567 <= not w15565 and not w15566;
w15568 <= w4401 and w11524;
w15569 <= w7778 and not w15568;
w15570 <= not w15567 and w15569;
w15571 <= w7778 and not w15570;
w15572 <= not w15568 and not w15570;
w15573 <= not w15567 and w15572;
w15574 <= not w15571 and not w15573;
w15575 <= not w15564 and not w15574;
w15576 <= not w15564 and not w15575;
w15577 <= not w15574 and not w15575;
w15578 <= not w15576 and not w15577;
w15579 <= not w15424 and not w15427;
w15580 <= w15578 and w15579;
w15581 <= not w15578 and not w15579;
w15582 <= not w15580 and not w15581;
w15583 <= not w15407 and not w15409;
w15584 <= w2949 and w8793;
w15585 <= w2404 and w9895;
w15586 <= w3618 and w9315;
w15587 <= not w15585 and not w15586;
w15588 <= not w15584 and not w15587;
w15589 <= not w15584 and not w15588;
w15590 <= a(33) and a(58);
w15591 <= not w8114 and not w15590;
w15592 <= w15589 and not w15591;
w15593 <= a(60) and not w15588;
w15594 <= a(31) and w15593;
w15595 <= not w15592 and not w15594;
w15596 <= w4889 and w7239;
w15597 <= w5236 and w10711;
w15598 <= w4371 and w7505;
w15599 <= not w15597 and not w15598;
w15600 <= not w15596 and not w15599;
w15601 <= a(37) and not w15600;
w15602 <= a(54) and w15601;
w15603 <= not w15596 and not w15600;
w15604 <= a(38) and a(53);
w15605 <= a(39) and a(52);
w15606 <= not w15604 and not w15605;
w15607 <= w15603 and not w15606;
w15608 <= not w15602 and not w15607;
w15609 <= not w15493 and not w15608;
w15610 <= not w15493 and not w15609;
w15611 <= not w15608 and not w15609;
w15612 <= not w15610 and not w15611;
w15613 <= not w15595 and not w15612;
w15614 <= not w15595 and not w15613;
w15615 <= not w15612 and not w15613;
w15616 <= not w15614 and not w15615;
w15617 <= not w15583 and not w15616;
w15618 <= not w15583 and not w15617;
w15619 <= not w15616 and not w15617;
w15620 <= not w15618 and not w15619;
w15621 <= w15582 and not w15620;
w15622 <= not w15582 and w15620;
w15623 <= w15453 and w15512;
w15624 <= not w15453 and not w15512;
w15625 <= not w15623 and not w15624;
w15626 <= not w15521 and not w15525;
w15627 <= not w15625 and w15626;
w15628 <= w15625 and not w15626;
w15629 <= not w15627 and not w15628;
w15630 <= not w15499 and not w15505;
w15631 <= not w15629 and w15630;
w15632 <= w15629 and not w15630;
w15633 <= not w15631 and not w15632;
w15634 <= a(40) and a(51);
w15635 <= a(41) and a(50);
w15636 <= not w15634 and not w15635;
w15637 <= w5219 and w6370;
w15638 <= a(63) and not w15637;
w15639 <= a(28) and w15638;
w15640 <= not w15636 and w15639;
w15641 <= not w15637 and not w15640;
w15642 <= not w15636 and w15641;
w15643 <= a(63) and not w15640;
w15644 <= a(28) and w15643;
w15645 <= not w15642 and not w15644;
w15646 <= a(43) and a(48);
w15647 <= a(44) and a(47);
w15648 <= not w15646 and not w15647;
w15649 <= w5102 and w6058;
w15650 <= a(56) and not w15649;
w15651 <= a(35) and w15650;
w15652 <= not w15648 and w15651;
w15653 <= a(56) and not w15652;
w15654 <= a(35) and w15653;
w15655 <= not w15649 and not w15652;
w15656 <= not w15648 and w15655;
w15657 <= not w15654 and not w15656;
w15658 <= not w15645 and not w15657;
w15659 <= not w15645 and not w15658;
w15660 <= not w15657 and not w15658;
w15661 <= not w15659 and not w15660;
w15662 <= a(46) and a(62);
w15663 <= a(29) and w15662;
w15664 <= w5366 and not w15663;
w15665 <= w5366 and not w15664;
w15666 <= not w15663 and not w15664;
w15667 <= a(29) and a(62);
w15668 <= not a(46) and not w15667;
w15669 <= w15666 and not w15668;
w15670 <= not w15665 and not w15669;
w15671 <= not w15661 and not w15670;
w15672 <= not w15661 and not w15671;
w15673 <= not w15670 and not w15671;
w15674 <= not w15672 and not w15673;
w15675 <= not w15633 and w15674;
w15676 <= w15633 and not w15674;
w15677 <= not w15675 and not w15676;
w15678 <= not w15412 and not w15416;
w15679 <= w15677 and not w15678;
w15680 <= not w15677 and w15678;
w15681 <= not w15679 and not w15680;
w15682 <= not w15622 and w15681;
w15683 <= not w15621 and w15682;
w15684 <= w15681 and not w15683;
w15685 <= not w15622 and not w15683;
w15686 <= not w15621 and w15685;
w15687 <= not w15684 and not w15686;
w15688 <= not w15480 and not w15548;
w15689 <= not w15540 and not w15544;
w15690 <= not w15431 and not w15477;
w15691 <= a(30) and a(61);
w15692 <= not w15469 and w15691;
w15693 <= w15469 and not w15691;
w15694 <= not w15692 and not w15693;
w15695 <= w15441 and not w15694;
w15696 <= not w15441 and w15694;
w15697 <= not w15695 and not w15696;
w15698 <= not w15532 and not w15536;
w15699 <= not w15458 and not w15473;
w15700 <= w15698 and w15699;
w15701 <= not w15698 and not w15699;
w15702 <= not w15700 and not w15701;
w15703 <= w15697 and w15702;
w15704 <= not w15697 and not w15702;
w15705 <= not w15703 and not w15704;
w15706 <= not w15690 and w15705;
w15707 <= not w15690 and not w15706;
w15708 <= w15705 and not w15706;
w15709 <= not w15707 and not w15708;
w15710 <= not w15689 and not w15709;
w15711 <= not w15689 and not w15710;
w15712 <= not w15709 and not w15710;
w15713 <= not w15711 and not w15712;
w15714 <= not w15688 and not w15713;
w15715 <= not w15688 and not w15714;
w15716 <= not w15713 and not w15714;
w15717 <= not w15715 and not w15716;
w15718 <= not w15687 and w15717;
w15719 <= w15687 and not w15717;
w15720 <= not w15718 and not w15719;
w15721 <= not w15563 and not w15720;
w15722 <= w15563 and w15720;
w15723 <= not w15721 and not w15722;
w15724 <= not w15562 and not w15723;
w15725 <= w15562 and w15723;
w15726 <= not w15724 and not w15725;
w15727 <= not w15562 and not w15722;
w15728 <= not w15721 and not w15727;
w15729 <= not w15706 and not w15710;
w15730 <= not w15617 and not w15621;
w15731 <= not w15701 and not w15703;
w15732 <= w2671 and w9527;
w15733 <= a(61) and not w15732;
w15734 <= a(31) and w15733;
w15735 <= a(62) and not w15732;
w15736 <= a(30) and w15735;
w15737 <= not w15734 and not w15736;
w15738 <= not w15666 and not w15737;
w15739 <= not w15666 and not w15738;
w15740 <= not w15737 and not w15738;
w15741 <= not w15739 and not w15740;
w15742 <= w5219 and w6774;
w15743 <= w3790 and w7038;
w15744 <= w3977 and w7239;
w15745 <= not w15743 and not w15744;
w15746 <= not w15742 and not w15745;
w15747 <= a(53) and not w15746;
w15748 <= a(39) and w15747;
w15749 <= a(40) and a(52);
w15750 <= a(41) and a(51);
w15751 <= not w15749 and not w15750;
w15752 <= not w15742 and not w15746;
w15753 <= not w15751 and w15752;
w15754 <= not w15748 and not w15753;
w15755 <= not w15741 and not w15754;
w15756 <= not w15741 and not w15755;
w15757 <= not w15754 and not w15755;
w15758 <= not w15756 and not w15757;
w15759 <= not w15692 and not w15696;
w15760 <= w15758 and w15759;
w15761 <= not w15758 and not w15759;
w15762 <= not w15760 and not w15761;
w15763 <= a(42) and a(50);
w15764 <= a(34) and w15763;
w15765 <= a(58) and w15764;
w15766 <= w3125 and w8242;
w15767 <= not w15765 and not w15766;
w15768 <= a(35) and a(57);
w15769 <= w15763 and w15768;
w15770 <= not w15767 and not w15769;
w15771 <= not w15769 and not w15770;
w15772 <= not w15763 and not w15768;
w15773 <= w15771 and not w15772;
w15774 <= a(58) and not w15770;
w15775 <= a(34) and w15774;
w15776 <= not w15773 and not w15775;
w15777 <= w5519 and w6058;
w15778 <= w4617 and w6060;
w15779 <= w5102 and w6062;
w15780 <= not w15778 and not w15779;
w15781 <= not w15777 and not w15780;
w15782 <= a(49) and not w15781;
w15783 <= a(43) and w15782;
w15784 <= not w15777 and not w15781;
w15785 <= a(44) and a(48);
w15786 <= not w5056 and not w15785;
w15787 <= w15784 and not w15786;
w15788 <= not w15783 and not w15787;
w15789 <= not w15776 and not w15788;
w15790 <= not w15776 and not w15789;
w15791 <= not w15788 and not w15789;
w15792 <= not w15790 and not w15791;
w15793 <= a(36) and a(56);
w15794 <= a(33) and a(59);
w15795 <= not w13462 and not w15794;
w15796 <= w13462 and w15794;
w15797 <= w15793 and not w15796;
w15798 <= not w15795 and w15797;
w15799 <= w15793 and not w15798;
w15800 <= not w15796 and not w15798;
w15801 <= not w15795 and w15800;
w15802 <= not w15799 and not w15801;
w15803 <= not w15792 and not w15802;
w15804 <= not w15792 and not w15803;
w15805 <= not w15802 and not w15803;
w15806 <= not w15804 and not w15805;
w15807 <= not w15762 and w15806;
w15808 <= w15762 and not w15806;
w15809 <= not w15807 and not w15808;
w15810 <= not w15731 and w15809;
w15811 <= w15731 and not w15809;
w15812 <= not w15810 and not w15811;
w15813 <= not w15730 and w15812;
w15814 <= w15730 and not w15812;
w15815 <= not w15813 and not w15814;
w15816 <= not w15729 and w15815;
w15817 <= w15729 and not w15815;
w15818 <= not w15816 and not w15817;
w15819 <= not w15679 and not w15683;
w15820 <= not w15609 and not w15613;
w15821 <= not w15624 and not w15628;
w15822 <= w15820 and w15821;
w15823 <= not w15820 and not w15821;
w15824 <= not w15822 and not w15823;
w15825 <= not w15658 and not w15671;
w15826 <= not w15824 and w15825;
w15827 <= w15824 and not w15825;
w15828 <= not w15826 and not w15827;
w15829 <= not w15632 and not w15676;
w15830 <= not w15575 and not w15581;
w15831 <= w15589 and w15603;
w15832 <= not w15589 and not w15603;
w15833 <= not w15831 and not w15832;
w15834 <= w15641 and not w15833;
w15835 <= not w15641 and w15833;
w15836 <= not w15834 and not w15835;
w15837 <= w15572 and w15655;
w15838 <= not w15572 and not w15655;
w15839 <= not w15837 and not w15838;
w15840 <= w4371 and w7507;
w15841 <= a(37) and a(55);
w15842 <= a(38) and a(54);
w15843 <= not w15841 and not w15842;
w15844 <= not w15840 and not w15843;
w15845 <= a(60) and w15844;
w15846 <= a(32) and w15845;
w15847 <= a(60) and not w15846;
w15848 <= a(32) and w15847;
w15849 <= not w15840 and not w15846;
w15850 <= not w15843 and w15849;
w15851 <= not w15848 and not w15850;
w15852 <= w15839 and not w15851;
w15853 <= w15839 and not w15852;
w15854 <= not w15851 and not w15852;
w15855 <= not w15853 and not w15854;
w15856 <= not w15836 and w15855;
w15857 <= w15836 and not w15855;
w15858 <= not w15856 and not w15857;
w15859 <= not w15830 and w15858;
w15860 <= w15830 and not w15858;
w15861 <= not w15859 and not w15860;
w15862 <= not w15829 and w15861;
w15863 <= w15829 and not w15861;
w15864 <= not w15862 and not w15863;
w15865 <= w15828 and w15864;
w15866 <= not w15828 and not w15864;
w15867 <= not w15865 and not w15866;
w15868 <= not w15819 and w15867;
w15869 <= w15819 and not w15867;
w15870 <= not w15868 and not w15869;
w15871 <= w15818 and w15870;
w15872 <= not w15818 and not w15870;
w15873 <= not w15871 and not w15872;
w15874 <= not w15687 and not w15717;
w15875 <= not w15714 and not w15874;
w15876 <= not w15873 and w15875;
w15877 <= w15873 and not w15875;
w15878 <= not w15876 and not w15877;
w15879 <= w15728 and not w15878;
w15880 <= not w15728 and not w15876;
w15881 <= not w15877 and w15880;
w15882 <= not w15879 and not w15881;
w15883 <= not w15877 and not w15880;
w15884 <= not w15868 and not w15871;
w15885 <= not w15813 and not w15816;
w15886 <= not w15838 and not w15852;
w15887 <= not w15832 and not w15835;
w15888 <= w15886 and w15887;
w15889 <= not w15886 and not w15887;
w15890 <= not w15888 and not w15889;
w15891 <= not w15789 and not w15803;
w15892 <= not w15890 and w15891;
w15893 <= w15890 and not w15891;
w15894 <= not w15892 and not w15893;
w15895 <= not w15857 and not w15859;
w15896 <= w15894 and not w15895;
w15897 <= not w15894 and w15895;
w15898 <= not w15896 and not w15897;
w15899 <= not w15755 and not w15761;
w15900 <= w15771 and w15784;
w15901 <= not w15771 and not w15784;
w15902 <= not w15900 and not w15901;
w15903 <= w15752 and not w15902;
w15904 <= not w15752 and w15902;
w15905 <= not w15903 and not w15904;
w15906 <= w15800 and w15849;
w15907 <= not w15800 and not w15849;
w15908 <= not w15906 and not w15907;
w15909 <= not w15732 and not w15738;
w15910 <= not w15908 and w15909;
w15911 <= w15908 and not w15909;
w15912 <= not w15910 and not w15911;
w15913 <= w15905 and w15912;
w15914 <= not w15905 and not w15912;
w15915 <= not w15913 and not w15914;
w15916 <= not w15899 and w15915;
w15917 <= w15899 and not w15915;
w15918 <= not w15916 and not w15917;
w15919 <= w15898 and w15918;
w15920 <= not w15898 and not w15918;
w15921 <= not w15919 and not w15920;
w15922 <= w15885 and not w15921;
w15923 <= not w15885 and w15921;
w15924 <= not w15922 and not w15923;
w15925 <= not w15862 and not w15865;
w15926 <= not w15808 and not w15810;
w15927 <= not w15823 and not w15827;
w15928 <= w2949 and w9318;
w15929 <= w9281 and w11440;
w15930 <= w2294 and w9715;
w15931 <= not w15929 and not w15930;
w15932 <= not w15928 and not w15931;
w15933 <= not w15928 and not w15932;
w15934 <= a(32) and a(61);
w15935 <= a(33) and a(60);
w15936 <= not w15934 and not w15935;
w15937 <= w15933 and not w15936;
w15938 <= a(63) and not w15932;
w15939 <= a(30) and w15938;
w15940 <= not w15937 and not w15939;
w15941 <= w8742 and w13536;
w15942 <= w3634 and w8242;
w15943 <= a(39) and a(54);
w15944 <= w15009 and w15943;
w15945 <= not w15942 and not w15944;
w15946 <= not w15941 and not w15945;
w15947 <= w15009 and not w15946;
w15948 <= not w15941 and not w15946;
w15949 <= a(36) and a(57);
w15950 <= not w15943 and not w15949;
w15951 <= w15948 and not w15950;
w15952 <= not w15947 and not w15951;
w15953 <= not w15940 and not w15952;
w15954 <= not w15940 and not w15953;
w15955 <= not w15952 and not w15953;
w15956 <= not w15954 and not w15955;
w15957 <= a(40) and a(53);
w15958 <= a(41) and a(52);
w15959 <= not w15957 and not w15958;
w15960 <= w5219 and w7239;
w15961 <= w14994 and not w15960;
w15962 <= not w15959 and w15961;
w15963 <= w14994 and not w15962;
w15964 <= not w15960 and not w15962;
w15965 <= not w15959 and w15964;
w15966 <= not w15963 and not w15965;
w15967 <= not w15956 and not w15966;
w15968 <= not w15956 and not w15967;
w15969 <= not w15966 and not w15967;
w15970 <= not w15968 and not w15969;
w15971 <= a(38) and a(55);
w15972 <= not w7961 and not w15971;
w15973 <= a(45) and a(55);
w15974 <= w6748 and w15973;
w15975 <= w5952 and w9472;
w15976 <= w4371 and w8967;
w15977 <= not w15975 and not w15976;
w15978 <= not w15974 and not w15977;
w15979 <= not w15974 and not w15978;
w15980 <= not w15972 and w15979;
w15981 <= a(56) and not w15978;
w15982 <= a(37) and w15981;
w15983 <= not w15980 and not w15982;
w15984 <= w5102 and w6131;
w15985 <= w4445 and w9740;
w15986 <= w4824 and w6370;
w15987 <= not w15985 and not w15986;
w15988 <= not w15984 and not w15987;
w15989 <= a(51) and not w15988;
w15990 <= a(42) and w15989;
w15991 <= not w15984 and not w15988;
w15992 <= a(43) and a(50);
w15993 <= not w8058 and not w15992;
w15994 <= w15991 and not w15993;
w15995 <= not w15990 and not w15994;
w15996 <= not w15983 and not w15995;
w15997 <= not w15983 and not w15996;
w15998 <= not w15995 and not w15996;
w15999 <= not w15997 and not w15998;
w16000 <= a(47) and a(62);
w16001 <= a(31) and w16000;
w16002 <= w5472 and not w16001;
w16003 <= w5472 and not w16002;
w16004 <= not w16001 and not w16002;
w16005 <= a(31) and a(62);
w16006 <= not a(47) and not w16005;
w16007 <= w16004 and not w16006;
w16008 <= not w16003 and not w16007;
w16009 <= not w15999 and not w16008;
w16010 <= not w15999 and not w16009;
w16011 <= not w16008 and not w16009;
w16012 <= not w16010 and not w16011;
w16013 <= w15970 and w16012;
w16014 <= not w15970 and not w16012;
w16015 <= not w16013 and not w16014;
w16016 <= not w15927 and w16015;
w16017 <= w15927 and not w16015;
w16018 <= not w16016 and not w16017;
w16019 <= not w15926 and w16018;
w16020 <= w15926 and not w16018;
w16021 <= not w16019 and not w16020;
w16022 <= w15925 and not w16021;
w16023 <= not w15925 and w16021;
w16024 <= not w16022 and not w16023;
w16025 <= w15924 and w16024;
w16026 <= not w15924 and not w16024;
w16027 <= not w16025 and not w16026;
w16028 <= not w15884 and w16027;
w16029 <= w15884 and not w16027;
w16030 <= not w16028 and not w16029;
w16031 <= not w15883 and not w16030;
w16032 <= w15883 and w16030;
w16033 <= not w16031 and not w16032;
w16034 <= not w16019 and not w16023;
w16035 <= not w16014 and not w16016;
w16036 <= not w15907 and not w15911;
w16037 <= not w15901 and not w15904;
w16038 <= w16036 and w16037;
w16039 <= not w16036 and not w16037;
w16040 <= not w16038 and not w16039;
w16041 <= not w15953 and not w15967;
w16042 <= not w16040 and w16041;
w16043 <= w16040 and not w16041;
w16044 <= not w16042 and not w16043;
w16045 <= not w15913 and not w15916;
w16046 <= w16044 and not w16045;
w16047 <= not w16044 and w16045;
w16048 <= not w16046 and not w16047;
w16049 <= not w16035 and w16048;
w16050 <= w16035 and not w16048;
w16051 <= not w16049 and not w16050;
w16052 <= w16034 and not w16051;
w16053 <= not w16034 and w16051;
w16054 <= not w16052 and not w16053;
w16055 <= a(43) and a(51);
w16056 <= not w8060 and not w16055;
w16057 <= w5102 and w6370;
w16058 <= a(36) and not w16057;
w16059 <= a(58) and w16058;
w16060 <= not w16056 and w16059;
w16061 <= not w16057 and not w16060;
w16062 <= not w16056 and w16061;
w16063 <= a(58) and not w16060;
w16064 <= a(36) and w16063;
w16065 <= not w16062 and not w16064;
w16066 <= w5150 and w7239;
w16067 <= w6259 and w10711;
w16068 <= w5219 and w7505;
w16069 <= not w16067 and not w16068;
w16070 <= not w16066 and not w16069;
w16071 <= a(54) and not w16070;
w16072 <= a(40) and w16071;
w16073 <= a(42) and a(52);
w16074 <= not w8045 and not w16073;
w16075 <= not w16066 and not w16070;
w16076 <= not w16074 and w16075;
w16077 <= not w16072 and not w16076;
w16078 <= not w16065 and not w16077;
w16079 <= not w16065 and not w16078;
w16080 <= not w16077 and not w16078;
w16081 <= not w16079 and not w16080;
w16082 <= w8309 and w14375;
w16083 <= w5366 and w6062;
w16084 <= not w16082 and not w16083;
w16085 <= w8384 and w14375;
w16086 <= not w16084 and not w16085;
w16087 <= w8309 and not w16086;
w16088 <= not w16085 and not w16086;
w16089 <= not w8384 and not w14375;
w16090 <= w16088 and not w16089;
w16091 <= not w16087 and not w16090;
w16092 <= not w16081 and not w16091;
w16093 <= not w16081 and not w16092;
w16094 <= not w16091 and not w16092;
w16095 <= not w16093 and not w16094;
w16096 <= not w15889 and not w15893;
w16097 <= w16095 and w16096;
w16098 <= not w16095 and not w16096;
w16099 <= not w16097 and not w16098;
w16100 <= w2778 and w8711;
w16101 <= a(59) and a(62);
w16102 <= w6629 and w16101;
w16103 <= w2949 and w9527;
w16104 <= not w16102 and not w16103;
w16105 <= not w16100 and not w16104;
w16106 <= a(62) and not w16105;
w16107 <= a(32) and w16106;
w16108 <= not w16100 and not w16105;
w16109 <= a(33) and a(61);
w16110 <= a(35) and a(59);
w16111 <= not w16109 and not w16110;
w16112 <= w16108 and not w16111;
w16113 <= not w16107 and not w16112;
w16114 <= w15991 and not w16113;
w16115 <= not w15991 and w16113;
w16116 <= not w16114 and not w16115;
w16117 <= w5236 and w11524;
w16118 <= w11421 and w13018;
w16119 <= not w16117 and not w16118;
w16120 <= a(34) and a(60);
w16121 <= a(39) and a(55);
w16122 <= w16120 and w16121;
w16123 <= not w16119 and not w16122;
w16124 <= a(57) and not w16123;
w16125 <= a(37) and w16124;
w16126 <= not w16122 and not w16123;
w16127 <= not w16120 and not w16121;
w16128 <= w16126 and not w16127;
w16129 <= not w16125 and not w16128;
w16130 <= not w16116 and not w16129;
w16131 <= w16116 and w16129;
w16132 <= not w16130 and not w16131;
w16133 <= w16099 and w16132;
w16134 <= not w16099 and not w16132;
w16135 <= not w15896 and not w15919;
w16136 <= w12844 and not w16004;
w16137 <= not w12844 and w16004;
w16138 <= not w16136 and not w16137;
w16139 <= w15979 and not w16138;
w16140 <= not w15979 and w16138;
w16141 <= not w16139 and not w16140;
w16142 <= not w15996 and not w16009;
w16143 <= not w16141 and w16142;
w16144 <= w16141 and not w16142;
w16145 <= not w16143 and not w16144;
w16146 <= w15933 and w15948;
w16147 <= not w15933 and not w15948;
w16148 <= not w16146 and not w16147;
w16149 <= w15964 and not w16148;
w16150 <= not w15964 and w16148;
w16151 <= not w16149 and not w16150;
w16152 <= w16145 and w16151;
w16153 <= not w16145 and not w16151;
w16154 <= not w16152 and not w16153;
w16155 <= not w16135 and w16154;
w16156 <= w16135 and not w16154;
w16157 <= not w16155 and not w16156;
w16158 <= not w16134 and w16157;
w16159 <= not w16133 and w16158;
w16160 <= w16157 and not w16159;
w16161 <= not w16134 and not w16159;
w16162 <= not w16133 and w16161;
w16163 <= not w16160 and not w16162;
w16164 <= not w16054 and w16163;
w16165 <= w16054 and not w16163;
w16166 <= not w16164 and not w16165;
w16167 <= not w15923 and not w16025;
w16168 <= not w16166 and w16167;
w16169 <= w16166 and not w16167;
w16170 <= not w16168 and not w16169;
w16171 <= not w15883 and not w16029;
w16172 <= not w16028 and not w16171;
w16173 <= not w16170 and w16172;
w16174 <= w16170 and not w16172;
w16175 <= not w16173 and not w16174;
w16176 <= not w16155 and not w16159;
w16177 <= not w16098 and not w16133;
w16178 <= w3634 and w9315;
w16179 <= a(59) and not w16178;
w16180 <= a(36) and w16179;
w16181 <= a(60) and not w16178;
w16182 <= a(35) and w16181;
w16183 <= not w16180 and not w16182;
w16184 <= not w16088 and not w16183;
w16185 <= not w16088 and not w16184;
w16186 <= not w16183 and not w16184;
w16187 <= not w16185 and not w16186;
w16188 <= not w16136 and not w16140;
w16189 <= w16187 and w16188;
w16190 <= not w16187 and not w16188;
w16191 <= not w16189 and not w16190;
w16192 <= not w16147 and not w16150;
w16193 <= not w16191 and w16192;
w16194 <= w16191 and not w16192;
w16195 <= not w16193 and not w16194;
w16196 <= not w16144 and not w16152;
w16197 <= w16195 and not w16196;
w16198 <= not w16195 and w16196;
w16199 <= not w16197 and not w16198;
w16200 <= not w16177 and w16199;
w16201 <= w16177 and not w16199;
w16202 <= not w16200 and not w16201;
w16203 <= w16176 and not w16202;
w16204 <= not w16176 and w16202;
w16205 <= not w16203 and not w16204;
w16206 <= a(48) and a(62);
w16207 <= a(33) and w16206;
w16208 <= w6058 and not w16207;
w16209 <= not w16207 and not w16208;
w16210 <= a(33) and a(62);
w16211 <= not a(48) and not w16210;
w16212 <= w16209 and not w16211;
w16213 <= w6058 and not w16208;
w16214 <= not w16212 and not w16213;
w16215 <= w5366 and w6131;
w16216 <= a(46) and a(49);
w16217 <= not w8312 and not w16216;
w16218 <= not w16215 and not w16217;
w16219 <= a(56) and w16218;
w16220 <= a(39) and w16219;
w16221 <= a(56) and not w16220;
w16222 <= a(39) and w16221;
w16223 <= not w16215 and not w16220;
w16224 <= not w16217 and w16223;
w16225 <= not w16222 and not w16224;
w16226 <= not w16214 and not w16225;
w16227 <= not w16214 and not w16226;
w16228 <= not w16225 and not w16226;
w16229 <= not w16227 and not w16228;
w16230 <= w5102 and w6774;
w16231 <= w4445 and w7038;
w16232 <= w4824 and w7239;
w16233 <= not w16231 and not w16232;
w16234 <= not w16230 and not w16233;
w16235 <= a(53) and not w16234;
w16236 <= a(42) and w16235;
w16237 <= a(43) and a(52);
w16238 <= not w8292 and not w16237;
w16239 <= not w16230 and not w16234;
w16240 <= not w16238 and w16239;
w16241 <= not w16236 and not w16240;
w16242 <= not w16229 and not w16241;
w16243 <= not w16229 and not w16242;
w16244 <= not w16241 and not w16242;
w16245 <= not w16243 and not w16244;
w16246 <= not w16039 and not w16043;
w16247 <= w16245 and w16246;
w16248 <= not w16245 and not w16246;
w16249 <= not w16247 and not w16248;
w16250 <= a(32) and a(63);
w16251 <= a(34) and a(61);
w16252 <= not w16250 and not w16251;
w16253 <= w3896 and w9715;
w16254 <= a(54) and not w16253;
w16255 <= a(41) and w16254;
w16256 <= not w16252 and w16255;
w16257 <= not w16253 and not w16256;
w16258 <= not w16252 and w16257;
w16259 <= a(54) and not w16256;
w16260 <= a(41) and w16259;
w16261 <= not w16258 and not w16260;
w16262 <= w3609 and w11524;
w16263 <= a(55) and a(58);
w16264 <= w5501 and w16263;
w16265 <= w4371 and w8242;
w16266 <= not w16264 and not w16265;
w16267 <= not w16262 and not w16266;
w16268 <= a(37) and not w16267;
w16269 <= a(58) and w16268;
w16270 <= not w16262 and not w16267;
w16271 <= a(38) and a(57);
w16272 <= a(40) and a(55);
w16273 <= not w16271 and not w16272;
w16274 <= w16270 and not w16273;
w16275 <= not w16269 and not w16274;
w16276 <= not w16061 and not w16275;
w16277 <= not w16061 and not w16276;
w16278 <= not w16275 and not w16276;
w16279 <= not w16277 and not w16278;
w16280 <= not w16261 and not w16279;
w16281 <= not w16261 and not w16280;
w16282 <= not w16279 and not w16280;
w16283 <= not w16281 and not w16282;
w16284 <= w16249 and not w16283;
w16285 <= w16249 and not w16284;
w16286 <= not w16283 and not w16284;
w16287 <= not w16285 and not w16286;
w16288 <= not w16046 and not w16049;
w16289 <= w16108 and w16126;
w16290 <= not w16108 and not w16126;
w16291 <= not w16289 and not w16290;
w16292 <= w16075 and not w16291;
w16293 <= not w16075 and w16291;
w16294 <= not w16292 and not w16293;
w16295 <= not w16078 and not w16092;
w16296 <= not w15991 and not w16113;
w16297 <= not w16130 and not w16296;
w16298 <= w16295 and w16297;
w16299 <= not w16295 and not w16297;
w16300 <= not w16298 and not w16299;
w16301 <= w16294 and w16300;
w16302 <= not w16294 and not w16300;
w16303 <= not w16301 and not w16302;
w16304 <= not w16288 and w16303;
w16305 <= w16288 and not w16303;
w16306 <= not w16304 and not w16305;
w16307 <= w16287 and w16306;
w16308 <= not w16287 and not w16306;
w16309 <= not w16307 and not w16308;
w16310 <= w16205 and not w16309;
w16311 <= w16205 and not w16310;
w16312 <= not w16309 and not w16310;
w16313 <= not w16311 and not w16312;
w16314 <= not w16053 and not w16165;
w16315 <= not w16313 and not w16314;
w16316 <= w16313 and w16314;
w16317 <= not w16315 and not w16316;
w16318 <= not w16168 and not w16172;
w16319 <= not w16169 and not w16318;
w16320 <= not w16317 and w16319;
w16321 <= w16317 and not w16319;
w16322 <= not w16320 and not w16321;
w16323 <= not w16316 and not w16319;
w16324 <= not w16315 and not w16323;
w16325 <= not w16204 and not w16310;
w16326 <= not w16248 and not w16284;
w16327 <= w5501 and w13676;
w16328 <= w3493 and w9315;
w16329 <= a(40) and a(60);
w16330 <= w15793 and w16329;
w16331 <= not w16328 and not w16330;
w16332 <= not w16327 and not w16331;
w16333 <= not w16327 and not w16332;
w16334 <= a(37) and a(59);
w16335 <= a(40) and a(56);
w16336 <= not w16334 and not w16335;
w16337 <= w16333 and not w16336;
w16338 <= a(60) and not w16332;
w16339 <= a(36) and w16338;
w16340 <= not w16337 and not w16339;
w16341 <= a(38) and a(58);
w16342 <= a(39) and a(57);
w16343 <= not w16341 and not w16342;
w16344 <= w4889 and w8242;
w16345 <= w8506 and not w16344;
w16346 <= not w16343 and w16345;
w16347 <= w8506 and not w16346;
w16348 <= not w16344 and not w16346;
w16349 <= not w16343 and w16348;
w16350 <= not w16347 and not w16349;
w16351 <= not w16340 and not w16350;
w16352 <= not w16340 and not w16351;
w16353 <= not w16350 and not w16351;
w16354 <= not w16352 and not w16353;
w16355 <= a(45) and a(51);
w16356 <= w5472 and w6131;
w16357 <= w6060 and w16355;
w16358 <= w5366 and w6370;
w16359 <= not w16357 and not w16358;
w16360 <= not w16356 and not w16359;
w16361 <= w16355 and not w16360;
w16362 <= not w16356 and not w16360;
w16363 <= a(46) and a(50);
w16364 <= not w6060 and not w16363;
w16365 <= w16362 and not w16364;
w16366 <= not w16361 and not w16365;
w16367 <= not w16354 and not w16366;
w16368 <= not w16354 and not w16367;
w16369 <= not w16366 and not w16367;
w16370 <= not w16368 and not w16369;
w16371 <= not w16299 and not w16301;
w16372 <= not w16370 and not w16371;
w16373 <= not w16370 and not w16372;
w16374 <= not w16371 and not w16372;
w16375 <= not w16373 and not w16374;
w16376 <= not w16326 and not w16375;
w16377 <= not w16326 and not w16376;
w16378 <= not w16375 and not w16376;
w16379 <= not w16377 and not w16378;
w16380 <= not w16287 and w16306;
w16381 <= not w16304 and not w16380;
w16382 <= not w16379 and not w16381;
w16383 <= not w16379 and not w16382;
w16384 <= not w16381 and not w16382;
w16385 <= not w16383 and not w16384;
w16386 <= not w16197 and not w16200;
w16387 <= w16209 and w16223;
w16388 <= not w16209 and not w16223;
w16389 <= not w16387 and not w16388;
w16390 <= w16239 and not w16389;
w16391 <= not w16239 and w16389;
w16392 <= not w16390 and not w16391;
w16393 <= not w16276 and not w16280;
w16394 <= not w16226 and not w16242;
w16395 <= w16393 and w16394;
w16396 <= not w16393 and not w16394;
w16397 <= not w16395 and not w16396;
w16398 <= w16392 and w16397;
w16399 <= not w16392 and not w16397;
w16400 <= not w16398 and not w16399;
w16401 <= not w16386 and w16400;
w16402 <= w16386 and not w16400;
w16403 <= not w16401 and not w16402;
w16404 <= w3125 and w9527;
w16405 <= w2778 and w9715;
w16406 <= w3956 and w9598;
w16407 <= not w16405 and not w16406;
w16408 <= not w16404 and not w16407;
w16409 <= not w16404 and not w16408;
w16410 <= a(34) and a(62);
w16411 <= a(35) and a(61);
w16412 <= not w16410 and not w16411;
w16413 <= w16409 and not w16412;
w16414 <= a(63) and not w16408;
w16415 <= a(33) and w16414;
w16416 <= not w16413 and not w16415;
w16417 <= w4824 and w7505;
w16418 <= a(43) and a(53);
w16419 <= w8400 and w16418;
w16420 <= w5150 and w7507;
w16421 <= not w16419 and not w16420;
w16422 <= not w16417 and not w16421;
w16423 <= w8400 and not w16422;
w16424 <= a(42) and a(54);
w16425 <= not w16418 and not w16424;
w16426 <= not w16417 and not w16422;
w16427 <= not w16425 and w16426;
w16428 <= not w16423 and not w16427;
w16429 <= not w16416 and not w16428;
w16430 <= not w16416 and not w16429;
w16431 <= not w16428 and not w16429;
w16432 <= not w16430 and not w16431;
w16433 <= not w16290 and not w16293;
w16434 <= w16432 and w16433;
w16435 <= not w16432 and not w16433;
w16436 <= not w16434 and not w16435;
w16437 <= w16257 and w16270;
w16438 <= not w16257 and not w16270;
w16439 <= not w16437 and not w16438;
w16440 <= not w16178 and not w16184;
w16441 <= not w16439 and w16440;
w16442 <= w16439 and not w16440;
w16443 <= not w16441 and not w16442;
w16444 <= not w16190 and not w16194;
w16445 <= not w16443 and w16444;
w16446 <= w16443 and not w16444;
w16447 <= not w16445 and not w16446;
w16448 <= w16436 and w16447;
w16449 <= not w16436 and not w16447;
w16450 <= not w16448 and not w16449;
w16451 <= w16403 and w16450;
w16452 <= not w16403 and not w16450;
w16453 <= not w16451 and not w16452;
w16454 <= not w16385 and w16453;
w16455 <= not w16384 and not w16453;
w16456 <= not w16383 and w16455;
w16457 <= not w16454 and not w16456;
w16458 <= w16325 and not w16457;
w16459 <= not w16325 and w16457;
w16460 <= not w16458 and not w16459;
w16461 <= w16324 and not w16460;
w16462 <= not w16324 and not w16458;
w16463 <= not w16459 and w16462;
w16464 <= not w16461 and not w16463;
w16465 <= not w16459 and not w16462;
w16466 <= not w16382 and not w16454;
w16467 <= not w16372 and not w16376;
w16468 <= a(36) and a(61);
w16469 <= not w16362 and w16468;
w16470 <= w16362 and not w16468;
w16471 <= not w16469 and not w16470;
w16472 <= w16348 and not w16471;
w16473 <= not w16348 and w16471;
w16474 <= not w16472 and not w16473;
w16475 <= not w16351 and not w16367;
w16476 <= not w16438 and not w16442;
w16477 <= w16475 and w16476;
w16478 <= not w16475 and not w16476;
w16479 <= not w16477 and not w16478;
w16480 <= w16474 and w16479;
w16481 <= not w16474 and not w16479;
w16482 <= not w16480 and not w16481;
w16483 <= a(49) and a(62);
w16484 <= a(35) and w16483;
w16485 <= w6062 and not w16484;
w16486 <= not w16484 and not w16485;
w16487 <= a(35) and a(62);
w16488 <= not a(49) and not w16487;
w16489 <= w16486 and not w16488;
w16490 <= w6062 and not w16485;
w16491 <= not w16489 and not w16490;
w16492 <= a(47) and a(50);
w16493 <= not w8660 and not w16492;
w16494 <= w5472 and w6370;
w16495 <= a(57) and not w16494;
w16496 <= a(40) and w16495;
w16497 <= not w16493 and w16496;
w16498 <= a(57) and not w16497;
w16499 <= a(40) and w16498;
w16500 <= not w16494 and not w16497;
w16501 <= not w16493 and w16500;
w16502 <= not w16499 and not w16501;
w16503 <= not w16491 and not w16502;
w16504 <= not w16491 and not w16503;
w16505 <= not w16502 and not w16503;
w16506 <= not w16504 and not w16505;
w16507 <= not w16388 and not w16391;
w16508 <= w16506 and w16507;
w16509 <= not w16506 and not w16507;
w16510 <= not w16508 and not w16509;
w16511 <= w16333 and w16409;
w16512 <= not w16333 and not w16409;
w16513 <= not w16511 and not w16512;
w16514 <= w16426 and not w16513;
w16515 <= not w16426 and w16513;
w16516 <= not w16514 and not w16515;
w16517 <= not w16429 and not w16435;
w16518 <= not w16516 and w16517;
w16519 <= w16516 and not w16517;
w16520 <= not w16518 and not w16519;
w16521 <= w16510 and w16520;
w16522 <= not w16510 and not w16520;
w16523 <= not w16521 and not w16522;
w16524 <= w16482 and w16523;
w16525 <= not w16482 and not w16523;
w16526 <= not w16524 and not w16525;
w16527 <= w16467 and not w16526;
w16528 <= not w16467 and w16526;
w16529 <= not w16527 and not w16528;
w16530 <= not w16446 and not w16448;
w16531 <= w5150 and w8967;
w16532 <= a(34) and a(63);
w16533 <= a(41) and a(56);
w16534 <= w16532 and w16533;
w16535 <= not w16531 and not w16534;
w16536 <= a(42) and a(55);
w16537 <= w16532 and w16536;
w16538 <= not w16535 and not w16537;
w16539 <= not w16537 and not w16538;
w16540 <= not w16532 and not w16536;
w16541 <= w16539 and not w16540;
w16542 <= w16533 and not w16538;
w16543 <= not w16541 and not w16542;
w16544 <= w4889 and w8793;
w16545 <= w5236 and w9895;
w16546 <= w4371 and w9315;
w16547 <= not w16545 and not w16546;
w16548 <= not w16544 and not w16547;
w16549 <= a(60) and not w16548;
w16550 <= a(37) and w16549;
w16551 <= not w16544 and not w16548;
w16552 <= a(38) and a(59);
w16553 <= a(39) and a(58);
w16554 <= not w16552 and not w16553;
w16555 <= w16551 and not w16554;
w16556 <= not w16550 and not w16555;
w16557 <= not w16543 and not w16556;
w16558 <= not w16543 and not w16557;
w16559 <= not w16556 and not w16557;
w16560 <= not w16558 and not w16559;
w16561 <= w5519 and w7239;
w16562 <= w4617 and w10711;
w16563 <= w5102 and w7505;
w16564 <= not w16562 and not w16563;
w16565 <= not w16561 and not w16564;
w16566 <= a(54) and not w16565;
w16567 <= a(43) and w16566;
w16568 <= a(44) and a(53);
w16569 <= not w8914 and not w16568;
w16570 <= not w16561 and not w16565;
w16571 <= not w16569 and w16570;
w16572 <= not w16567 and not w16571;
w16573 <= not w16560 and not w16572;
w16574 <= not w16560 and not w16573;
w16575 <= not w16572 and not w16573;
w16576 <= not w16574 and not w16575;
w16577 <= not w16396 and not w16398;
w16578 <= not w16576 and not w16577;
w16579 <= not w16576 and not w16578;
w16580 <= not w16577 and not w16578;
w16581 <= not w16579 and not w16580;
w16582 <= not w16530 and not w16581;
w16583 <= not w16530 and not w16582;
w16584 <= not w16581 and not w16582;
w16585 <= not w16583 and not w16584;
w16586 <= not w16401 and not w16451;
w16587 <= w16585 and w16586;
w16588 <= not w16585 and not w16586;
w16589 <= not w16587 and not w16588;
w16590 <= w16529 and w16589;
w16591 <= not w16529 and not w16589;
w16592 <= not w16590 and not w16591;
w16593 <= not w16466 and w16592;
w16594 <= w16466 and not w16592;
w16595 <= not w16593 and not w16594;
w16596 <= not w16465 and not w16595;
w16597 <= w16465 and w16595;
w16598 <= not w16596 and not w16597;
w16599 <= not w16588 and not w16590;
w16600 <= not w16578 and not w16582;
w16601 <= not w16512 and not w16515;
w16602 <= not w16469 and not w16473;
w16603 <= w16601 and w16602;
w16604 <= not w16601 and not w16602;
w16605 <= not w16603 and not w16604;
w16606 <= not w16557 and not w16573;
w16607 <= not w16605 and w16606;
w16608 <= w16605 and not w16606;
w16609 <= not w16607 and not w16608;
w16610 <= w16539 and w16551;
w16611 <= not w16539 and not w16551;
w16612 <= not w16610 and not w16611;
w16613 <= w16570 and not w16612;
w16614 <= not w16570 and w16612;
w16615 <= not w16613 and not w16614;
w16616 <= not w16503 and not w16509;
w16617 <= not w16615 and w16616;
w16618 <= w16615 and not w16616;
w16619 <= not w16617 and not w16618;
w16620 <= a(39) and a(59);
w16621 <= a(40) and a(58);
w16622 <= not w16620 and not w16621;
w16623 <= w3977 and w8793;
w16624 <= a(45) and not w16623;
w16625 <= a(53) and w16624;
w16626 <= not w16622 and w16625;
w16627 <= not w16623 and not w16626;
w16628 <= not w16622 and w16627;
w16629 <= a(53) and not w16626;
w16630 <= a(45) and w16629;
w16631 <= not w16628 and not w16630;
w16632 <= w6058 and w6370;
w16633 <= w5472 and w6774;
w16634 <= a(48) and a(52);
w16635 <= w16363 and w16634;
w16636 <= not w16633 and not w16635;
w16637 <= not w16632 and not w16636;
w16638 <= a(52) and not w16637;
w16639 <= a(46) and w16638;
w16640 <= not w16632 and not w16637;
w16641 <= not w5694 and not w8933;
w16642 <= w16640 and not w16641;
w16643 <= not w16639 and not w16642;
w16644 <= not w16631 and not w16643;
w16645 <= not w16631 and not w16644;
w16646 <= not w16643 and not w16644;
w16647 <= not w16645 and not w16646;
w16648 <= w3493 and w9527;
w16649 <= a(37) and a(61);
w16650 <= not w11394 and not w16649;
w16651 <= not w16648 and not w16650;
w16652 <= not w16486 and w16651;
w16653 <= w16486 and not w16651;
w16654 <= not w16652 and not w16653;
w16655 <= w16647 and w16654;
w16656 <= not w16647 and not w16654;
w16657 <= not w16655 and not w16656;
w16658 <= w16619 and not w16657;
w16659 <= w16619 and not w16658;
w16660 <= not w16657 and not w16658;
w16661 <= not w16659 and not w16660;
w16662 <= w16609 and not w16661;
w16663 <= not w16609 and w16661;
w16664 <= not w16600 and not w16663;
w16665 <= not w16662 and w16664;
w16666 <= not w16600 and not w16665;
w16667 <= not w16662 and not w16665;
w16668 <= not w16663 and w16667;
w16669 <= not w16666 and not w16668;
w16670 <= not w16524 and not w16528;
w16671 <= not w16519 and not w16521;
w16672 <= w5102 and w7507;
w16673 <= a(43) and a(55);
w16674 <= a(44) and a(54);
w16675 <= not w16673 and not w16674;
w16676 <= not w16672 and not w16675;
w16677 <= a(35) and a(63);
w16678 <= not w16676 and not w16677;
w16679 <= w16676 and w16677;
w16680 <= not w16678 and not w16679;
w16681 <= not w16500 and w16680;
w16682 <= w16500 and not w16680;
w16683 <= not w16681 and not w16682;
w16684 <= a(38) and a(60);
w16685 <= a(41) and a(57);
w16686 <= a(42) and a(56);
w16687 <= not w16685 and not w16686;
w16688 <= w5150 and w8006;
w16689 <= w16684 and not w16688;
w16690 <= not w16687 and w16689;
w16691 <= w16684 and not w16690;
w16692 <= not w16688 and not w16690;
w16693 <= not w16687 and w16692;
w16694 <= not w16691 and not w16693;
w16695 <= w16683 and not w16694;
w16696 <= w16683 and not w16695;
w16697 <= not w16694 and not w16695;
w16698 <= not w16696 and not w16697;
w16699 <= not w16478 and not w16480;
w16700 <= not w16698 and not w16699;
w16701 <= not w16698 and not w16700;
w16702 <= not w16699 and not w16700;
w16703 <= not w16701 and not w16702;
w16704 <= not w16671 and not w16703;
w16705 <= w16671 and not w16702;
w16706 <= not w16701 and w16705;
w16707 <= not w16704 and not w16706;
w16708 <= not w16670 and w16707;
w16709 <= not w16670 and not w16708;
w16710 <= w16707 and not w16708;
w16711 <= not w16709 and not w16710;
w16712 <= not w16669 and not w16711;
w16713 <= w16669 and not w16710;
w16714 <= not w16709 and w16713;
w16715 <= not w16712 and not w16714;
w16716 <= w16599 and not w16715;
w16717 <= not w16599 and w16715;
w16718 <= not w16716 and not w16717;
w16719 <= not w16465 and not w16594;
w16720 <= not w16593 and not w16719;
w16721 <= not w16718 and w16720;
w16722 <= w16718 and not w16720;
w16723 <= not w16721 and not w16722;
w16724 <= not w16708 and not w16712;
w16725 <= not w16700 and not w16704;
w16726 <= not w16611 and not w16614;
w16727 <= a(50) and a(62);
w16728 <= a(37) and w16727;
w16729 <= w6131 and not w16728;
w16730 <= w6131 and not w16729;
w16731 <= not w16728 and not w16729;
w16732 <= a(37) and a(62);
w16733 <= not a(50) and not w16732;
w16734 <= w16731 and not w16733;
w16735 <= not w16730 and not w16734;
w16736 <= not w16726 and not w16735;
w16737 <= not w16726 and not w16736;
w16738 <= not w16735 and not w16736;
w16739 <= not w16737 and not w16738;
w16740 <= not w16681 and not w16695;
w16741 <= w16739 and w16740;
w16742 <= not w16739 and not w16740;
w16743 <= not w16741 and not w16742;
w16744 <= not w16648 and not w16652;
w16745 <= w16692 and w16744;
w16746 <= not w16692 and not w16744;
w16747 <= not w16745 and not w16746;
w16748 <= w4889 and w9318;
w16749 <= w8742 and w11440;
w16750 <= w3336 and w9715;
w16751 <= not w16749 and not w16750;
w16752 <= not w16748 and not w16751;
w16753 <= a(63) and not w16752;
w16754 <= a(36) and w16753;
w16755 <= not w16748 and not w16752;
w16756 <= a(38) and a(61);
w16757 <= a(39) and a(60);
w16758 <= not w16756 and not w16757;
w16759 <= w16755 and not w16758;
w16760 <= not w16754 and not w16759;
w16761 <= w16747 and not w16760;
w16762 <= w16747 and not w16761;
w16763 <= not w16760 and not w16761;
w16764 <= not w16762 and not w16763;
w16765 <= w16627 and w16640;
w16766 <= not w16627 and not w16640;
w16767 <= not w16765 and not w16766;
w16768 <= not w16672 and not w16679;
w16769 <= not w16767 and w16768;
w16770 <= w16767 and not w16768;
w16771 <= not w16769 and not w16770;
w16772 <= not w16647 and w16654;
w16773 <= not w16644 and not w16772;
w16774 <= w16771 and not w16773;
w16775 <= not w16771 and w16773;
w16776 <= not w16774 and not w16775;
w16777 <= not w16764 and not w16776;
w16778 <= w16764 and w16776;
w16779 <= not w16777 and not w16778;
w16780 <= w16743 and not w16779;
w16781 <= not w16743 and w16779;
w16782 <= not w16780 and not w16781;
w16783 <= not w16725 and w16782;
w16784 <= w16725 and not w16782;
w16785 <= not w16783 and not w16784;
w16786 <= a(41) and a(58);
w16787 <= not w9296 and not w16786;
w16788 <= w5219 and w8793;
w16789 <= a(44) and a(59);
w16790 <= w16272 and w16789;
w16791 <= not w16788 and not w16790;
w16792 <= w9296 and w16786;
w16793 <= not w16791 and not w16792;
w16794 <= not w16792 and not w16793;
w16795 <= not w16787 and w16794;
w16796 <= a(59) and not w16793;
w16797 <= a(40) and w16796;
w16798 <= not w16795 and not w16797;
w16799 <= w5472 and w7239;
w16800 <= w5056 and w10711;
w16801 <= w5366 and w7505;
w16802 <= not w16800 and not w16801;
w16803 <= not w16799 and not w16802;
w16804 <= a(54) and not w16803;
w16805 <= a(45) and w16804;
w16806 <= not w16799 and not w16803;
w16807 <= a(46) and a(53);
w16808 <= not w9234 and not w16807;
w16809 <= w16806 and not w16808;
w16810 <= not w16805 and not w16809;
w16811 <= not w16798 and not w16810;
w16812 <= not w16798 and not w16811;
w16813 <= not w16810 and not w16811;
w16814 <= not w16812 and not w16813;
w16815 <= a(48) and a(51);
w16816 <= a(42) and a(57);
w16817 <= a(43) and a(56);
w16818 <= not w16816 and not w16817;
w16819 <= w4824 and w8006;
w16820 <= w16815 and not w16819;
w16821 <= not w16818 and w16820;
w16822 <= w16815 and not w16821;
w16823 <= not w16819 and not w16821;
w16824 <= not w16818 and w16823;
w16825 <= not w16822 and not w16824;
w16826 <= not w16814 and not w16825;
w16827 <= not w16814 and not w16826;
w16828 <= not w16825 and not w16826;
w16829 <= not w16827 and not w16828;
w16830 <= not w16604 and not w16608;
w16831 <= w16829 and w16830;
w16832 <= not w16829 and not w16830;
w16833 <= not w16831 and not w16832;
w16834 <= not w16618 and not w16658;
w16835 <= not w16833 and w16834;
w16836 <= w16833 and not w16834;
w16837 <= not w16835 and not w16836;
w16838 <= not w16667 and w16837;
w16839 <= w16837 and not w16838;
w16840 <= not w16667 and not w16838;
w16841 <= not w16839 and not w16840;
w16842 <= w16785 and not w16841;
w16843 <= not w16785 and not w16840;
w16844 <= not w16839 and w16843;
w16845 <= not w16842 and not w16844;
w16846 <= not w16724 and w16845;
w16847 <= w16724 and not w16845;
w16848 <= not w16846 and not w16847;
w16849 <= not w16716 and not w16720;
w16850 <= not w16717 and not w16849;
w16851 <= not w16848 and w16850;
w16852 <= w16848 and not w16850;
w16853 <= not w16851 and not w16852;
w16854 <= not w16847 and not w16850;
w16855 <= not w16846 and not w16854;
w16856 <= not w16838 and not w16842;
w16857 <= not w16766 and not w16770;
w16858 <= w6062 and w6774;
w16859 <= w6060 and w7038;
w16860 <= w6058 and w7239;
w16861 <= not w16859 and not w16860;
w16862 <= not w16858 and not w16861;
w16863 <= a(53) and not w16862;
w16864 <= a(47) and w16863;
w16865 <= not w16858 and not w16862;
w16866 <= not w9740 and not w16634;
w16867 <= w16865 and not w16866;
w16868 <= not w16864 and not w16867;
w16869 <= not w16857 and not w16868;
w16870 <= not w16857 and not w16869;
w16871 <= not w16868 and not w16869;
w16872 <= not w16870 and not w16871;
w16873 <= not w16746 and not w16761;
w16874 <= w16872 and w16873;
w16875 <= not w16872 and not w16873;
w16876 <= not w16874 and not w16875;
w16877 <= not w16832 and not w16836;
w16878 <= not w16876 and w16877;
w16879 <= w16876 and not w16877;
w16880 <= not w16878 and not w16879;
w16881 <= w16755 and w16806;
w16882 <= not w16755 and not w16806;
w16883 <= not w16881 and not w16882;
w16884 <= w16794 and not w16883;
w16885 <= not w16794 and w16883;
w16886 <= not w16884 and not w16885;
w16887 <= not w16811 and not w16826;
w16888 <= not w16886 and w16887;
w16889 <= w16886 and not w16887;
w16890 <= not w16888 and not w16889;
w16891 <= a(37) and a(63);
w16892 <= not w16731 and w16891;
w16893 <= w16731 and not w16891;
w16894 <= not w16892 and not w16893;
w16895 <= w16823 and not w16894;
w16896 <= not w16823 and w16894;
w16897 <= not w16895 and not w16896;
w16898 <= w16890 and w16897;
w16899 <= not w16890 and not w16897;
w16900 <= not w16898 and not w16899;
w16901 <= w16880 and w16900;
w16902 <= not w16880 and not w16900;
w16903 <= not w16901 and not w16902;
w16904 <= not w16780 and not w16783;
w16905 <= w3977 and w9318;
w16906 <= w13350 and w16684;
w16907 <= w4889 and w9527;
w16908 <= not w16906 and not w16907;
w16909 <= not w16905 and not w16908;
w16910 <= not w16905 and not w16909;
w16911 <= a(39) and a(61);
w16912 <= not w16329 and not w16911;
w16913 <= w16910 and not w16912;
w16914 <= w12377 and not w16909;
w16915 <= not w16913 and not w16914;
w16916 <= w5519 and w8967;
w16917 <= w4617 and w11524;
w16918 <= w5102 and w8006;
w16919 <= not w16917 and not w16918;
w16920 <= not w16916 and not w16919;
w16921 <= w10109 and not w16920;
w16922 <= not w9299 and not w15973;
w16923 <= not w16916 and not w16920;
w16924 <= not w16922 and w16923;
w16925 <= not w16921 and not w16924;
w16926 <= not w16915 and not w16925;
w16927 <= not w16915 and not w16926;
w16928 <= not w16925 and not w16926;
w16929 <= not w16927 and not w16928;
w16930 <= a(41) and a(59);
w16931 <= a(42) and a(58);
w16932 <= not w16930 and not w16931;
w16933 <= w5150 and w8793;
w16934 <= w9220 and not w16933;
w16935 <= not w16932 and w16934;
w16936 <= w9220 and not w16935;
w16937 <= not w16933 and not w16935;
w16938 <= not w16932 and w16937;
w16939 <= not w16936 and not w16938;
w16940 <= not w16929 and not w16939;
w16941 <= not w16929 and not w16940;
w16942 <= not w16939 and not w16940;
w16943 <= not w16941 and not w16942;
w16944 <= not w16736 and not w16742;
w16945 <= w16943 and w16944;
w16946 <= not w16943 and not w16944;
w16947 <= not w16945 and not w16946;
w16948 <= not w16764 and w16776;
w16949 <= not w16774 and not w16948;
w16950 <= w16947 and not w16949;
w16951 <= not w16947 and w16949;
w16952 <= not w16950 and not w16951;
w16953 <= not w16904 and w16952;
w16954 <= w16904 and not w16952;
w16955 <= not w16953 and not w16954;
w16956 <= w16903 and w16955;
w16957 <= not w16903 and not w16955;
w16958 <= not w16956 and not w16957;
w16959 <= not w16856 and w16958;
w16960 <= w16856 and not w16958;
w16961 <= not w16959 and not w16960;
w16962 <= w16855 and not w16961;
w16963 <= not w16855 and not w16960;
w16964 <= not w16959 and w16963;
w16965 <= not w16962 and not w16964;
w16966 <= not w16959 and not w16963;
w16967 <= not w16953 and not w16956;
w16968 <= not w16879 and not w16901;
w16969 <= a(46) and a(55);
w16970 <= a(47) and a(54);
w16971 <= not w16969 and not w16970;
w16972 <= w5472 and w7507;
w16973 <= a(38) and not w16972;
w16974 <= a(63) and w16973;
w16975 <= not w16971 and w16974;
w16976 <= not w16972 and not w16975;
w16977 <= not w16971 and w16976;
w16978 <= a(63) and not w16975;
w16979 <= a(38) and w16978;
w16980 <= not w16977 and not w16979;
w16981 <= w4617 and w7748;
w16982 <= w13676 and w14973;
w16983 <= w4824 and w8793;
w16984 <= not w16982 and not w16983;
w16985 <= not w16981 and not w16984;
w16986 <= a(59) and not w16985;
w16987 <= a(42) and w16986;
w16988 <= not w16981 and not w16985;
w16989 <= a(43) and a(58);
w16990 <= a(45) and a(56);
w16991 <= not w16989 and not w16990;
w16992 <= w16988 and not w16991;
w16993 <= not w16987 and not w16992;
w16994 <= not w16980 and not w16993;
w16995 <= not w16980 and not w16994;
w16996 <= not w16993 and not w16994;
w16997 <= not w16995 and not w16996;
w16998 <= w8506 and w12407;
w16999 <= w6062 and w7239;
w17000 <= a(44) and a(57);
w17001 <= w10245 and w17000;
w17002 <= not w16999 and not w17001;
w17003 <= not w16998 and not w17002;
w17004 <= w10245 and not w17003;
w17005 <= not w16998 and not w17003;
w17006 <= a(49) and a(52);
w17007 <= not w17000 and not w17006;
w17008 <= w17005 and not w17007;
w17009 <= not w17004 and not w17008;
w17010 <= not w16997 and not w17009;
w17011 <= not w16997 and not w17010;
w17012 <= not w17009 and not w17010;
w17013 <= not w17011 and not w17012;
w17014 <= not w16869 and not w16875;
w17015 <= w17013 and w17014;
w17016 <= not w17013 and not w17014;
w17017 <= not w17015 and not w17016;
w17018 <= not w16892 and not w16896;
w17019 <= w5219 and w9318;
w17020 <= a(60) and not w17019;
w17021 <= a(41) and w17020;
w17022 <= a(61) and not w17019;
w17023 <= a(40) and w17022;
w17024 <= not w17021 and not w17023;
w17025 <= not w16865 and not w17024;
w17026 <= not w16865 and not w17025;
w17027 <= not w17024 and not w17025;
w17028 <= not w17026 and not w17027;
w17029 <= a(62) and w7580;
w17030 <= w6370 and not w17029;
w17031 <= not w17029 and not w17030;
w17032 <= a(39) and a(62);
w17033 <= not a(51) and not w17032;
w17034 <= w17031 and not w17033;
w17035 <= w6370 and not w17030;
w17036 <= not w17034 and not w17035;
w17037 <= not w17028 and not w17036;
w17038 <= not w17028 and not w17037;
w17039 <= not w17036 and not w17037;
w17040 <= not w17038 and not w17039;
w17041 <= not w17018 and not w17040;
w17042 <= not w17018 and not w17041;
w17043 <= not w17040 and not w17041;
w17044 <= not w17042 and not w17043;
w17045 <= w17017 and not w17044;
w17046 <= not w17017 and w17044;
w17047 <= not w16968 and not w17046;
w17048 <= not w17045 and w17047;
w17049 <= not w16968 and not w17048;
w17050 <= not w17046 and not w17048;
w17051 <= not w17045 and w17050;
w17052 <= not w17049 and not w17051;
w17053 <= not w16946 and not w16950;
w17054 <= not w16889 and not w16898;
w17055 <= not w17053 and not w17054;
w17056 <= not w17053 and not w17055;
w17057 <= not w17054 and not w17055;
w17058 <= not w17056 and not w17057;
w17059 <= w16910 and w16937;
w17060 <= not w16910 and not w16937;
w17061 <= not w17059 and not w17060;
w17062 <= w16923 and not w17061;
w17063 <= not w16923 and w17061;
w17064 <= not w17062 and not w17063;
w17065 <= not w16926 and not w16940;
w17066 <= not w16882 and not w16885;
w17067 <= w17065 and w17066;
w17068 <= not w17065 and not w17066;
w17069 <= not w17067 and not w17068;
w17070 <= w17064 and w17069;
w17071 <= not w17064 and not w17069;
w17072 <= not w17070 and not w17071;
w17073 <= not w17058 and w17072;
w17074 <= not w17058 and not w17073;
w17075 <= w17072 and not w17073;
w17076 <= not w17074 and not w17075;
w17077 <= not w17052 and w17076;
w17078 <= w17052 and not w17076;
w17079 <= not w17077 and not w17078;
w17080 <= not w16967 and not w17079;
w17081 <= w16967 and w17079;
w17082 <= not w17080 and not w17081;
w17083 <= not w16966 and not w17082;
w17084 <= w16966 and w17082;
w17085 <= not w17083 and not w17084;
w17086 <= not w16966 and not w17081;
w17087 <= not w17080 and not w17086;
w17088 <= not w17052 and not w17076;
w17089 <= not w17048 and not w17088;
w17090 <= not w17055 and not w17073;
w17091 <= not w17019 and not w17025;
w17092 <= w16988 and w17091;
w17093 <= not w16988 and not w17091;
w17094 <= not w17092 and not w17093;
w17095 <= w5150 and w9318;
w17096 <= w11440 and w13777;
w17097 <= w3790 and w9715;
w17098 <= not w17096 and not w17097;
w17099 <= not w17095 and not w17098;
w17100 <= a(63) and not w17099;
w17101 <= a(39) and w17100;
w17102 <= not w17095 and not w17099;
w17103 <= a(41) and a(61);
w17104 <= a(42) and a(60);
w17105 <= not w17103 and not w17104;
w17106 <= w17102 and not w17105;
w17107 <= not w17101 and not w17106;
w17108 <= w17094 and not w17107;
w17109 <= w17094 and not w17108;
w17110 <= not w17107 and not w17108;
w17111 <= not w17109 and not w17110;
w17112 <= not w17037 and not w17041;
w17113 <= w17111 and w17112;
w17114 <= not w17111 and not w17112;
w17115 <= not w17113 and not w17114;
w17116 <= a(43) and a(59);
w17117 <= a(44) and a(58);
w17118 <= not w17116 and not w17117;
w17119 <= w5102 and w8793;
w17120 <= w13350 and not w17119;
w17121 <= not w17118 and w17120;
w17122 <= not w17119 and not w17121;
w17123 <= not w17118 and w17122;
w17124 <= w13350 and not w17121;
w17125 <= not w17123 and not w17124;
w17126 <= w5472 and w8967;
w17127 <= w5056 and w11524;
w17128 <= w5366 and w8006;
w17129 <= not w17127 and not w17128;
w17130 <= not w17126 and not w17129;
w17131 <= a(57) and not w17130;
w17132 <= a(45) and w17131;
w17133 <= a(46) and a(56);
w17134 <= a(47) and a(55);
w17135 <= not w17133 and not w17134;
w17136 <= not w17126 and not w17130;
w17137 <= not w17135 and w17136;
w17138 <= not w17132 and not w17137;
w17139 <= not w17125 and not w17138;
w17140 <= not w17125 and not w17139;
w17141 <= not w17138 and not w17139;
w17142 <= not w17140 and not w17141;
w17143 <= w6131 and w7239;
w17144 <= w5694 and w10711;
w17145 <= w6062 and w7505;
w17146 <= not w17144 and not w17145;
w17147 <= not w17143 and not w17146;
w17148 <= a(54) and not w17147;
w17149 <= a(48) and w17148;
w17150 <= not w17143 and not w17147;
w17151 <= a(49) and a(53);
w17152 <= not w6772 and not w17151;
w17153 <= w17150 and not w17152;
w17154 <= not w17149 and not w17153;
w17155 <= not w17142 and not w17154;
w17156 <= not w17142 and not w17155;
w17157 <= not w17154 and not w17155;
w17158 <= not w17156 and not w17157;
w17159 <= w17115 and not w17158;
w17160 <= not w17115 and w17158;
w17161 <= not w17090 and not w17160;
w17162 <= not w17159 and w17161;
w17163 <= not w17090 and not w17162;
w17164 <= not w17160 and not w17162;
w17165 <= not w17159 and w17164;
w17166 <= not w17163 and not w17165;
w17167 <= w17005 and w17031;
w17168 <= not w17005 and not w17031;
w17169 <= not w17167 and not w17168;
w17170 <= w16976 and not w17169;
w17171 <= not w16976 and w17169;
w17172 <= not w17170 and not w17171;
w17173 <= not w17060 and not w17063;
w17174 <= not w17172 and w17173;
w17175 <= w17172 and not w17173;
w17176 <= not w17174 and not w17175;
w17177 <= not w16994 and not w17010;
w17178 <= not w17176 and w17177;
w17179 <= w17176 and not w17177;
w17180 <= not w17178 and not w17179;
w17181 <= not w17016 and not w17045;
w17182 <= not w17068 and not w17070;
w17183 <= not w17181 and not w17182;
w17184 <= not w17181 and not w17183;
w17185 <= not w17182 and not w17183;
w17186 <= not w17184 and not w17185;
w17187 <= w17180 and not w17186;
w17188 <= not w17180 and w17186;
w17189 <= not w17166 and not w17188;
w17190 <= not w17187 and w17189;
w17191 <= not w17166 and not w17190;
w17192 <= not w17188 and not w17190;
w17193 <= not w17187 and w17192;
w17194 <= not w17191 and not w17193;
w17195 <= w17089 and w17194;
w17196 <= not w17089 and not w17194;
w17197 <= not w17195 and not w17196;
w17198 <= w17087 and not w17197;
w17199 <= not w17087 and not w17195;
w17200 <= not w17196 and w17199;
w17201 <= not w17198 and not w17200;
w17202 <= not w17196 and not w17199;
w17203 <= not w17183 and not w17187;
w17204 <= a(46) and a(57);
w17205 <= a(47) and a(56);
w17206 <= not w17204 and not w17205;
w17207 <= w5472 and w8006;
w17208 <= a(43) and not w17207;
w17209 <= a(60) and w17208;
w17210 <= not w17206 and w17209;
w17211 <= not w17207 and not w17210;
w17212 <= not w17206 and w17211;
w17213 <= a(60) and not w17210;
w17214 <= a(43) and w17213;
w17215 <= not w17212 and not w17214;
w17216 <= w6131 and w7505;
w17217 <= w5694 and w7503;
w17218 <= w6062 and w7507;
w17219 <= not w17217 and not w17218;
w17220 <= not w17216 and not w17219;
w17221 <= a(55) and not w17220;
w17222 <= a(48) and w17221;
w17223 <= not w17216 and not w17220;
w17224 <= a(50) and a(53);
w17225 <= not w11919 and not w17224;
w17226 <= w17223 and not w17225;
w17227 <= not w17222 and not w17226;
w17228 <= not w17215 and not w17227;
w17229 <= not w17215 and not w17228;
w17230 <= not w17227 and not w17228;
w17231 <= not w17229 and not w17230;
w17232 <= a(52) and w13666;
w17233 <= w6774 and not w17232;
w17234 <= w6774 and not w17233;
w17235 <= not w17232 and not w17233;
w17236 <= not a(52) and not w13666;
w17237 <= w17235 and not w17236;
w17238 <= not w17234 and not w17237;
w17239 <= not w17231 and not w17238;
w17240 <= not w17231 and not w17239;
w17241 <= not w17238 and not w17239;
w17242 <= not w17240 and not w17241;
w17243 <= a(40) and a(63);
w17244 <= not w17150 and w17243;
w17245 <= w17150 and not w17243;
w17246 <= not w17244 and not w17245;
w17247 <= w17136 and not w17246;
w17248 <= not w17136 and w17246;
w17249 <= not w17247 and not w17248;
w17250 <= w17102 and w17122;
w17251 <= not w17102 and not w17122;
w17252 <= not w17250 and not w17251;
w17253 <= w5519 and w8793;
w17254 <= w4445 and w8711;
w17255 <= a(45) and a(61);
w17256 <= w16931 and w17255;
w17257 <= not w17254 and not w17256;
w17258 <= not w17253 and not w17257;
w17259 <= a(61) and not w17258;
w17260 <= a(42) and w17259;
w17261 <= a(45) and a(58);
w17262 <= not w16789 and not w17261;
w17263 <= not w17253 and not w17258;
w17264 <= not w17262 and w17263;
w17265 <= not w17260 and not w17264;
w17266 <= w17252 and not w17265;
w17267 <= w17252 and not w17266;
w17268 <= not w17265 and not w17266;
w17269 <= not w17267 and not w17268;
w17270 <= not w17249 and w17269;
w17271 <= w17249 and not w17269;
w17272 <= not w17270 and not w17271;
w17273 <= not w17242 and w17272;
w17274 <= not w17242 and not w17273;
w17275 <= w17272 and not w17273;
w17276 <= not w17274 and not w17275;
w17277 <= not w17203 and not w17276;
w17278 <= not w17203 and not w17277;
w17279 <= not w17276 and not w17277;
w17280 <= not w17278 and not w17279;
w17281 <= not w17093 and not w17108;
w17282 <= not w17168 and not w17171;
w17283 <= w17281 and w17282;
w17284 <= not w17281 and not w17282;
w17285 <= not w17283 and not w17284;
w17286 <= not w17139 and not w17155;
w17287 <= not w17285 and w17286;
w17288 <= w17285 and not w17286;
w17289 <= not w17287 and not w17288;
w17290 <= not w17114 and not w17159;
w17291 <= not w17175 and not w17179;
w17292 <= w17290 and w17291;
w17293 <= not w17290 and not w17291;
w17294 <= not w17292 and not w17293;
w17295 <= w17289 and w17294;
w17296 <= not w17289 and not w17294;
w17297 <= not w17295 and not w17296;
w17298 <= not w17280 and w17297;
w17299 <= not w17280 and not w17298;
w17300 <= w17297 and not w17298;
w17301 <= not w17299 and not w17300;
w17302 <= not w17162 and not w17190;
w17303 <= not w17301 and not w17302;
w17304 <= w17301 and w17302;
w17305 <= not w17303 and not w17304;
w17306 <= not w17202 and not w17305;
w17307 <= w17202 and w17305;
w17308 <= not w17306 and not w17307;
w17309 <= not w17202 and not w17304;
w17310 <= not w17303 and not w17309;
w17311 <= not w17277 and not w17298;
w17312 <= not w17293 and not w17295;
w17313 <= w17211 and w17223;
w17314 <= not w17211 and not w17223;
w17315 <= not w17313 and not w17314;
w17316 <= w17263 and not w17315;
w17317 <= not w17263 and w17315;
w17318 <= not w17316 and not w17317;
w17319 <= not w17228 and not w17239;
w17320 <= not w17318 and w17319;
w17321 <= w17318 and not w17319;
w17322 <= not w17320 and not w17321;
w17323 <= a(43) and a(61);
w17324 <= a(45) and a(59);
w17325 <= not w17323 and not w17324;
w17326 <= w4617 and w8711;
w17327 <= w5102 and w9318;
w17328 <= w5519 and w9315;
w17329 <= not w17327 and not w17328;
w17330 <= not w17326 and not w17329;
w17331 <= not w17326 and not w17330;
w17332 <= not w17325 and w17331;
w17333 <= a(60) and not w17330;
w17334 <= a(44) and w17333;
w17335 <= not w17332 and not w17334;
w17336 <= w6058 and w8006;
w17337 <= w5472 and w8242;
w17338 <= a(48) and a(58);
w17339 <= w17133 and w17338;
w17340 <= not w17337 and not w17339;
w17341 <= not w17336 and not w17340;
w17342 <= a(58) and not w17341;
w17343 <= a(46) and w17342;
w17344 <= not w17336 and not w17341;
w17345 <= a(47) and a(57);
w17346 <= not w9472 and not w17345;
w17347 <= w17344 and not w17346;
w17348 <= not w17343 and not w17347;
w17349 <= not w17335 and not w17348;
w17350 <= not w17335 and not w17349;
w17351 <= not w17348 and not w17349;
w17352 <= not w17350 and not w17351;
w17353 <= w6370 and w7505;
w17354 <= w7038 and w9607;
w17355 <= w6131 and w7507;
w17356 <= not w17354 and not w17355;
w17357 <= not w17353 and not w17356;
w17358 <= w9607 and not w17357;
w17359 <= not w17353 and not w17357;
w17360 <= a(50) and a(54);
w17361 <= not w7038 and not w17360;
w17362 <= w17359 and not w17361;
w17363 <= not w17358 and not w17362;
w17364 <= not w17352 and not w17363;
w17365 <= not w17352 and not w17364;
w17366 <= not w17363 and not w17364;
w17367 <= not w17365 and not w17366;
w17368 <= w17322 and not w17367;
w17369 <= not w17322 and w17367;
w17370 <= not w17312 and not w17369;
w17371 <= not w17368 and w17370;
w17372 <= not w17312 and not w17371;
w17373 <= not w17369 and not w17371;
w17374 <= not w17368 and w17373;
w17375 <= not w17372 and not w17374;
w17376 <= not w17271 and not w17273;
w17377 <= not w17284 and not w17288;
w17378 <= w17376 and w17377;
w17379 <= not w17376 and not w17377;
w17380 <= not w17378 and not w17379;
w17381 <= not w17244 and not w17248;
w17382 <= w5150 and w9598;
w17383 <= a(41) and a(63);
w17384 <= not w14174 and not w17383;
w17385 <= not w17382 and not w17384;
w17386 <= not w17235 and w17385;
w17387 <= w17235 and not w17385;
w17388 <= not w17386 and not w17387;
w17389 <= w17381 and not w17388;
w17390 <= not w17381 and w17388;
w17391 <= not w17389 and not w17390;
w17392 <= not w17251 and not w17266;
w17393 <= not w17391 and w17392;
w17394 <= w17391 and not w17392;
w17395 <= not w17393 and not w17394;
w17396 <= w17380 and w17395;
w17397 <= not w17380 and not w17395;
w17398 <= not w17396 and not w17397;
w17399 <= not w17375 and w17398;
w17400 <= not w17375 and not w17399;
w17401 <= w17398 and not w17399;
w17402 <= not w17400 and not w17401;
w17403 <= not w17311 and not w17402;
w17404 <= w17311 and w17402;
w17405 <= not w17403 and not w17404;
w17406 <= not w17310 and w17405;
w17407 <= w17310 and not w17405;
w17408 <= not w17406 and not w17407;
w17409 <= w17344 and w17359;
w17410 <= not w17344 and not w17359;
w17411 <= not w17409 and not w17410;
w17412 <= w17331 and not w17411;
w17413 <= not w17331 and w17411;
w17414 <= not w17412 and not w17413;
w17415 <= not w17349 and not w17364;
w17416 <= not w17414 and w17415;
w17417 <= w17414 and not w17415;
w17418 <= not w17416 and not w17417;
w17419 <= not w17390 and not w17394;
w17420 <= not w17418 and w17419;
w17421 <= w17418 and not w17419;
w17422 <= not w17420 and not w17421;
w17423 <= not w17379 and not w17396;
w17424 <= w17422 and not w17423;
w17425 <= not w17422 and w17423;
w17426 <= not w17424 and not w17425;
w17427 <= not w17321 and not w17368;
w17428 <= a(62) and w16418;
w17429 <= w7239 and not w17428;
w17430 <= not w17428 and not w17429;
w17431 <= not a(53) and not w14538;
w17432 <= w17430 and not w17431;
w17433 <= w7239 and not w17429;
w17434 <= not w17432 and not w17433;
w17435 <= w6370 and w7507;
w17436 <= w7227 and w9740;
w17437 <= w6131 and w8967;
w17438 <= not w17436 and not w17437;
w17439 <= not w17435 and not w17438;
w17440 <= a(56) and not w17439;
w17441 <= a(49) and w17440;
w17442 <= a(51) and a(54);
w17443 <= a(50) and a(55);
w17444 <= not w17442 and not w17443;
w17445 <= not w17435 and not w17439;
w17446 <= not w17444 and w17445;
w17447 <= not w17441 and not w17446;
w17448 <= not w17434 and not w17447;
w17449 <= not w17434 and not w17448;
w17450 <= not w17447 and not w17448;
w17451 <= not w17449 and not w17450;
w17452 <= not w17314 and not w17317;
w17453 <= w17451 and w17452;
w17454 <= not w17451 and not w17452;
w17455 <= not w17453 and not w17454;
w17456 <= w5519 and w9318;
w17457 <= w11440 and w14973;
w17458 <= w4445 and w9715;
w17459 <= not w17457 and not w17458;
w17460 <= not w17456 and not w17459;
w17461 <= a(42) and not w17460;
w17462 <= a(63) and w17461;
w17463 <= not w17456 and not w17460;
w17464 <= a(44) and a(61);
w17465 <= a(45) and a(60);
w17466 <= not w17464 and not w17465;
w17467 <= w17463 and not w17466;
w17468 <= not w17462 and not w17467;
w17469 <= not w17382 and not w17386;
w17470 <= not w17468 and w17469;
w17471 <= w17468 and not w17469;
w17472 <= not w17470 and not w17471;
w17473 <= w6058 and w8242;
w17474 <= w8384 and w8791;
w17475 <= w5472 and w8793;
w17476 <= not w17474 and not w17475;
w17477 <= not w17473 and not w17476;
w17478 <= a(59) and not w17477;
w17479 <= a(46) and w17478;
w17480 <= not w17473 and not w17477;
w17481 <= a(47) and a(58);
w17482 <= a(48) and a(57);
w17483 <= not w17481 and not w17482;
w17484 <= w17480 and not w17483;
w17485 <= not w17479 and not w17484;
w17486 <= not w17472 and not w17485;
w17487 <= w17472 and w17485;
w17488 <= not w17486 and not w17487;
w17489 <= not w17455 and not w17488;
w17490 <= w17455 and w17488;
w17491 <= not w17489 and not w17490;
w17492 <= not w17427 and w17491;
w17493 <= w17427 and not w17491;
w17494 <= not w17492 and not w17493;
w17495 <= w17426 and w17494;
w17496 <= not w17426 and not w17494;
w17497 <= not w17495 and not w17496;
w17498 <= not w17371 and not w17399;
w17499 <= not w17497 and w17498;
w17500 <= w17497 and not w17498;
w17501 <= not w17499 and not w17500;
w17502 <= not w17310 and not w17404;
w17503 <= not w17403 and not w17502;
w17504 <= not w17501 and w17503;
w17505 <= w17501 and not w17503;
w17506 <= not w17504 and not w17505;
w17507 <= not w17499 and not w17503;
w17508 <= not w17500 and not w17507;
w17509 <= not w17424 and not w17495;
w17510 <= not w17417 and not w17421;
w17511 <= w6062 and w8242;
w17512 <= w6060 and w8791;
w17513 <= w6058 and w8793;
w17514 <= not w17512 and not w17513;
w17515 <= not w17511 and not w17514;
w17516 <= not w17511 and not w17515;
w17517 <= not w12407 and not w17338;
w17518 <= w17516 and not w17517;
w17519 <= a(59) and not w17515;
w17520 <= a(47) and w17519;
w17521 <= not w17518 and not w17520;
w17522 <= w6774 and w7507;
w17523 <= w6772 and w7227;
w17524 <= w6370 and w8967;
w17525 <= not w17523 and not w17524;
w17526 <= not w17522 and not w17525;
w17527 <= a(56) and not w17526;
w17528 <= a(50) and w17527;
w17529 <= not w17522 and not w17526;
w17530 <= a(51) and a(55);
w17531 <= not w10711 and not w17530;
w17532 <= w17529 and not w17531;
w17533 <= not w17528 and not w17532;
w17534 <= not w17521 and not w17533;
w17535 <= not w17521 and not w17534;
w17536 <= not w17533 and not w17534;
w17537 <= not w17535 and not w17536;
w17538 <= not w17410 and not w17413;
w17539 <= w17537 and w17538;
w17540 <= not w17537 and not w17538;
w17541 <= not w17539 and not w17540;
w17542 <= w17463 and w17480;
w17543 <= not w17463 and not w17480;
w17544 <= not w17542 and not w17543;
w17545 <= w5366 and w9318;
w17546 <= w5519 and w9527;
w17547 <= a(46) and a(60);
w17548 <= w14913 and w17547;
w17549 <= not w17546 and not w17548;
w17550 <= not w17545 and not w17549;
w17551 <= w14913 and not w17550;
w17552 <= not w17545 and not w17550;
w17553 <= not w17255 and not w17547;
w17554 <= w17552 and not w17553;
w17555 <= not w17551 and not w17554;
w17556 <= w17544 and not w17555;
w17557 <= w17544 and not w17556;
w17558 <= not w17555 and not w17556;
w17559 <= not w17557 and not w17558;
w17560 <= w17541 and not w17559;
w17561 <= not w17541 and w17559;
w17562 <= not w17510 and not w17561;
w17563 <= not w17560 and w17562;
w17564 <= not w17510 and not w17563;
w17565 <= not w17560 and not w17563;
w17566 <= not w17561 and w17565;
w17567 <= not w17564 and not w17566;
w17568 <= a(43) and a(63);
w17569 <= not w17430 and w17568;
w17570 <= w17430 and not w17568;
w17571 <= not w17569 and not w17570;
w17572 <= w17445 and not w17571;
w17573 <= not w17445 and w17571;
w17574 <= not w17572 and not w17573;
w17575 <= not w17468 and not w17469;
w17576 <= not w17486 and not w17575;
w17577 <= not w17574 and w17576;
w17578 <= w17574 and not w17576;
w17579 <= not w17577 and not w17578;
w17580 <= not w17448 and not w17454;
w17581 <= not w17579 and w17580;
w17582 <= w17579 and not w17580;
w17583 <= not w17581 and not w17582;
w17584 <= not w17490 and not w17492;
w17585 <= w17583 and not w17584;
w17586 <= not w17583 and w17584;
w17587 <= not w17585 and not w17586;
w17588 <= w17567 and w17587;
w17589 <= not w17567 and not w17587;
w17590 <= not w17588 and not w17589;
w17591 <= not w17509 and not w17590;
w17592 <= w17509 and w17590;
w17593 <= not w17591 and not w17592;
w17594 <= w17508 and not w17593;
w17595 <= not w17508 and not w17592;
w17596 <= not w17591 and w17595;
w17597 <= not w17594 and not w17596;
w17598 <= not w17591 and not w17595;
w17599 <= not w17567 and w17587;
w17600 <= not w17585 and not w17599;
w17601 <= not w17578 and not w17582;
w17602 <= w17516 and w17552;
w17603 <= not w17516 and not w17552;
w17604 <= not w17602 and not w17603;
w17605 <= a(58) and a(63);
w17606 <= w8058 and w17605;
w17607 <= w6062 and w8793;
w17608 <= a(59) and a(63);
w17609 <= w15785 and w17608;
w17610 <= not w17607 and not w17609;
w17611 <= not w17606 and not w17610;
w17612 <= a(59) and not w17611;
w17613 <= a(48) and w17612;
w17614 <= a(44) and a(63);
w17615 <= a(49) and a(58);
w17616 <= not w17614 and not w17615;
w17617 <= not w17606 and not w17611;
w17618 <= not w17616 and w17617;
w17619 <= not w17613 and not w17618;
w17620 <= w17604 and not w17619;
w17621 <= w17604 and not w17620;
w17622 <= not w17619 and not w17620;
w17623 <= not w17621 and not w17622;
w17624 <= a(54) and w15269;
w17625 <= w7505 and not w17624;
w17626 <= not w17624 and not w17625;
w17627 <= not a(54) and not w15269;
w17628 <= w17626 and not w17627;
w17629 <= w7505 and not w17625;
w17630 <= not w17628 and not w17629;
w17631 <= w6774 and w8967;
w17632 <= w6772 and w11524;
w17633 <= w6370 and w8006;
w17634 <= not w17632 and not w17633;
w17635 <= not w17631 and not w17634;
w17636 <= a(57) and not w17635;
w17637 <= a(50) and w17636;
w17638 <= not w17631 and not w17635;
w17639 <= a(51) and a(56);
w17640 <= not w12194 and not w17639;
w17641 <= w17638 and not w17640;
w17642 <= not w17637 and not w17641;
w17643 <= not w17630 and not w17642;
w17644 <= not w17630 and not w17643;
w17645 <= not w17642 and not w17643;
w17646 <= not w17644 and not w17645;
w17647 <= w5472 and w9318;
w17648 <= a(60) and not w17647;
w17649 <= a(47) and w17648;
w17650 <= a(46) and not w17647;
w17651 <= a(61) and w17650;
w17652 <= not w17649 and not w17651;
w17653 <= not w17529 and not w17652;
w17654 <= not w17529 and not w17653;
w17655 <= not w17652 and not w17653;
w17656 <= not w17654 and not w17655;
w17657 <= not w17646 and w17656;
w17658 <= w17646 and not w17656;
w17659 <= not w17657 and not w17658;
w17660 <= not w17623 and not w17659;
w17661 <= w17623 and w17659;
w17662 <= not w17660 and not w17661;
w17663 <= w17601 and not w17662;
w17664 <= not w17601 and w17662;
w17665 <= not w17663 and not w17664;
w17666 <= not w17543 and not w17556;
w17667 <= not w17569 and not w17573;
w17668 <= w17666 and w17667;
w17669 <= not w17666 and not w17667;
w17670 <= not w17668 and not w17669;
w17671 <= not w17534 and not w17540;
w17672 <= not w17670 and w17671;
w17673 <= w17670 and not w17671;
w17674 <= not w17672 and not w17673;
w17675 <= not w17565 and w17674;
w17676 <= w17565 and not w17674;
w17677 <= not w17675 and not w17676;
w17678 <= w17665 and w17677;
w17679 <= not w17665 and not w17677;
w17680 <= not w17678 and not w17679;
w17681 <= w17600 and not w17680;
w17682 <= not w17600 and w17680;
w17683 <= not w17681 and not w17682;
w17684 <= not w17598 and not w17683;
w17685 <= w17598 and w17683;
w17686 <= not w17684 and not w17685;
w17687 <= not w17598 and not w17681;
w17688 <= not w17682 and not w17687;
w17689 <= not w17675 and not w17678;
w17690 <= not w17603 and not w17620;
w17691 <= w7239 and w8967;
w17692 <= w7038 and w11524;
w17693 <= w6774 and w8006;
w17694 <= not w17692 and not w17693;
w17695 <= not w17691 and not w17694;
w17696 <= w14223 and not w17695;
w17697 <= not w17691 and not w17695;
w17698 <= a(52) and a(56);
w17699 <= not w7503 and not w17698;
w17700 <= w17697 and not w17699;
w17701 <= not w17696 and not w17700;
w17702 <= not w17690 and not w17701;
w17703 <= not w17690 and not w17702;
w17704 <= not w17701 and not w17702;
w17705 <= not w17703 and not w17704;
w17706 <= not w17646 and not w17656;
w17707 <= not w17643 and not w17706;
w17708 <= not w17705 and not w17707;
w17709 <= not w17705 and not w17708;
w17710 <= not w17707 and not w17708;
w17711 <= not w17709 and not w17710;
w17712 <= not w17660 and not w17664;
w17713 <= w17711 and w17712;
w17714 <= not w17711 and not w17712;
w17715 <= not w17713 and not w17714;
w17716 <= w17626 and w17638;
w17717 <= not w17626 and not w17638;
w17718 <= not w17716 and not w17717;
w17719 <= w17617 and not w17718;
w17720 <= not w17617 and w17718;
w17721 <= not w17719 and not w17720;
w17722 <= not w17669 and not w17673;
w17723 <= not w17721 and w17722;
w17724 <= w17721 and not w17722;
w17725 <= not w17723 and not w17724;
w17726 <= w5472 and w9527;
w17727 <= w5056 and w9715;
w17728 <= w5366 and w9598;
w17729 <= not w17727 and not w17728;
w17730 <= not w17726 and not w17729;
w17731 <= a(45) and not w17730;
w17732 <= a(63) and w17731;
w17733 <= not w17726 and not w17730;
w17734 <= a(47) and a(61);
w17735 <= not w15662 and not w17734;
w17736 <= w17733 and not w17735;
w17737 <= not w17732 and not w17736;
w17738 <= not w17647 and not w17653;
w17739 <= not w17737 and w17738;
w17740 <= w17737 and not w17738;
w17741 <= not w17739 and not w17740;
w17742 <= w6131 and w8793;
w17743 <= w5694 and w9895;
w17744 <= w6062 and w9315;
w17745 <= not w17743 and not w17744;
w17746 <= not w17742 and not w17745;
w17747 <= a(60) and not w17746;
w17748 <= a(48) and w17747;
w17749 <= a(49) and a(59);
w17750 <= a(50) and a(58);
w17751 <= not w17749 and not w17750;
w17752 <= not w17742 and not w17746;
w17753 <= not w17751 and w17752;
w17754 <= not w17748 and not w17753;
w17755 <= not w17741 and not w17754;
w17756 <= w17741 and w17754;
w17757 <= not w17755 and not w17756;
w17758 <= w17725 and w17757;
w17759 <= not w17725 and not w17757;
w17760 <= w17715 and not w17759;
w17761 <= not w17758 and w17760;
w17762 <= w17715 and not w17761;
w17763 <= not w17759 and not w17761;
w17764 <= not w17758 and w17763;
w17765 <= not w17762 and not w17764;
w17766 <= w17689 and w17765;
w17767 <= not w17689 and not w17765;
w17768 <= not w17766 and not w17767;
w17769 <= w17688 and not w17768;
w17770 <= not w17688 and not w17766;
w17771 <= not w17767 and w17770;
w17772 <= not w17769 and not w17771;
w17773 <= not w17767 and not w17770;
w17774 <= not w17717 and not w17720;
w17775 <= a(55) and w16000;
w17776 <= w7507 and not w17775;
w17777 <= w7507 and not w17776;
w17778 <= not w17775 and not w17776;
w17779 <= not a(55) and not w16000;
w17780 <= w17778 and not w17779;
w17781 <= not w17777 and not w17780;
w17782 <= not w17774 and not w17781;
w17783 <= not w17774 and not w17782;
w17784 <= not w17781 and not w17782;
w17785 <= not w17783 and not w17784;
w17786 <= not w17737 and not w17738;
w17787 <= not w17755 and not w17786;
w17788 <= w17785 and w17787;
w17789 <= not w17785 and not w17787;
w17790 <= not w17788 and not w17789;
w17791 <= not w17724 and not w17758;
w17792 <= w17790 and not w17791;
w17793 <= not w17790 and w17791;
w17794 <= not w17792 and not w17793;
w17795 <= a(46) and a(63);
w17796 <= not w17697 and w17795;
w17797 <= w17697 and not w17795;
w17798 <= not w17796 and not w17797;
w17799 <= w17752 and not w17798;
w17800 <= not w17752 and w17798;
w17801 <= not w17799 and not w17800;
w17802 <= not w17702 and not w17708;
w17803 <= not w17801 and w17802;
w17804 <= w17801 and not w17802;
w17805 <= not w17803 and not w17804;
w17806 <= w6131 and w9315;
w17807 <= w5694 and w8711;
w17808 <= w6062 and w9318;
w17809 <= not w17807 and not w17808;
w17810 <= not w17806 and not w17809;
w17811 <= a(48) and not w17810;
w17812 <= a(61) and w17811;
w17813 <= not w17806 and not w17810;
w17814 <= a(49) and a(60);
w17815 <= a(50) and a(59);
w17816 <= not w17814 and not w17815;
w17817 <= w17813 and not w17816;
w17818 <= not w17812 and not w17817;
w17819 <= w17733 and not w17818;
w17820 <= not w17733 and w17818;
w17821 <= not w17819 and not w17820;
w17822 <= a(51) and a(58);
w17823 <= w7239 and w8006;
w17824 <= w7038 and w7748;
w17825 <= w6774 and w8242;
w17826 <= not w17824 and not w17825;
w17827 <= not w17823 and not w17826;
w17828 <= w17822 and not w17827;
w17829 <= not w17823 and not w17827;
w17830 <= a(52) and a(57);
w17831 <= not w13094 and not w17830;
w17832 <= w17829 and not w17831;
w17833 <= not w17828 and not w17832;
w17834 <= not w17821 and not w17833;
w17835 <= w17821 and w17833;
w17836 <= not w17834 and not w17835;
w17837 <= w17805 and w17836;
w17838 <= not w17805 and not w17836;
w17839 <= w17794 and not w17838;
w17840 <= not w17837 and w17839;
w17841 <= w17794 and not w17840;
w17842 <= not w17838 and not w17840;
w17843 <= not w17837 and w17842;
w17844 <= not w17841 and not w17843;
w17845 <= not w17714 and not w17761;
w17846 <= not w17844 and not w17845;
w17847 <= w17844 and w17845;
w17848 <= not w17846 and not w17847;
w17849 <= not w17773 and not w17848;
w17850 <= w17773 and w17848;
w17851 <= not w17849 and not w17850;
w17852 <= not w17773 and not w17847;
w17853 <= not w17846 and not w17852;
w17854 <= not w17792 and not w17840;
w17855 <= w17813 and w17829;
w17856 <= not w17813 and not w17829;
w17857 <= not w17855 and not w17856;
w17858 <= w6370 and w9315;
w17859 <= w8711 and w9740;
w17860 <= w6131 and w9318;
w17861 <= not w17859 and not w17860;
w17862 <= not w17858 and not w17861;
w17863 <= a(61) and not w17862;
w17864 <= a(49) and w17863;
w17865 <= not w17858 and not w17862;
w17866 <= a(50) and a(60);
w17867 <= a(51) and a(59);
w17868 <= not w17866 and not w17867;
w17869 <= w17865 and not w17868;
w17870 <= not w17864 and not w17869;
w17871 <= w17857 and not w17870;
w17872 <= w17857 and not w17871;
w17873 <= not w17870 and not w17871;
w17874 <= not w17872 and not w17873;
w17875 <= not w17733 and not w17818;
w17876 <= not w17834 and not w17875;
w17877 <= w17874 and w17876;
w17878 <= not w17874 and not w17876;
w17879 <= not w17877 and not w17878;
w17880 <= not w17782 and not w17789;
w17881 <= not w17879 and w17880;
w17882 <= w17879 and not w17880;
w17883 <= not w17881 and not w17882;
w17884 <= w7505 and w8006;
w17885 <= w7239 and w8242;
w17886 <= a(54) and a(58);
w17887 <= w17698 and w17886;
w17888 <= not w17885 and not w17887;
w17889 <= not w17884 and not w17888;
w17890 <= a(58) and not w17889;
w17891 <= a(52) and w17890;
w17892 <= not w17884 and not w17889;
w17893 <= a(53) and a(57);
w17894 <= not w7227 and not w17893;
w17895 <= w17892 and not w17894;
w17896 <= not w17891 and not w17895;
w17897 <= w6058 and w9598;
w17898 <= a(47) and a(63);
w17899 <= not w16206 and not w17898;
w17900 <= not w17897 and not w17899;
w17901 <= not w17778 and w17900;
w17902 <= w17778 and not w17900;
w17903 <= not w17901 and not w17902;
w17904 <= not w17896 and w17903;
w17905 <= w17903 and not w17904;
w17906 <= not w17896 and not w17904;
w17907 <= not w17905 and not w17906;
w17908 <= not w17796 and not w17800;
w17909 <= w17907 and w17908;
w17910 <= not w17907 and not w17908;
w17911 <= not w17909 and not w17910;
w17912 <= not w17804 and not w17837;
w17913 <= w17911 and not w17912;
w17914 <= w17911 and not w17913;
w17915 <= not w17912 and not w17913;
w17916 <= not w17914 and not w17915;
w17917 <= w17883 and not w17916;
w17918 <= not w17883 and not w17915;
w17919 <= not w17914 and w17918;
w17920 <= not w17917 and not w17919;
w17921 <= w17854 and not w17920;
w17922 <= not w17854 and w17920;
w17923 <= not w17921 and not w17922;
w17924 <= w17853 and not w17923;
w17925 <= not w17853 and not w17921;
w17926 <= not w17922 and w17925;
w17927 <= not w17924 and not w17926;
w17928 <= not w17922 and not w17925;
w17929 <= not w17913 and not w17917;
w17930 <= w17865 and w17892;
w17931 <= not w17865 and not w17892;
w17932 <= not w17930 and not w17931;
w17933 <= not w17897 and not w17901;
w17934 <= not w17932 and w17933;
w17935 <= w17932 and not w17933;
w17936 <= not w17934 and not w17935;
w17937 <= not w17856 and not w17871;
w17938 <= not w17936 and w17937;
w17939 <= w17936 and not w17937;
w17940 <= not w17938 and not w17939;
w17941 <= not w17904 and not w17910;
w17942 <= not w17940 and w17941;
w17943 <= w17940 and not w17941;
w17944 <= not w17942 and not w17943;
w17945 <= w6370 and w9318;
w17946 <= w11440 and w16815;
w17947 <= w5694 and w9715;
w17948 <= not w17946 and not w17947;
w17949 <= not w17945 and not w17948;
w17950 <= not w17945 and not w17949;
w17951 <= a(50) and a(61);
w17952 <= a(51) and a(60);
w17953 <= not w17951 and not w17952;
w17954 <= w17950 and not w17953;
w17955 <= a(63) and not w17949;
w17956 <= a(48) and w17955;
w17957 <= not w17954 and not w17956;
w17958 <= a(56) and a(62);
w17959 <= a(49) and w17958;
w17960 <= w8967 and not w17959;
w17961 <= w8967 and not w17960;
w17962 <= not w17959 and not w17960;
w17963 <= not a(56) and not w16483;
w17964 <= w17962 and not w17963;
w17965 <= not w17961 and not w17964;
w17966 <= not w17957 and not w17965;
w17967 <= not w17957 and not w17966;
w17968 <= not w17965 and not w17966;
w17969 <= not w17967 and not w17968;
w17970 <= w7505 and w8242;
w17971 <= w8791 and w10711;
w17972 <= w7239 and w8793;
w17973 <= not w17971 and not w17972;
w17974 <= not w17970 and not w17973;
w17975 <= a(59) and not w17974;
w17976 <= a(52) and w17975;
w17977 <= a(53) and a(58);
w17978 <= not w13536 and not w17977;
w17979 <= not w17970 and not w17974;
w17980 <= not w17978 and w17979;
w17981 <= not w17976 and not w17980;
w17982 <= not w17969 and not w17981;
w17983 <= not w17969 and not w17982;
w17984 <= not w17981 and not w17982;
w17985 <= not w17983 and not w17984;
w17986 <= not w17878 and not w17882;
w17987 <= w17985 and w17986;
w17988 <= not w17985 and not w17986;
w17989 <= not w17987 and not w17988;
w17990 <= w17944 and w17989;
w17991 <= not w17944 and not w17989;
w17992 <= not w17990 and not w17991;
w17993 <= not w17929 and w17992;
w17994 <= w17929 and not w17992;
w17995 <= not w17993 and not w17994;
w17996 <= not w17928 and not w17995;
w17997 <= w17928 and w17995;
w17998 <= not w17996 and not w17997;
w17999 <= not w17928 and not w17994;
w18000 <= not w17993 and not w17999;
w18001 <= not w17988 and not w17990;
w18002 <= not w17939 and not w17943;
w18003 <= a(52) and w11440;
w18004 <= a(51) and w9715;
w18005 <= not w18003 and not w18004;
w18006 <= w6774 and w9318;
w18007 <= a(49) and not w18006;
w18008 <= not w18005 and w18007;
w18009 <= a(49) and not w18008;
w18010 <= a(63) and w18009;
w18011 <= not w18006 and not w18008;
w18012 <= a(51) and a(61);
w18013 <= a(52) and a(60);
w18014 <= not w18012 and not w18013;
w18015 <= w18011 and not w18014;
w18016 <= not w18010 and not w18015;
w18017 <= w17950 and not w18016;
w18018 <= not w17950 and w18016;
w18019 <= not w18017 and not w18018;
w18020 <= w7507 and w8242;
w18021 <= w7505 and w8793;
w18022 <= a(55) and a(59);
w18023 <= w17893 and w18022;
w18024 <= not w18021 and not w18023;
w18025 <= not w18020 and not w18024;
w18026 <= a(59) and not w18025;
w18027 <= a(53) and w18026;
w18028 <= not w18020 and not w18025;
w18029 <= not w11524 and not w17886;
w18030 <= w18028 and not w18029;
w18031 <= not w18027 and not w18030;
w18032 <= not w18019 and not w18031;
w18033 <= w18019 and w18031;
w18034 <= not w18032 and not w18033;
w18035 <= w18002 and not w18034;
w18036 <= not w18002 and w18034;
w18037 <= not w18035 and not w18036;
w18038 <= w16727 and not w17962;
w18039 <= not w16727 and w17962;
w18040 <= not w18038 and not w18039;
w18041 <= w17979 and not w18040;
w18042 <= not w17979 and w18040;
w18043 <= not w18041 and not w18042;
w18044 <= not w17931 and not w17935;
w18045 <= not w17966 and not w17982;
w18046 <= w18044 and w18045;
w18047 <= not w18044 and not w18045;
w18048 <= not w18046 and not w18047;
w18049 <= w18043 and w18048;
w18050 <= not w18043 and not w18048;
w18051 <= not w18049 and not w18050;
w18052 <= w18037 and w18051;
w18053 <= not w18037 and not w18051;
w18054 <= not w18052 and not w18053;
w18055 <= w18001 and not w18054;
w18056 <= not w18001 and w18054;
w18057 <= not w18055 and not w18056;
w18058 <= w18000 and not w18057;
w18059 <= not w18000 and not w18055;
w18060 <= not w18056 and w18059;
w18061 <= not w18058 and not w18060;
w18062 <= not w18056 and not w18059;
w18063 <= not w18036 and not w18052;
w18064 <= w7239 and w9318;
w18065 <= a(60) and not w18064;
w18066 <= a(53) and w18065;
w18067 <= a(52) and not w18064;
w18068 <= a(61) and w18067;
w18069 <= not w18066 and not w18068;
w18070 <= not w18028 and not w18069;
w18071 <= not w18028 and not w18070;
w18072 <= not w18069 and not w18070;
w18073 <= not w18071 and not w18072;
w18074 <= not w18038 and not w18042;
w18075 <= w18073 and w18074;
w18076 <= not w18073 and not w18074;
w18077 <= not w18075 and not w18076;
w18078 <= not w17950 and not w18016;
w18079 <= not w18032 and not w18078;
w18080 <= not w18077 and w18079;
w18081 <= w18077 and not w18079;
w18082 <= not w18080 and not w18081;
w18083 <= not w18047 and not w18049;
w18084 <= a(54) and a(59);
w18085 <= not w16263 and not w18084;
w18086 <= w7507 and w8793;
w18087 <= a(50) and not w18086;
w18088 <= a(63) and w18087;
w18089 <= not w18085 and w18088;
w18090 <= a(50) and not w18089;
w18091 <= a(63) and w18090;
w18092 <= not w18086 and not w18089;
w18093 <= not w18085 and w18092;
w18094 <= not w18091 and not w18093;
w18095 <= w18011 and not w18094;
w18096 <= not w18011 and w18094;
w18097 <= not w18095 and not w18096;
w18098 <= a(62) and w14223;
w18099 <= w8006 and not w18098;
w18100 <= w8006 and not w18099;
w18101 <= not w18098 and not w18099;
w18102 <= not a(57) and not w13887;
w18103 <= w18101 and not w18102;
w18104 <= not w18100 and not w18103;
w18105 <= not w18097 and not w18104;
w18106 <= w18097 and w18104;
w18107 <= not w18105 and not w18106;
w18108 <= not w18083 and w18107;
w18109 <= w18083 and not w18107;
w18110 <= not w18108 and not w18109;
w18111 <= not w18082 and not w18110;
w18112 <= w18082 and w18110;
w18113 <= not w18111 and not w18112;
w18114 <= w18063 and not w18113;
w18115 <= not w18063 and w18113;
w18116 <= not w18114 and not w18115;
w18117 <= not w18062 and not w18116;
w18118 <= w18062 and w18116;
w18119 <= not w18117 and not w18118;
w18120 <= not w18062 and not w18114;
w18121 <= not w18115 and not w18120;
w18122 <= not w18108 and not w18112;
w18123 <= w18092 and w18101;
w18124 <= not w18092 and not w18101;
w18125 <= not w18123 and not w18124;
w18126 <= not w18064 and not w18070;
w18127 <= not w18125 and w18126;
w18128 <= w18125 and not w18126;
w18129 <= not w18127 and not w18128;
w18130 <= not w18076 and not w18081;
w18131 <= not w18129 and w18130;
w18132 <= w18129 and not w18130;
w18133 <= not w18131 and not w18132;
w18134 <= a(52) and a(62);
w18135 <= a(53) and a(61);
w18136 <= not w18134 and not w18135;
w18137 <= w7239 and w9527;
w18138 <= w6774 and w9598;
w18139 <= w7038 and w9715;
w18140 <= not w18138 and not w18139;
w18141 <= not w18137 and not w18140;
w18142 <= not w18137 and not w18141;
w18143 <= not w18136 and w18142;
w18144 <= a(63) and not w18141;
w18145 <= a(51) and w18144;
w18146 <= not w18143 and not w18145;
w18147 <= w8793 and w8967;
w18148 <= w7227 and w9895;
w18149 <= w7507 and w9315;
w18150 <= not w18148 and not w18149;
w18151 <= not w18147 and not w18150;
w18152 <= a(60) and not w18151;
w18153 <= a(54) and w18152;
w18154 <= not w18147 and not w18151;
w18155 <= not w7748 and not w18022;
w18156 <= w18154 and not w18155;
w18157 <= not w18153 and not w18156;
w18158 <= not w18146 and not w18157;
w18159 <= not w18146 and not w18158;
w18160 <= not w18157 and not w18158;
w18161 <= not w18159 and not w18160;
w18162 <= not w18011 and not w18094;
w18163 <= not w18105 and not w18162;
w18164 <= w18161 and w18163;
w18165 <= not w18161 and not w18163;
w18166 <= not w18164 and not w18165;
w18167 <= w18133 and w18166;
w18168 <= not w18133 and not w18166;
w18169 <= not w18167 and not w18168;
w18170 <= w18122 and not w18169;
w18171 <= not w18122 and w18169;
w18172 <= not w18170 and not w18171;
w18173 <= w18121 and not w18172;
w18174 <= not w18121 and not w18170;
w18175 <= not w18171 and w18174;
w18176 <= not w18173 and not w18175;
w18177 <= not w18171 and not w18174;
w18178 <= not w18132 and not w18167;
w18179 <= a(53) and a(62);
w18180 <= a(58) and w18179;
w18181 <= w8242 and not w18180;
w18182 <= not w18180 and not w18181;
w18183 <= not a(58) and not w18179;
w18184 <= w18182 and not w18183;
w18185 <= w8242 and not w18181;
w18186 <= not w18184 and not w18185;
w18187 <= w8967 and w9315;
w18188 <= w7227 and w8711;
w18189 <= w7507 and w9318;
w18190 <= not w18188 and not w18189;
w18191 <= not w18187 and not w18190;
w18192 <= a(61) and not w18191;
w18193 <= a(54) and w18192;
w18194 <= not w18187 and not w18191;
w18195 <= a(55) and a(60);
w18196 <= not w13676 and not w18195;
w18197 <= w18194 and not w18196;
w18198 <= not w18193 and not w18197;
w18199 <= not w18186 and not w18198;
w18200 <= not w18186 and not w18199;
w18201 <= not w18198 and not w18199;
w18202 <= not w18200 and not w18201;
w18203 <= not w18124 and not w18128;
w18204 <= w18202 and w18203;
w18205 <= not w18202 and not w18203;
w18206 <= not w18204 and not w18205;
w18207 <= a(52) and a(63);
w18208 <= not w18154 and w18207;
w18209 <= w18154 and not w18207;
w18210 <= not w18208 and not w18209;
w18211 <= w18142 and not w18210;
w18212 <= not w18142 and w18210;
w18213 <= not w18211 and not w18212;
w18214 <= not w18158 and not w18165;
w18215 <= not w18213 and w18214;
w18216 <= w18213 and not w18214;
w18217 <= not w18215 and not w18216;
w18218 <= w18206 and w18217;
w18219 <= not w18206 and not w18217;
w18220 <= not w18218 and not w18219;
w18221 <= not w18178 and w18220;
w18222 <= w18178 and not w18220;
w18223 <= not w18221 and not w18222;
w18224 <= not w18177 and not w18223;
w18225 <= w18177 and w18223;
w18226 <= not w18224 and not w18225;
w18227 <= not w18177 and not w18222;
w18228 <= not w18221 and not w18227;
w18229 <= not w18199 and not w18205;
w18230 <= not w18208 and not w18212;
w18231 <= w18229 and w18230;
w18232 <= not w18229 and not w18230;
w18233 <= not w18231 and not w18232;
w18234 <= w7505 and w9598;
w18235 <= a(62) and not w18234;
w18236 <= a(54) and w18235;
w18237 <= a(53) and not w18234;
w18238 <= a(63) and w18237;
w18239 <= not w18236 and not w18238;
w18240 <= not w18182 and not w18239;
w18241 <= not w18182 and not w18240;
w18242 <= not w18239 and not w18240;
w18243 <= not w18241 and not w18242;
w18244 <= w8006 and w9315;
w18245 <= w8711 and w11524;
w18246 <= w8967 and w9318;
w18247 <= not w18245 and not w18246;
w18248 <= not w18244 and not w18247;
w18249 <= a(55) and not w18248;
w18250 <= a(61) and w18249;
w18251 <= not w18244 and not w18248;
w18252 <= a(56) and a(60);
w18253 <= not w8791 and not w18252;
w18254 <= w18251 and not w18253;
w18255 <= not w18250 and not w18254;
w18256 <= not w18194 and not w18255;
w18257 <= not w18194 and not w18256;
w18258 <= not w18255 and not w18256;
w18259 <= not w18257 and not w18258;
w18260 <= not w18243 and not w18259;
w18261 <= w18243 and not w18258;
w18262 <= not w18257 and w18261;
w18263 <= not w18260 and not w18262;
w18264 <= w18233 and w18263;
w18265 <= not w18233 and not w18263;
w18266 <= not w18264 and not w18265;
w18267 <= not w18216 and not w18218;
w18268 <= not w18266 and w18267;
w18269 <= w18266 and not w18267;
w18270 <= not w18268 and not w18269;
w18271 <= w18228 and not w18270;
w18272 <= not w18228 and not w18268;
w18273 <= not w18269 and w18272;
w18274 <= not w18271 and not w18273;
w18275 <= not w18269 and not w18272;
w18276 <= not w18232 and not w18264;
w18277 <= not w18234 and not w18240;
w18278 <= w18251 and w18277;
w18279 <= not w18251 and not w18277;
w18280 <= not w18278 and not w18279;
w18281 <= w8006 and w9318;
w18282 <= w11440 and w13536;
w18283 <= w7227 and w9715;
w18284 <= not w18282 and not w18283;
w18285 <= not w18281 and not w18284;
w18286 <= a(63) and not w18285;
w18287 <= a(54) and w18286;
w18288 <= a(56) and a(61);
w18289 <= not w13018 and not w18288;
w18290 <= not w18281 and not w18285;
w18291 <= not w18289 and w18290;
w18292 <= not w18287 and not w18291;
w18293 <= w18280 and not w18292;
w18294 <= w18280 and not w18293;
w18295 <= not w18292 and not w18293;
w18296 <= not w18294 and not w18295;
w18297 <= not w18256 and not w18260;
w18298 <= a(55) and w16101;
w18299 <= w8793 and not w18298;
w18300 <= w8793 and not w18299;
w18301 <= not w18298 and not w18299;
w18302 <= a(55) and a(62);
w18303 <= not a(59) and not w18302;
w18304 <= w18301 and not w18303;
w18305 <= not w18300 and not w18304;
w18306 <= not w18297 and not w18305;
w18307 <= not w18297 and not w18306;
w18308 <= not w18305 and not w18306;
w18309 <= not w18307 and not w18308;
w18310 <= not w18296 and w18309;
w18311 <= w18296 and not w18309;
w18312 <= not w18310 and not w18311;
w18313 <= not w18276 and not w18312;
w18314 <= w18276 and w18312;
w18315 <= not w18313 and not w18314;
w18316 <= not w18275 and not w18315;
w18317 <= w18275 and w18315;
w18318 <= not w18316 and not w18317;
w18319 <= a(55) and a(63);
w18320 <= not w18301 and w18319;
w18321 <= w18301 and not w18319;
w18322 <= not w18320 and not w18321;
w18323 <= w18290 and not w18322;
w18324 <= not w18290 and w18322;
w18325 <= not w18323 and not w18324;
w18326 <= not w18279 and not w18293;
w18327 <= w8242 and w9318;
w18328 <= w9895 and w17958;
w18329 <= w8006 and w9527;
w18330 <= not w18328 and not w18329;
w18331 <= not w18327 and not w18330;
w18332 <= w17958 and not w18331;
w18333 <= not w18327 and not w18331;
w18334 <= a(57) and a(61);
w18335 <= not w9895 and not w18334;
w18336 <= w18333 and not w18335;
w18337 <= not w18332 and not w18336;
w18338 <= not w18326 and not w18337;
w18339 <= not w18326 and not w18338;
w18340 <= not w18337 and not w18338;
w18341 <= not w18339 and not w18340;
w18342 <= not w18325 and w18341;
w18343 <= w18325 and not w18341;
w18344 <= not w18342 and not w18343;
w18345 <= not w18296 and not w18309;
w18346 <= not w18306 and not w18345;
w18347 <= not w18344 and w18346;
w18348 <= w18344 and not w18346;
w18349 <= not w18347 and not w18348;
w18350 <= not w18275 and not w18314;
w18351 <= not w18313 and not w18350;
w18352 <= not w18349 and w18351;
w18353 <= w18349 and not w18351;
w18354 <= not w18352 and not w18353;
w18355 <= w7748 and w9715;
w18356 <= a(61) and not w18355;
w18357 <= a(58) and w18356;
w18358 <= a(56) and not w18355;
w18359 <= a(63) and w18358;
w18360 <= not w18357 and not w18359;
w18361 <= not w18333 and not w18360;
w18362 <= not w18333 and not w18361;
w18363 <= not w18360 and not w18361;
w18364 <= not w18362 and not w18363;
w18365 <= a(57) and w8891;
w18366 <= w9315 and not w18365;
w18367 <= w9315 and not w18366;
w18368 <= not w18365 and not w18366;
w18369 <= a(57) and a(62);
w18370 <= not a(60) and not w18369;
w18371 <= w18368 and not w18370;
w18372 <= not w18367 and not w18371;
w18373 <= not w18364 and not w18372;
w18374 <= not w18364 and not w18373;
w18375 <= not w18372 and not w18373;
w18376 <= not w18374 and not w18375;
w18377 <= not w18320 and not w18324;
w18378 <= w18376 and w18377;
w18379 <= not w18376 and not w18377;
w18380 <= not w18378 and not w18379;
w18381 <= not w18338 and not w18343;
w18382 <= w18380 and not w18381;
w18383 <= not w18380 and w18381;
w18384 <= not w18382 and not w18383;
w18385 <= not w18347 and not w18351;
w18386 <= not w18348 and not w18385;
w18387 <= not w18384 and w18386;
w18388 <= w18384 and not w18386;
w18389 <= not w18387 and not w18388;
w18390 <= not w18383 and not w18386;
w18391 <= not w18382 and not w18390;
w18392 <= not w18373 and not w18379;
w18393 <= not w18355 and not w18361;
w18394 <= w18368 and w18393;
w18395 <= not w18368 and not w18393;
w18396 <= not w18394 and not w18395;
w18397 <= w8793 and w9527;
w18398 <= w8791 and w9715;
w18399 <= w8242 and w9598;
w18400 <= not w18398 and not w18399;
w18401 <= not w18397 and not w18400;
w18402 <= a(63) and not w18401;
w18403 <= a(57) and w18402;
w18404 <= not w18397 and not w18401;
w18405 <= a(58) and a(62);
w18406 <= not w8711 and not w18405;
w18407 <= w18404 and not w18406;
w18408 <= not w18403 and not w18407;
w18409 <= w18396 and not w18408;
w18410 <= not w18396 and w18408;
w18411 <= not w18409 and not w18410;
w18412 <= w18392 and not w18411;
w18413 <= not w18392 and w18411;
w18414 <= not w18412 and not w18413;
w18415 <= w18391 and not w18414;
w18416 <= not w18391 and not w18412;
w18417 <= not w18413 and w18416;
w18418 <= not w18415 and not w18417;
w18419 <= not a(60) and a(61);
w18420 <= not w16101 and not w18419;
w18421 <= w16101 and w18419;
w18422 <= not w18420 and not w18421;
w18423 <= w17605 and not w18404;
w18424 <= not w17605 and w18404;
w18425 <= not w18423 and not w18424;
w18426 <= not w18422 and not w18425;
w18427 <= w18422 and w18425;
w18428 <= not w18426 and not w18427;
w18429 <= not w18395 and not w18409;
w18430 <= not w18428 and w18429;
w18431 <= w18428 and not w18429;
w18432 <= not w18430 and not w18431;
w18433 <= not w18413 and not w18416;
w18434 <= not w18432 and w18433;
w18435 <= w18432 and not w18433;
w18436 <= not w18434 and not w18435;
w18437 <= not w18430 and not w18433;
w18438 <= not w18431 and not w18437;
w18439 <= not w8891 and not w17608;
w18440 <= w9315 and w9598;
w18441 <= not w9318 and not w18421;
w18442 <= not w18440 and not w18441;
w18443 <= not w18439 and w18442;
w18444 <= not w18440 and not w18443;
w18445 <= not w18439 and w18444;
w18446 <= not w18441 and not w18443;
w18447 <= not w18445 and not w18446;
w18448 <= not w18423 and not w18427;
w18449 <= w18447 and w18448;
w18450 <= not w18447 and not w18448;
w18451 <= not w18449 and not w18450;
w18452 <= w18438 and not w18451;
w18453 <= not w18438 and not w18449;
w18454 <= not w18450 and w18453;
w18455 <= not w18452 and not w18454;
w18456 <= not a(61) and a(62);
w18457 <= not w11440 and not w18456;
w18458 <= w11440 and w18456;
w18459 <= not w18457 and not w18458;
w18460 <= w18444 and not w18459;
w18461 <= not w18444 and w18459;
w18462 <= not w18460 and not w18461;
w18463 <= not w18450 and not w18453;
w18464 <= not w18462 and w18463;
w18465 <= w18462 and not w18463;
w18466 <= not w18464 and not w18465;
w18467 <= not w18460 and not w18463;
w18468 <= not w18461 and not w18467;
w18469 <= a(62) and w9715;
w18470 <= not w9527 and not w9715;
w18471 <= not w18458 and w18470;
w18472 <= not w18469 and not w18471;
w18473 <= not w18468 and w18472;
w18474 <= w18468 and not w18472;
w18475 <= not w18473 and not w18474;
w18476 <= not a(62) and a(63);
w18477 <= not w18468 and not w18471;
w18478 <= not w18469 and not w18477;
w18479 <= not w18476 and w18478;
w18480 <= w18476 and not w18478;
w18481 <= not w18479 and not w18480;
w18482 <= a(63) and not w18478;
w18483 <= not w9598 and not w18482;
one <= '1';
asquared(0) <= a(0);-- level 0
asquared(1) <= not one;-- level 0
asquared(2) <= w1;-- level 2
asquared(3) <= w5;-- level 3
asquared(4) <= not w14;-- level 6
asquared(5) <= w28;-- level 7
asquared(6) <= w48;-- level 11
asquared(7) <= w70;-- level 13
asquared(8) <= w103;-- level 15
asquared(9) <= w136;-- level 16
asquared(10) <= w180;-- level 18
asquared(11) <= w226;-- level 21
asquared(12) <= w278;-- level 22
asquared(13) <= w331;-- level 25
asquared(14) <= w386;-- level 26
asquared(15) <= w451;-- level 29
asquared(16) <= not w521;-- level 30
asquared(17) <= w596;-- level 32
asquared(18) <= w678;-- level 34
asquared(19) <= w762;-- level 37
asquared(20) <= w849;-- level 38
asquared(21) <= w942;-- level 40
asquared(22) <= w1038;-- level 42
asquared(23) <= w1134;-- level 45
asquared(24) <= w1236;-- level 46
asquared(25) <= w1348;-- level 49
asquared(26) <= w1465;-- level 50
asquared(27) <= w1585;-- level 52
asquared(28) <= w1705;-- level 54
asquared(29) <= w1831;-- level 56
asquared(30) <= w1969;-- level 58
asquared(31) <= w2103;-- level 60
asquared(32) <= w2251;-- level 62
asquared(33) <= w2391;-- level 64
asquared(34) <= w2547;-- level 66
asquared(35) <= w2703;-- level 69
asquared(36) <= not w2862;-- level 70
asquared(37) <= w3029;-- level 72
asquared(38) <= w3206;-- level 74
asquared(39) <= w3381;-- level 76
asquared(40) <= w3563;-- level 78
asquared(41) <= w3744;-- level 81
asquared(42) <= w3933;-- level 82
asquared(43) <= w4129;-- level 84
asquared(44) <= w4333;-- level 86
asquared(45) <= w4536;-- level 88
asquared(46) <= w4754;-- level 90
asquared(47) <= w4960;-- level 92
asquared(48) <= w5197;-- level 94
asquared(49) <= w5421;-- level 97
asquared(50) <= w5647;-- level 98
asquared(51) <= w5882;-- level 101
asquared(52) <= not w6122;-- level 102
asquared(53) <= w6362;-- level 105
asquared(54) <= not w6605;-- level 106
asquared(55) <= w6859;-- level 108
asquared(56) <= w7125;-- level 110
asquared(57) <= w7391;-- level 112
asquared(58) <= w7664;-- level 114
asquared(59) <= w7927;-- level 117
asquared(60) <= w8207;-- level 118
asquared(61) <= w8489;-- level 120
asquared(62) <= w8782;-- level 122
asquared(63) <= w9076;-- level 125
asquared(64) <= not w9374;-- level 126
asquared(65) <= w9664;-- level 129
asquared(66) <= not w9954;-- level 130
asquared(67) <= w10237;-- level 132
asquared(68) <= w10516;-- level 134
asquared(69) <= w10783;-- level 136
asquared(70) <= w11053;-- level 138
asquared(71) <= w11322;-- level 141
asquared(72) <= not w11576;-- level 142
asquared(73) <= w11823;-- level 145
asquared(74) <= not w12071;-- level 146
asquared(75) <= w12307;-- level 148
asquared(76) <= w12552;-- level 150
asquared(77) <= w12781;-- level 152
asquared(78) <= w13010;-- level 154
asquared(79) <= w13233;-- level 156
asquared(80) <= w13452;-- level 158
asquared(81) <= w13661;-- level 161
asquared(82) <= not w13879;-- level 162
asquared(83) <= w14084;-- level 164
asquared(84) <= w14289;-- level 166
asquared(85) <= w14487;-- level 168
asquared(86) <= not w14683;-- level 170
asquared(87) <= w14862;-- level 173
asquared(88) <= not w15045;-- level 174
asquared(89) <= w15216;-- level 176
asquared(90) <= w15391;-- level 178
asquared(91) <= w15561;-- level 181
asquared(92) <= not w15726;-- level 182
asquared(93) <= w15882;-- level 185
asquared(94) <= not w16033;-- level 186
asquared(95) <= w16175;-- level 188
asquared(96) <= w16322;-- level 190
asquared(97) <= w16464;-- level 193
asquared(98) <= not w16598;-- level 194
asquared(99) <= w16723;-- level 196
asquared(100) <= w16853;-- level 198
asquared(101) <= w16965;-- level 201
asquared(102) <= not w17085;-- level 202
asquared(103) <= w17201;-- level 205
asquared(104) <= not w17308;-- level 206
asquared(105) <= w17408;-- level 208
asquared(106) <= w17506;-- level 210
asquared(107) <= w17597;-- level 213
asquared(108) <= not w17686;-- level 214
asquared(109) <= w17772;-- level 217
asquared(110) <= not w17851;-- level 218
asquared(111) <= w17927;-- level 221
asquared(112) <= not w17998;-- level 222
asquared(113) <= w18061;-- level 225
asquared(114) <= not w18119;-- level 226
asquared(115) <= w18176;-- level 229
asquared(116) <= not w18226;-- level 230
asquared(117) <= w18274;-- level 233
asquared(118) <= not w18318;-- level 234
asquared(119) <= w18354;-- level 236
asquared(120) <= w18389;-- level 238
asquared(121) <= w18418;-- level 241
asquared(122) <= w18436;-- level 242
asquared(123) <= w18455;-- level 245
asquared(124) <= w18466;-- level 246
asquared(125) <= w18475;-- level 248
asquared(126) <= w18481;-- level 250
asquared(127) <= not w18483;-- level 250
end Behavioral;