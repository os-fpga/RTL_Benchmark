.INIT({   1'b0, INIT[2047*8 +: 8], 1'b0, INIT[2046*8 +: 8], 1'b0, INIT[2043*8 +: 8], 1'b0, INIT[2042*8 +: 8], 
          1'b0, INIT[2039*8 +: 8], 1'b0, INIT[2038*8 +: 8], 1'b0, INIT[2035*8 +: 8], 1'b0, INIT[2034*8 +: 8], 
          1'b0, INIT[2031*8 +: 8], 1'b0, INIT[2030*8 +: 8], 1'b0, INIT[2027*8 +: 8], 1'b0, INIT[2026*8 +: 8], 
          1'b0, INIT[2023*8 +: 8], 1'b0, INIT[2022*8 +: 8], 1'b0, INIT[2019*8 +: 8], 1'b0, INIT[2018*8 +: 8], 
          1'b0, INIT[2015*8 +: 8], 1'b0, INIT[2014*8 +: 8], 1'b0, INIT[2011*8 +: 8], 1'b0, INIT[2010*8 +: 8], 
          1'b0, INIT[2007*8 +: 8], 1'b0, INIT[2006*8 +: 8], 1'b0, INIT[2003*8 +: 8], 1'b0, INIT[2002*8 +: 8], 
          1'b0, INIT[1999*8 +: 8], 1'b0, INIT[1998*8 +: 8], 1'b0, INIT[1995*8 +: 8], 1'b0, INIT[1994*8 +: 8], 
          1'b0, INIT[1991*8 +: 8], 1'b0, INIT[1990*8 +: 8], 1'b0, INIT[1987*8 +: 8], 1'b0, INIT[1986*8 +: 8], 
          1'b0, INIT[1983*8 +: 8], 1'b0, INIT[1982*8 +: 8], 1'b0, INIT[1979*8 +: 8], 1'b0, INIT[1978*8 +: 8], 
          1'b0, INIT[1975*8 +: 8], 1'b0, INIT[1974*8 +: 8], 1'b0, INIT[1971*8 +: 8], 1'b0, INIT[1970*8 +: 8], 
          1'b0, INIT[1967*8 +: 8], 1'b0, INIT[1966*8 +: 8], 1'b0, INIT[1963*8 +: 8], 1'b0, INIT[1962*8 +: 8], 
          1'b0, INIT[1959*8 +: 8], 1'b0, INIT[1958*8 +: 8], 1'b0, INIT[1955*8 +: 8], 1'b0, INIT[1954*8 +: 8], 
          1'b0, INIT[1951*8 +: 8], 1'b0, INIT[1950*8 +: 8], 1'b0, INIT[1947*8 +: 8], 1'b0, INIT[1946*8 +: 8], 
          1'b0, INIT[1943*8 +: 8], 1'b0, INIT[1942*8 +: 8], 1'b0, INIT[1939*8 +: 8], 1'b0, INIT[1938*8 +: 8], 
          1'b0, INIT[1935*8 +: 8], 1'b0, INIT[1934*8 +: 8], 1'b0, INIT[1931*8 +: 8], 1'b0, INIT[1930*8 +: 8], 
          1'b0, INIT[1927*8 +: 8], 1'b0, INIT[1926*8 +: 8], 1'b0, INIT[1923*8 +: 8], 1'b0, INIT[1922*8 +: 8], 
          1'b0, INIT[1919*8 +: 8], 1'b0, INIT[1918*8 +: 8], 1'b0, INIT[1915*8 +: 8], 1'b0, INIT[1914*8 +: 8], 
          1'b0, INIT[1911*8 +: 8], 1'b0, INIT[1910*8 +: 8], 1'b0, INIT[1907*8 +: 8], 1'b0, INIT[1906*8 +: 8], 
          1'b0, INIT[1903*8 +: 8], 1'b0, INIT[1902*8 +: 8], 1'b0, INIT[1899*8 +: 8], 1'b0, INIT[1898*8 +: 8], 
          1'b0, INIT[1895*8 +: 8], 1'b0, INIT[1894*8 +: 8], 1'b0, INIT[1891*8 +: 8], 1'b0, INIT[1890*8 +: 8], 
          1'b0, INIT[1887*8 +: 8], 1'b0, INIT[1886*8 +: 8], 1'b0, INIT[1883*8 +: 8], 1'b0, INIT[1882*8 +: 8], 
          1'b0, INIT[1879*8 +: 8], 1'b0, INIT[1878*8 +: 8], 1'b0, INIT[1875*8 +: 8], 1'b0, INIT[1874*8 +: 8], 
          1'b0, INIT[1871*8 +: 8], 1'b0, INIT[1870*8 +: 8], 1'b0, INIT[1867*8 +: 8], 1'b0, INIT[1866*8 +: 8], 
          1'b0, INIT[1863*8 +: 8], 1'b0, INIT[1862*8 +: 8], 1'b0, INIT[1859*8 +: 8], 1'b0, INIT[1858*8 +: 8], 
          1'b0, INIT[1855*8 +: 8], 1'b0, INIT[1854*8 +: 8], 1'b0, INIT[1851*8 +: 8], 1'b0, INIT[1850*8 +: 8], 
          1'b0, INIT[1847*8 +: 8], 1'b0, INIT[1846*8 +: 8], 1'b0, INIT[1843*8 +: 8], 1'b0, INIT[1842*8 +: 8], 
          1'b0, INIT[1839*8 +: 8], 1'b0, INIT[1838*8 +: 8], 1'b0, INIT[1835*8 +: 8], 1'b0, INIT[1834*8 +: 8], 
          1'b0, INIT[1831*8 +: 8], 1'b0, INIT[1830*8 +: 8], 1'b0, INIT[1827*8 +: 8], 1'b0, INIT[1826*8 +: 8], 
          1'b0, INIT[1823*8 +: 8], 1'b0, INIT[1822*8 +: 8], 1'b0, INIT[1819*8 +: 8], 1'b0, INIT[1818*8 +: 8], 
          1'b0, INIT[1815*8 +: 8], 1'b0, INIT[1814*8 +: 8], 1'b0, INIT[1811*8 +: 8], 1'b0, INIT[1810*8 +: 8], 
          1'b0, INIT[1807*8 +: 8], 1'b0, INIT[1806*8 +: 8], 1'b0, INIT[1803*8 +: 8], 1'b0, INIT[1802*8 +: 8], 
          1'b0, INIT[1799*8 +: 8], 1'b0, INIT[1798*8 +: 8], 1'b0, INIT[1795*8 +: 8], 1'b0, INIT[1794*8 +: 8], 
          1'b0, INIT[1791*8 +: 8], 1'b0, INIT[1790*8 +: 8], 1'b0, INIT[1787*8 +: 8], 1'b0, INIT[1786*8 +: 8], 
          1'b0, INIT[1783*8 +: 8], 1'b0, INIT[1782*8 +: 8], 1'b0, INIT[1779*8 +: 8], 1'b0, INIT[1778*8 +: 8], 
          1'b0, INIT[1775*8 +: 8], 1'b0, INIT[1774*8 +: 8], 1'b0, INIT[1771*8 +: 8], 1'b0, INIT[1770*8 +: 8], 
          1'b0, INIT[1767*8 +: 8], 1'b0, INIT[1766*8 +: 8], 1'b0, INIT[1763*8 +: 8], 1'b0, INIT[1762*8 +: 8], 
          1'b0, INIT[1759*8 +: 8], 1'b0, INIT[1758*8 +: 8], 1'b0, INIT[1755*8 +: 8], 1'b0, INIT[1754*8 +: 8], 
          1'b0, INIT[1751*8 +: 8], 1'b0, INIT[1750*8 +: 8], 1'b0, INIT[1747*8 +: 8], 1'b0, INIT[1746*8 +: 8], 
          1'b0, INIT[1743*8 +: 8], 1'b0, INIT[1742*8 +: 8], 1'b0, INIT[1739*8 +: 8], 1'b0, INIT[1738*8 +: 8], 
          1'b0, INIT[1735*8 +: 8], 1'b0, INIT[1734*8 +: 8], 1'b0, INIT[1731*8 +: 8], 1'b0, INIT[1730*8 +: 8], 
          1'b0, INIT[1727*8 +: 8], 1'b0, INIT[1726*8 +: 8], 1'b0, INIT[1723*8 +: 8], 1'b0, INIT[1722*8 +: 8], 
          1'b0, INIT[1719*8 +: 8], 1'b0, INIT[1718*8 +: 8], 1'b0, INIT[1715*8 +: 8], 1'b0, INIT[1714*8 +: 8], 
          1'b0, INIT[1711*8 +: 8], 1'b0, INIT[1710*8 +: 8], 1'b0, INIT[1707*8 +: 8], 1'b0, INIT[1706*8 +: 8], 
          1'b0, INIT[1703*8 +: 8], 1'b0, INIT[1702*8 +: 8], 1'b0, INIT[1699*8 +: 8], 1'b0, INIT[1698*8 +: 8], 
          1'b0, INIT[1695*8 +: 8], 1'b0, INIT[1694*8 +: 8], 1'b0, INIT[1691*8 +: 8], 1'b0, INIT[1690*8 +: 8], 
          1'b0, INIT[1687*8 +: 8], 1'b0, INIT[1686*8 +: 8], 1'b0, INIT[1683*8 +: 8], 1'b0, INIT[1682*8 +: 8], 
          1'b0, INIT[1679*8 +: 8], 1'b0, INIT[1678*8 +: 8], 1'b0, INIT[1675*8 +: 8], 1'b0, INIT[1674*8 +: 8], 
          1'b0, INIT[1671*8 +: 8], 1'b0, INIT[1670*8 +: 8], 1'b0, INIT[1667*8 +: 8], 1'b0, INIT[1666*8 +: 8], 
          1'b0, INIT[1663*8 +: 8], 1'b0, INIT[1662*8 +: 8], 1'b0, INIT[1659*8 +: 8], 1'b0, INIT[1658*8 +: 8], 
          1'b0, INIT[1655*8 +: 8], 1'b0, INIT[1654*8 +: 8], 1'b0, INIT[1651*8 +: 8], 1'b0, INIT[1650*8 +: 8], 
          1'b0, INIT[1647*8 +: 8], 1'b0, INIT[1646*8 +: 8], 1'b0, INIT[1643*8 +: 8], 1'b0, INIT[1642*8 +: 8], 
          1'b0, INIT[1639*8 +: 8], 1'b0, INIT[1638*8 +: 8], 1'b0, INIT[1635*8 +: 8], 1'b0, INIT[1634*8 +: 8], 
          1'b0, INIT[1631*8 +: 8], 1'b0, INIT[1630*8 +: 8], 1'b0, INIT[1627*8 +: 8], 1'b0, INIT[1626*8 +: 8], 
          1'b0, INIT[1623*8 +: 8], 1'b0, INIT[1622*8 +: 8], 1'b0, INIT[1619*8 +: 8], 1'b0, INIT[1618*8 +: 8], 
          1'b0, INIT[1615*8 +: 8], 1'b0, INIT[1614*8 +: 8], 1'b0, INIT[1611*8 +: 8], 1'b0, INIT[1610*8 +: 8], 
          1'b0, INIT[1607*8 +: 8], 1'b0, INIT[1606*8 +: 8], 1'b0, INIT[1603*8 +: 8], 1'b0, INIT[1602*8 +: 8], 
          1'b0, INIT[1599*8 +: 8], 1'b0, INIT[1598*8 +: 8], 1'b0, INIT[1595*8 +: 8], 1'b0, INIT[1594*8 +: 8], 
          1'b0, INIT[1591*8 +: 8], 1'b0, INIT[1590*8 +: 8], 1'b0, INIT[1587*8 +: 8], 1'b0, INIT[1586*8 +: 8], 
          1'b0, INIT[1583*8 +: 8], 1'b0, INIT[1582*8 +: 8], 1'b0, INIT[1579*8 +: 8], 1'b0, INIT[1578*8 +: 8], 
          1'b0, INIT[1575*8 +: 8], 1'b0, INIT[1574*8 +: 8], 1'b0, INIT[1571*8 +: 8], 1'b0, INIT[1570*8 +: 8], 
          1'b0, INIT[1567*8 +: 8], 1'b0, INIT[1566*8 +: 8], 1'b0, INIT[1563*8 +: 8], 1'b0, INIT[1562*8 +: 8], 
          1'b0, INIT[1559*8 +: 8], 1'b0, INIT[1558*8 +: 8], 1'b0, INIT[1555*8 +: 8], 1'b0, INIT[1554*8 +: 8], 
          1'b0, INIT[1551*8 +: 8], 1'b0, INIT[1550*8 +: 8], 1'b0, INIT[1547*8 +: 8], 1'b0, INIT[1546*8 +: 8], 
          1'b0, INIT[1543*8 +: 8], 1'b0, INIT[1542*8 +: 8], 1'b0, INIT[1539*8 +: 8], 1'b0, INIT[1538*8 +: 8], 
          1'b0, INIT[1535*8 +: 8], 1'b0, INIT[1534*8 +: 8], 1'b0, INIT[1531*8 +: 8], 1'b0, INIT[1530*8 +: 8], 
          1'b0, INIT[1527*8 +: 8], 1'b0, INIT[1526*8 +: 8], 1'b0, INIT[1523*8 +: 8], 1'b0, INIT[1522*8 +: 8], 
          1'b0, INIT[1519*8 +: 8], 1'b0, INIT[1518*8 +: 8], 1'b0, INIT[1515*8 +: 8], 1'b0, INIT[1514*8 +: 8], 
          1'b0, INIT[1511*8 +: 8], 1'b0, INIT[1510*8 +: 8], 1'b0, INIT[1507*8 +: 8], 1'b0, INIT[1506*8 +: 8], 
          1'b0, INIT[1503*8 +: 8], 1'b0, INIT[1502*8 +: 8], 1'b0, INIT[1499*8 +: 8], 1'b0, INIT[1498*8 +: 8], 
          1'b0, INIT[1495*8 +: 8], 1'b0, INIT[1494*8 +: 8], 1'b0, INIT[1491*8 +: 8], 1'b0, INIT[1490*8 +: 8], 
          1'b0, INIT[1487*8 +: 8], 1'b0, INIT[1486*8 +: 8], 1'b0, INIT[1483*8 +: 8], 1'b0, INIT[1482*8 +: 8], 
          1'b0, INIT[1479*8 +: 8], 1'b0, INIT[1478*8 +: 8], 1'b0, INIT[1475*8 +: 8], 1'b0, INIT[1474*8 +: 8], 
          1'b0, INIT[1471*8 +: 8], 1'b0, INIT[1470*8 +: 8], 1'b0, INIT[1467*8 +: 8], 1'b0, INIT[1466*8 +: 8], 
          1'b0, INIT[1463*8 +: 8], 1'b0, INIT[1462*8 +: 8], 1'b0, INIT[1459*8 +: 8], 1'b0, INIT[1458*8 +: 8], 
          1'b0, INIT[1455*8 +: 8], 1'b0, INIT[1454*8 +: 8], 1'b0, INIT[1451*8 +: 8], 1'b0, INIT[1450*8 +: 8], 
          1'b0, INIT[1447*8 +: 8], 1'b0, INIT[1446*8 +: 8], 1'b0, INIT[1443*8 +: 8], 1'b0, INIT[1442*8 +: 8], 
          1'b0, INIT[1439*8 +: 8], 1'b0, INIT[1438*8 +: 8], 1'b0, INIT[1435*8 +: 8], 1'b0, INIT[1434*8 +: 8], 
          1'b0, INIT[1431*8 +: 8], 1'b0, INIT[1430*8 +: 8], 1'b0, INIT[1427*8 +: 8], 1'b0, INIT[1426*8 +: 8], 
          1'b0, INIT[1423*8 +: 8], 1'b0, INIT[1422*8 +: 8], 1'b0, INIT[1419*8 +: 8], 1'b0, INIT[1418*8 +: 8], 
          1'b0, INIT[1415*8 +: 8], 1'b0, INIT[1414*8 +: 8], 1'b0, INIT[1411*8 +: 8], 1'b0, INIT[1410*8 +: 8], 
          1'b0, INIT[1407*8 +: 8], 1'b0, INIT[1406*8 +: 8], 1'b0, INIT[1403*8 +: 8], 1'b0, INIT[1402*8 +: 8], 
          1'b0, INIT[1399*8 +: 8], 1'b0, INIT[1398*8 +: 8], 1'b0, INIT[1395*8 +: 8], 1'b0, INIT[1394*8 +: 8], 
          1'b0, INIT[1391*8 +: 8], 1'b0, INIT[1390*8 +: 8], 1'b0, INIT[1387*8 +: 8], 1'b0, INIT[1386*8 +: 8], 
          1'b0, INIT[1383*8 +: 8], 1'b0, INIT[1382*8 +: 8], 1'b0, INIT[1379*8 +: 8], 1'b0, INIT[1378*8 +: 8], 
          1'b0, INIT[1375*8 +: 8], 1'b0, INIT[1374*8 +: 8], 1'b0, INIT[1371*8 +: 8], 1'b0, INIT[1370*8 +: 8], 
          1'b0, INIT[1367*8 +: 8], 1'b0, INIT[1366*8 +: 8], 1'b0, INIT[1363*8 +: 8], 1'b0, INIT[1362*8 +: 8], 
          1'b0, INIT[1359*8 +: 8], 1'b0, INIT[1358*8 +: 8], 1'b0, INIT[1355*8 +: 8], 1'b0, INIT[1354*8 +: 8], 
          1'b0, INIT[1351*8 +: 8], 1'b0, INIT[1350*8 +: 8], 1'b0, INIT[1347*8 +: 8], 1'b0, INIT[1346*8 +: 8], 
          1'b0, INIT[1343*8 +: 8], 1'b0, INIT[1342*8 +: 8], 1'b0, INIT[1339*8 +: 8], 1'b0, INIT[1338*8 +: 8], 
          1'b0, INIT[1335*8 +: 8], 1'b0, INIT[1334*8 +: 8], 1'b0, INIT[1331*8 +: 8], 1'b0, INIT[1330*8 +: 8], 
          1'b0, INIT[1327*8 +: 8], 1'b0, INIT[1326*8 +: 8], 1'b0, INIT[1323*8 +: 8], 1'b0, INIT[1322*8 +: 8], 
          1'b0, INIT[1319*8 +: 8], 1'b0, INIT[1318*8 +: 8], 1'b0, INIT[1315*8 +: 8], 1'b0, INIT[1314*8 +: 8], 
          1'b0, INIT[1311*8 +: 8], 1'b0, INIT[1310*8 +: 8], 1'b0, INIT[1307*8 +: 8], 1'b0, INIT[1306*8 +: 8], 
          1'b0, INIT[1303*8 +: 8], 1'b0, INIT[1302*8 +: 8], 1'b0, INIT[1299*8 +: 8], 1'b0, INIT[1298*8 +: 8], 
          1'b0, INIT[1295*8 +: 8], 1'b0, INIT[1294*8 +: 8], 1'b0, INIT[1291*8 +: 8], 1'b0, INIT[1290*8 +: 8], 
          1'b0, INIT[1287*8 +: 8], 1'b0, INIT[1286*8 +: 8], 1'b0, INIT[1283*8 +: 8], 1'b0, INIT[1282*8 +: 8], 
          1'b0, INIT[1279*8 +: 8], 1'b0, INIT[1278*8 +: 8], 1'b0, INIT[1275*8 +: 8], 1'b0, INIT[1274*8 +: 8], 
          1'b0, INIT[1271*8 +: 8], 1'b0, INIT[1270*8 +: 8], 1'b0, INIT[1267*8 +: 8], 1'b0, INIT[1266*8 +: 8], 
          1'b0, INIT[1263*8 +: 8], 1'b0, INIT[1262*8 +: 8], 1'b0, INIT[1259*8 +: 8], 1'b0, INIT[1258*8 +: 8], 
          1'b0, INIT[1255*8 +: 8], 1'b0, INIT[1254*8 +: 8], 1'b0, INIT[1251*8 +: 8], 1'b0, INIT[1250*8 +: 8], 
          1'b0, INIT[1247*8 +: 8], 1'b0, INIT[1246*8 +: 8], 1'b0, INIT[1243*8 +: 8], 1'b0, INIT[1242*8 +: 8], 
          1'b0, INIT[1239*8 +: 8], 1'b0, INIT[1238*8 +: 8], 1'b0, INIT[1235*8 +: 8], 1'b0, INIT[1234*8 +: 8], 
          1'b0, INIT[1231*8 +: 8], 1'b0, INIT[1230*8 +: 8], 1'b0, INIT[1227*8 +: 8], 1'b0, INIT[1226*8 +: 8], 
          1'b0, INIT[1223*8 +: 8], 1'b0, INIT[1222*8 +: 8], 1'b0, INIT[1219*8 +: 8], 1'b0, INIT[1218*8 +: 8], 
          1'b0, INIT[1215*8 +: 8], 1'b0, INIT[1214*8 +: 8], 1'b0, INIT[1211*8 +: 8], 1'b0, INIT[1210*8 +: 8], 
          1'b0, INIT[1207*8 +: 8], 1'b0, INIT[1206*8 +: 8], 1'b0, INIT[1203*8 +: 8], 1'b0, INIT[1202*8 +: 8], 
          1'b0, INIT[1199*8 +: 8], 1'b0, INIT[1198*8 +: 8], 1'b0, INIT[1195*8 +: 8], 1'b0, INIT[1194*8 +: 8], 
          1'b0, INIT[1191*8 +: 8], 1'b0, INIT[1190*8 +: 8], 1'b0, INIT[1187*8 +: 8], 1'b0, INIT[1186*8 +: 8], 
          1'b0, INIT[1183*8 +: 8], 1'b0, INIT[1182*8 +: 8], 1'b0, INIT[1179*8 +: 8], 1'b0, INIT[1178*8 +: 8], 
          1'b0, INIT[1175*8 +: 8], 1'b0, INIT[1174*8 +: 8], 1'b0, INIT[1171*8 +: 8], 1'b0, INIT[1170*8 +: 8], 
          1'b0, INIT[1167*8 +: 8], 1'b0, INIT[1166*8 +: 8], 1'b0, INIT[1163*8 +: 8], 1'b0, INIT[1162*8 +: 8], 
          1'b0, INIT[1159*8 +: 8], 1'b0, INIT[1158*8 +: 8], 1'b0, INIT[1155*8 +: 8], 1'b0, INIT[1154*8 +: 8], 
          1'b0, INIT[1151*8 +: 8], 1'b0, INIT[1150*8 +: 8], 1'b0, INIT[1147*8 +: 8], 1'b0, INIT[1146*8 +: 8], 
          1'b0, INIT[1143*8 +: 8], 1'b0, INIT[1142*8 +: 8], 1'b0, INIT[1139*8 +: 8], 1'b0, INIT[1138*8 +: 8], 
          1'b0, INIT[1135*8 +: 8], 1'b0, INIT[1134*8 +: 8], 1'b0, INIT[1131*8 +: 8], 1'b0, INIT[1130*8 +: 8], 
          1'b0, INIT[1127*8 +: 8], 1'b0, INIT[1126*8 +: 8], 1'b0, INIT[1123*8 +: 8], 1'b0, INIT[1122*8 +: 8], 
          1'b0, INIT[1119*8 +: 8], 1'b0, INIT[1118*8 +: 8], 1'b0, INIT[1115*8 +: 8], 1'b0, INIT[1114*8 +: 8], 
          1'b0, INIT[1111*8 +: 8], 1'b0, INIT[1110*8 +: 8], 1'b0, INIT[1107*8 +: 8], 1'b0, INIT[1106*8 +: 8], 
          1'b0, INIT[1103*8 +: 8], 1'b0, INIT[1102*8 +: 8], 1'b0, INIT[1099*8 +: 8], 1'b0, INIT[1098*8 +: 8], 
          1'b0, INIT[1095*8 +: 8], 1'b0, INIT[1094*8 +: 8], 1'b0, INIT[1091*8 +: 8], 1'b0, INIT[1090*8 +: 8], 
          1'b0, INIT[1087*8 +: 8], 1'b0, INIT[1086*8 +: 8], 1'b0, INIT[1083*8 +: 8], 1'b0, INIT[1082*8 +: 8], 
          1'b0, INIT[1079*8 +: 8], 1'b0, INIT[1078*8 +: 8], 1'b0, INIT[1075*8 +: 8], 1'b0, INIT[1074*8 +: 8], 
          1'b0, INIT[1071*8 +: 8], 1'b0, INIT[1070*8 +: 8], 1'b0, INIT[1067*8 +: 8], 1'b0, INIT[1066*8 +: 8], 
          1'b0, INIT[1063*8 +: 8], 1'b0, INIT[1062*8 +: 8], 1'b0, INIT[1059*8 +: 8], 1'b0, INIT[1058*8 +: 8], 
          1'b0, INIT[1055*8 +: 8], 1'b0, INIT[1054*8 +: 8], 1'b0, INIT[1051*8 +: 8], 1'b0, INIT[1050*8 +: 8], 
          1'b0, INIT[1047*8 +: 8], 1'b0, INIT[1046*8 +: 8], 1'b0, INIT[1043*8 +: 8], 1'b0, INIT[1042*8 +: 8], 
          1'b0, INIT[1039*8 +: 8], 1'b0, INIT[1038*8 +: 8], 1'b0, INIT[1035*8 +: 8], 1'b0, INIT[1034*8 +: 8], 
          1'b0, INIT[1031*8 +: 8], 1'b0, INIT[1030*8 +: 8], 1'b0, INIT[1027*8 +: 8], 1'b0, INIT[1026*8 +: 8], 
          1'b0, INIT[1023*8 +: 8], 1'b0, INIT[1022*8 +: 8], 1'b0, INIT[1019*8 +: 8], 1'b0, INIT[1018*8 +: 8], 
          1'b0, INIT[1015*8 +: 8], 1'b0, INIT[1014*8 +: 8], 1'b0, INIT[1011*8 +: 8], 1'b0, INIT[1010*8 +: 8], 
          1'b0, INIT[1007*8 +: 8], 1'b0, INIT[1006*8 +: 8], 1'b0, INIT[1003*8 +: 8], 1'b0, INIT[1002*8 +: 8], 
          1'b0, INIT[ 999*8 +: 8], 1'b0, INIT[ 998*8 +: 8], 1'b0, INIT[ 995*8 +: 8], 1'b0, INIT[ 994*8 +: 8], 
          1'b0, INIT[ 991*8 +: 8], 1'b0, INIT[ 990*8 +: 8], 1'b0, INIT[ 987*8 +: 8], 1'b0, INIT[ 986*8 +: 8], 
          1'b0, INIT[ 983*8 +: 8], 1'b0, INIT[ 982*8 +: 8], 1'b0, INIT[ 979*8 +: 8], 1'b0, INIT[ 978*8 +: 8], 
          1'b0, INIT[ 975*8 +: 8], 1'b0, INIT[ 974*8 +: 8], 1'b0, INIT[ 971*8 +: 8], 1'b0, INIT[ 970*8 +: 8], 
          1'b0, INIT[ 967*8 +: 8], 1'b0, INIT[ 966*8 +: 8], 1'b0, INIT[ 963*8 +: 8], 1'b0, INIT[ 962*8 +: 8], 
          1'b0, INIT[ 959*8 +: 8], 1'b0, INIT[ 958*8 +: 8], 1'b0, INIT[ 955*8 +: 8], 1'b0, INIT[ 954*8 +: 8], 
          1'b0, INIT[ 951*8 +: 8], 1'b0, INIT[ 950*8 +: 8], 1'b0, INIT[ 947*8 +: 8], 1'b0, INIT[ 946*8 +: 8], 
          1'b0, INIT[ 943*8 +: 8], 1'b0, INIT[ 942*8 +: 8], 1'b0, INIT[ 939*8 +: 8], 1'b0, INIT[ 938*8 +: 8], 
          1'b0, INIT[ 935*8 +: 8], 1'b0, INIT[ 934*8 +: 8], 1'b0, INIT[ 931*8 +: 8], 1'b0, INIT[ 930*8 +: 8], 
          1'b0, INIT[ 927*8 +: 8], 1'b0, INIT[ 926*8 +: 8], 1'b0, INIT[ 923*8 +: 8], 1'b0, INIT[ 922*8 +: 8], 
          1'b0, INIT[ 919*8 +: 8], 1'b0, INIT[ 918*8 +: 8], 1'b0, INIT[ 915*8 +: 8], 1'b0, INIT[ 914*8 +: 8], 
          1'b0, INIT[ 911*8 +: 8], 1'b0, INIT[ 910*8 +: 8], 1'b0, INIT[ 907*8 +: 8], 1'b0, INIT[ 906*8 +: 8], 
          1'b0, INIT[ 903*8 +: 8], 1'b0, INIT[ 902*8 +: 8], 1'b0, INIT[ 899*8 +: 8], 1'b0, INIT[ 898*8 +: 8], 
          1'b0, INIT[ 895*8 +: 8], 1'b0, INIT[ 894*8 +: 8], 1'b0, INIT[ 891*8 +: 8], 1'b0, INIT[ 890*8 +: 8], 
          1'b0, INIT[ 887*8 +: 8], 1'b0, INIT[ 886*8 +: 8], 1'b0, INIT[ 883*8 +: 8], 1'b0, INIT[ 882*8 +: 8], 
          1'b0, INIT[ 879*8 +: 8], 1'b0, INIT[ 878*8 +: 8], 1'b0, INIT[ 875*8 +: 8], 1'b0, INIT[ 874*8 +: 8], 
          1'b0, INIT[ 871*8 +: 8], 1'b0, INIT[ 870*8 +: 8], 1'b0, INIT[ 867*8 +: 8], 1'b0, INIT[ 866*8 +: 8], 
          1'b0, INIT[ 863*8 +: 8], 1'b0, INIT[ 862*8 +: 8], 1'b0, INIT[ 859*8 +: 8], 1'b0, INIT[ 858*8 +: 8], 
          1'b0, INIT[ 855*8 +: 8], 1'b0, INIT[ 854*8 +: 8], 1'b0, INIT[ 851*8 +: 8], 1'b0, INIT[ 850*8 +: 8], 
          1'b0, INIT[ 847*8 +: 8], 1'b0, INIT[ 846*8 +: 8], 1'b0, INIT[ 843*8 +: 8], 1'b0, INIT[ 842*8 +: 8], 
          1'b0, INIT[ 839*8 +: 8], 1'b0, INIT[ 838*8 +: 8], 1'b0, INIT[ 835*8 +: 8], 1'b0, INIT[ 834*8 +: 8], 
          1'b0, INIT[ 831*8 +: 8], 1'b0, INIT[ 830*8 +: 8], 1'b0, INIT[ 827*8 +: 8], 1'b0, INIT[ 826*8 +: 8], 
          1'b0, INIT[ 823*8 +: 8], 1'b0, INIT[ 822*8 +: 8], 1'b0, INIT[ 819*8 +: 8], 1'b0, INIT[ 818*8 +: 8], 
          1'b0, INIT[ 815*8 +: 8], 1'b0, INIT[ 814*8 +: 8], 1'b0, INIT[ 811*8 +: 8], 1'b0, INIT[ 810*8 +: 8], 
          1'b0, INIT[ 807*8 +: 8], 1'b0, INIT[ 806*8 +: 8], 1'b0, INIT[ 803*8 +: 8], 1'b0, INIT[ 802*8 +: 8], 
          1'b0, INIT[ 799*8 +: 8], 1'b0, INIT[ 798*8 +: 8], 1'b0, INIT[ 795*8 +: 8], 1'b0, INIT[ 794*8 +: 8], 
          1'b0, INIT[ 791*8 +: 8], 1'b0, INIT[ 790*8 +: 8], 1'b0, INIT[ 787*8 +: 8], 1'b0, INIT[ 786*8 +: 8], 
          1'b0, INIT[ 783*8 +: 8], 1'b0, INIT[ 782*8 +: 8], 1'b0, INIT[ 779*8 +: 8], 1'b0, INIT[ 778*8 +: 8], 
          1'b0, INIT[ 775*8 +: 8], 1'b0, INIT[ 774*8 +: 8], 1'b0, INIT[ 771*8 +: 8], 1'b0, INIT[ 770*8 +: 8], 
          1'b0, INIT[ 767*8 +: 8], 1'b0, INIT[ 766*8 +: 8], 1'b0, INIT[ 763*8 +: 8], 1'b0, INIT[ 762*8 +: 8], 
          1'b0, INIT[ 759*8 +: 8], 1'b0, INIT[ 758*8 +: 8], 1'b0, INIT[ 755*8 +: 8], 1'b0, INIT[ 754*8 +: 8], 
          1'b0, INIT[ 751*8 +: 8], 1'b0, INIT[ 750*8 +: 8], 1'b0, INIT[ 747*8 +: 8], 1'b0, INIT[ 746*8 +: 8], 
          1'b0, INIT[ 743*8 +: 8], 1'b0, INIT[ 742*8 +: 8], 1'b0, INIT[ 739*8 +: 8], 1'b0, INIT[ 738*8 +: 8], 
          1'b0, INIT[ 735*8 +: 8], 1'b0, INIT[ 734*8 +: 8], 1'b0, INIT[ 731*8 +: 8], 1'b0, INIT[ 730*8 +: 8], 
          1'b0, INIT[ 727*8 +: 8], 1'b0, INIT[ 726*8 +: 8], 1'b0, INIT[ 723*8 +: 8], 1'b0, INIT[ 722*8 +: 8], 
          1'b0, INIT[ 719*8 +: 8], 1'b0, INIT[ 718*8 +: 8], 1'b0, INIT[ 715*8 +: 8], 1'b0, INIT[ 714*8 +: 8], 
          1'b0, INIT[ 711*8 +: 8], 1'b0, INIT[ 710*8 +: 8], 1'b0, INIT[ 707*8 +: 8], 1'b0, INIT[ 706*8 +: 8], 
          1'b0, INIT[ 703*8 +: 8], 1'b0, INIT[ 702*8 +: 8], 1'b0, INIT[ 699*8 +: 8], 1'b0, INIT[ 698*8 +: 8], 
          1'b0, INIT[ 695*8 +: 8], 1'b0, INIT[ 694*8 +: 8], 1'b0, INIT[ 691*8 +: 8], 1'b0, INIT[ 690*8 +: 8], 
          1'b0, INIT[ 687*8 +: 8], 1'b0, INIT[ 686*8 +: 8], 1'b0, INIT[ 683*8 +: 8], 1'b0, INIT[ 682*8 +: 8], 
          1'b0, INIT[ 679*8 +: 8], 1'b0, INIT[ 678*8 +: 8], 1'b0, INIT[ 675*8 +: 8], 1'b0, INIT[ 674*8 +: 8], 
          1'b0, INIT[ 671*8 +: 8], 1'b0, INIT[ 670*8 +: 8], 1'b0, INIT[ 667*8 +: 8], 1'b0, INIT[ 666*8 +: 8], 
          1'b0, INIT[ 663*8 +: 8], 1'b0, INIT[ 662*8 +: 8], 1'b0, INIT[ 659*8 +: 8], 1'b0, INIT[ 658*8 +: 8], 
          1'b0, INIT[ 655*8 +: 8], 1'b0, INIT[ 654*8 +: 8], 1'b0, INIT[ 651*8 +: 8], 1'b0, INIT[ 650*8 +: 8], 
          1'b0, INIT[ 647*8 +: 8], 1'b0, INIT[ 646*8 +: 8], 1'b0, INIT[ 643*8 +: 8], 1'b0, INIT[ 642*8 +: 8], 
          1'b0, INIT[ 639*8 +: 8], 1'b0, INIT[ 638*8 +: 8], 1'b0, INIT[ 635*8 +: 8], 1'b0, INIT[ 634*8 +: 8], 
          1'b0, INIT[ 631*8 +: 8], 1'b0, INIT[ 630*8 +: 8], 1'b0, INIT[ 627*8 +: 8], 1'b0, INIT[ 626*8 +: 8], 
          1'b0, INIT[ 623*8 +: 8], 1'b0, INIT[ 622*8 +: 8], 1'b0, INIT[ 619*8 +: 8], 1'b0, INIT[ 618*8 +: 8], 
          1'b0, INIT[ 615*8 +: 8], 1'b0, INIT[ 614*8 +: 8], 1'b0, INIT[ 611*8 +: 8], 1'b0, INIT[ 610*8 +: 8], 
          1'b0, INIT[ 607*8 +: 8], 1'b0, INIT[ 606*8 +: 8], 1'b0, INIT[ 603*8 +: 8], 1'b0, INIT[ 602*8 +: 8], 
          1'b0, INIT[ 599*8 +: 8], 1'b0, INIT[ 598*8 +: 8], 1'b0, INIT[ 595*8 +: 8], 1'b0, INIT[ 594*8 +: 8], 
          1'b0, INIT[ 591*8 +: 8], 1'b0, INIT[ 590*8 +: 8], 1'b0, INIT[ 587*8 +: 8], 1'b0, INIT[ 586*8 +: 8], 
          1'b0, INIT[ 583*8 +: 8], 1'b0, INIT[ 582*8 +: 8], 1'b0, INIT[ 579*8 +: 8], 1'b0, INIT[ 578*8 +: 8], 
          1'b0, INIT[ 575*8 +: 8], 1'b0, INIT[ 574*8 +: 8], 1'b0, INIT[ 571*8 +: 8], 1'b0, INIT[ 570*8 +: 8], 
          1'b0, INIT[ 567*8 +: 8], 1'b0, INIT[ 566*8 +: 8], 1'b0, INIT[ 563*8 +: 8], 1'b0, INIT[ 562*8 +: 8], 
          1'b0, INIT[ 559*8 +: 8], 1'b0, INIT[ 558*8 +: 8], 1'b0, INIT[ 555*8 +: 8], 1'b0, INIT[ 554*8 +: 8], 
          1'b0, INIT[ 551*8 +: 8], 1'b0, INIT[ 550*8 +: 8], 1'b0, INIT[ 547*8 +: 8], 1'b0, INIT[ 546*8 +: 8], 
          1'b0, INIT[ 543*8 +: 8], 1'b0, INIT[ 542*8 +: 8], 1'b0, INIT[ 539*8 +: 8], 1'b0, INIT[ 538*8 +: 8], 
          1'b0, INIT[ 535*8 +: 8], 1'b0, INIT[ 534*8 +: 8], 1'b0, INIT[ 531*8 +: 8], 1'b0, INIT[ 530*8 +: 8], 
          1'b0, INIT[ 527*8 +: 8], 1'b0, INIT[ 526*8 +: 8], 1'b0, INIT[ 523*8 +: 8], 1'b0, INIT[ 522*8 +: 8], 
          1'b0, INIT[ 519*8 +: 8], 1'b0, INIT[ 518*8 +: 8], 1'b0, INIT[ 515*8 +: 8], 1'b0, INIT[ 514*8 +: 8], 
          1'b0, INIT[ 511*8 +: 8], 1'b0, INIT[ 510*8 +: 8], 1'b0, INIT[ 507*8 +: 8], 1'b0, INIT[ 506*8 +: 8], 
          1'b0, INIT[ 503*8 +: 8], 1'b0, INIT[ 502*8 +: 8], 1'b0, INIT[ 499*8 +: 8], 1'b0, INIT[ 498*8 +: 8], 
          1'b0, INIT[ 495*8 +: 8], 1'b0, INIT[ 494*8 +: 8], 1'b0, INIT[ 491*8 +: 8], 1'b0, INIT[ 490*8 +: 8], 
          1'b0, INIT[ 487*8 +: 8], 1'b0, INIT[ 486*8 +: 8], 1'b0, INIT[ 483*8 +: 8], 1'b0, INIT[ 482*8 +: 8], 
          1'b0, INIT[ 479*8 +: 8], 1'b0, INIT[ 478*8 +: 8], 1'b0, INIT[ 475*8 +: 8], 1'b0, INIT[ 474*8 +: 8], 
          1'b0, INIT[ 471*8 +: 8], 1'b0, INIT[ 470*8 +: 8], 1'b0, INIT[ 467*8 +: 8], 1'b0, INIT[ 466*8 +: 8], 
          1'b0, INIT[ 463*8 +: 8], 1'b0, INIT[ 462*8 +: 8], 1'b0, INIT[ 459*8 +: 8], 1'b0, INIT[ 458*8 +: 8], 
          1'b0, INIT[ 455*8 +: 8], 1'b0, INIT[ 454*8 +: 8], 1'b0, INIT[ 451*8 +: 8], 1'b0, INIT[ 450*8 +: 8], 
          1'b0, INIT[ 447*8 +: 8], 1'b0, INIT[ 446*8 +: 8], 1'b0, INIT[ 443*8 +: 8], 1'b0, INIT[ 442*8 +: 8], 
          1'b0, INIT[ 439*8 +: 8], 1'b0, INIT[ 438*8 +: 8], 1'b0, INIT[ 435*8 +: 8], 1'b0, INIT[ 434*8 +: 8], 
          1'b0, INIT[ 431*8 +: 8], 1'b0, INIT[ 430*8 +: 8], 1'b0, INIT[ 427*8 +: 8], 1'b0, INIT[ 426*8 +: 8], 
          1'b0, INIT[ 423*8 +: 8], 1'b0, INIT[ 422*8 +: 8], 1'b0, INIT[ 419*8 +: 8], 1'b0, INIT[ 418*8 +: 8], 
          1'b0, INIT[ 415*8 +: 8], 1'b0, INIT[ 414*8 +: 8], 1'b0, INIT[ 411*8 +: 8], 1'b0, INIT[ 410*8 +: 8], 
          1'b0, INIT[ 407*8 +: 8], 1'b0, INIT[ 406*8 +: 8], 1'b0, INIT[ 403*8 +: 8], 1'b0, INIT[ 402*8 +: 8], 
          1'b0, INIT[ 399*8 +: 8], 1'b0, INIT[ 398*8 +: 8], 1'b0, INIT[ 395*8 +: 8], 1'b0, INIT[ 394*8 +: 8], 
          1'b0, INIT[ 391*8 +: 8], 1'b0, INIT[ 390*8 +: 8], 1'b0, INIT[ 387*8 +: 8], 1'b0, INIT[ 386*8 +: 8], 
          1'b0, INIT[ 383*8 +: 8], 1'b0, INIT[ 382*8 +: 8], 1'b0, INIT[ 379*8 +: 8], 1'b0, INIT[ 378*8 +: 8], 
          1'b0, INIT[ 375*8 +: 8], 1'b0, INIT[ 374*8 +: 8], 1'b0, INIT[ 371*8 +: 8], 1'b0, INIT[ 370*8 +: 8], 
          1'b0, INIT[ 367*8 +: 8], 1'b0, INIT[ 366*8 +: 8], 1'b0, INIT[ 363*8 +: 8], 1'b0, INIT[ 362*8 +: 8], 
          1'b0, INIT[ 359*8 +: 8], 1'b0, INIT[ 358*8 +: 8], 1'b0, INIT[ 355*8 +: 8], 1'b0, INIT[ 354*8 +: 8], 
          1'b0, INIT[ 351*8 +: 8], 1'b0, INIT[ 350*8 +: 8], 1'b0, INIT[ 347*8 +: 8], 1'b0, INIT[ 346*8 +: 8], 
          1'b0, INIT[ 343*8 +: 8], 1'b0, INIT[ 342*8 +: 8], 1'b0, INIT[ 339*8 +: 8], 1'b0, INIT[ 338*8 +: 8], 
          1'b0, INIT[ 335*8 +: 8], 1'b0, INIT[ 334*8 +: 8], 1'b0, INIT[ 331*8 +: 8], 1'b0, INIT[ 330*8 +: 8], 
          1'b0, INIT[ 327*8 +: 8], 1'b0, INIT[ 326*8 +: 8], 1'b0, INIT[ 323*8 +: 8], 1'b0, INIT[ 322*8 +: 8], 
          1'b0, INIT[ 319*8 +: 8], 1'b0, INIT[ 318*8 +: 8], 1'b0, INIT[ 315*8 +: 8], 1'b0, INIT[ 314*8 +: 8], 
          1'b0, INIT[ 311*8 +: 8], 1'b0, INIT[ 310*8 +: 8], 1'b0, INIT[ 307*8 +: 8], 1'b0, INIT[ 306*8 +: 8], 
          1'b0, INIT[ 303*8 +: 8], 1'b0, INIT[ 302*8 +: 8], 1'b0, INIT[ 299*8 +: 8], 1'b0, INIT[ 298*8 +: 8], 
          1'b0, INIT[ 295*8 +: 8], 1'b0, INIT[ 294*8 +: 8], 1'b0, INIT[ 291*8 +: 8], 1'b0, INIT[ 290*8 +: 8], 
          1'b0, INIT[ 287*8 +: 8], 1'b0, INIT[ 286*8 +: 8], 1'b0, INIT[ 283*8 +: 8], 1'b0, INIT[ 282*8 +: 8], 
          1'b0, INIT[ 279*8 +: 8], 1'b0, INIT[ 278*8 +: 8], 1'b0, INIT[ 275*8 +: 8], 1'b0, INIT[ 274*8 +: 8], 
          1'b0, INIT[ 271*8 +: 8], 1'b0, INIT[ 270*8 +: 8], 1'b0, INIT[ 267*8 +: 8], 1'b0, INIT[ 266*8 +: 8], 
          1'b0, INIT[ 263*8 +: 8], 1'b0, INIT[ 262*8 +: 8], 1'b0, INIT[ 259*8 +: 8], 1'b0, INIT[ 258*8 +: 8], 
          1'b0, INIT[ 255*8 +: 8], 1'b0, INIT[ 254*8 +: 8], 1'b0, INIT[ 251*8 +: 8], 1'b0, INIT[ 250*8 +: 8], 
          1'b0, INIT[ 247*8 +: 8], 1'b0, INIT[ 246*8 +: 8], 1'b0, INIT[ 243*8 +: 8], 1'b0, INIT[ 242*8 +: 8], 
          1'b0, INIT[ 239*8 +: 8], 1'b0, INIT[ 238*8 +: 8], 1'b0, INIT[ 235*8 +: 8], 1'b0, INIT[ 234*8 +: 8], 
          1'b0, INIT[ 231*8 +: 8], 1'b0, INIT[ 230*8 +: 8], 1'b0, INIT[ 227*8 +: 8], 1'b0, INIT[ 226*8 +: 8], 
          1'b0, INIT[ 223*8 +: 8], 1'b0, INIT[ 222*8 +: 8], 1'b0, INIT[ 219*8 +: 8], 1'b0, INIT[ 218*8 +: 8], 
          1'b0, INIT[ 215*8 +: 8], 1'b0, INIT[ 214*8 +: 8], 1'b0, INIT[ 211*8 +: 8], 1'b0, INIT[ 210*8 +: 8], 
          1'b0, INIT[ 207*8 +: 8], 1'b0, INIT[ 206*8 +: 8], 1'b0, INIT[ 203*8 +: 8], 1'b0, INIT[ 202*8 +: 8], 
          1'b0, INIT[ 199*8 +: 8], 1'b0, INIT[ 198*8 +: 8], 1'b0, INIT[ 195*8 +: 8], 1'b0, INIT[ 194*8 +: 8], 
          1'b0, INIT[ 191*8 +: 8], 1'b0, INIT[ 190*8 +: 8], 1'b0, INIT[ 187*8 +: 8], 1'b0, INIT[ 186*8 +: 8], 
          1'b0, INIT[ 183*8 +: 8], 1'b0, INIT[ 182*8 +: 8], 1'b0, INIT[ 179*8 +: 8], 1'b0, INIT[ 178*8 +: 8], 
          1'b0, INIT[ 175*8 +: 8], 1'b0, INIT[ 174*8 +: 8], 1'b0, INIT[ 171*8 +: 8], 1'b0, INIT[ 170*8 +: 8], 
          1'b0, INIT[ 167*8 +: 8], 1'b0, INIT[ 166*8 +: 8], 1'b0, INIT[ 163*8 +: 8], 1'b0, INIT[ 162*8 +: 8], 
          1'b0, INIT[ 159*8 +: 8], 1'b0, INIT[ 158*8 +: 8], 1'b0, INIT[ 155*8 +: 8], 1'b0, INIT[ 154*8 +: 8], 
          1'b0, INIT[ 151*8 +: 8], 1'b0, INIT[ 150*8 +: 8], 1'b0, INIT[ 147*8 +: 8], 1'b0, INIT[ 146*8 +: 8], 
          1'b0, INIT[ 143*8 +: 8], 1'b0, INIT[ 142*8 +: 8], 1'b0, INIT[ 139*8 +: 8], 1'b0, INIT[ 138*8 +: 8], 
          1'b0, INIT[ 135*8 +: 8], 1'b0, INIT[ 134*8 +: 8], 1'b0, INIT[ 131*8 +: 8], 1'b0, INIT[ 130*8 +: 8], 
          1'b0, INIT[ 127*8 +: 8], 1'b0, INIT[ 126*8 +: 8], 1'b0, INIT[ 123*8 +: 8], 1'b0, INIT[ 122*8 +: 8], 
          1'b0, INIT[ 119*8 +: 8], 1'b0, INIT[ 118*8 +: 8], 1'b0, INIT[ 115*8 +: 8], 1'b0, INIT[ 114*8 +: 8], 
          1'b0, INIT[ 111*8 +: 8], 1'b0, INIT[ 110*8 +: 8], 1'b0, INIT[ 107*8 +: 8], 1'b0, INIT[ 106*8 +: 8], 
          1'b0, INIT[ 103*8 +: 8], 1'b0, INIT[ 102*8 +: 8], 1'b0, INIT[  99*8 +: 8], 1'b0, INIT[  98*8 +: 8], 
          1'b0, INIT[  95*8 +: 8], 1'b0, INIT[  94*8 +: 8], 1'b0, INIT[  91*8 +: 8], 1'b0, INIT[  90*8 +: 8], 
          1'b0, INIT[  87*8 +: 8], 1'b0, INIT[  86*8 +: 8], 1'b0, INIT[  83*8 +: 8], 1'b0, INIT[  82*8 +: 8], 
          1'b0, INIT[  79*8 +: 8], 1'b0, INIT[  78*8 +: 8], 1'b0, INIT[  75*8 +: 8], 1'b0, INIT[  74*8 +: 8], 
          1'b0, INIT[  71*8 +: 8], 1'b0, INIT[  70*8 +: 8], 1'b0, INIT[  67*8 +: 8], 1'b0, INIT[  66*8 +: 8], 
          1'b0, INIT[  63*8 +: 8], 1'b0, INIT[  62*8 +: 8], 1'b0, INIT[  59*8 +: 8], 1'b0, INIT[  58*8 +: 8], 
          1'b0, INIT[  55*8 +: 8], 1'b0, INIT[  54*8 +: 8], 1'b0, INIT[  51*8 +: 8], 1'b0, INIT[  50*8 +: 8], 
          1'b0, INIT[  47*8 +: 8], 1'b0, INIT[  46*8 +: 8], 1'b0, INIT[  43*8 +: 8], 1'b0, INIT[  42*8 +: 8], 
          1'b0, INIT[  39*8 +: 8], 1'b0, INIT[  38*8 +: 8], 1'b0, INIT[  35*8 +: 8], 1'b0, INIT[  34*8 +: 8], 
          1'b0, INIT[  31*8 +: 8], 1'b0, INIT[  30*8 +: 8], 1'b0, INIT[  27*8 +: 8], 1'b0, INIT[  26*8 +: 8], 
          1'b0, INIT[  23*8 +: 8], 1'b0, INIT[  22*8 +: 8], 1'b0, INIT[  19*8 +: 8], 1'b0, INIT[  18*8 +: 8], 
          1'b0, INIT[  15*8 +: 8], 1'b0, INIT[  14*8 +: 8], 1'b0, INIT[  11*8 +: 8], 1'b0, INIT[  10*8 +: 8], 
          1'b0, INIT[   7*8 +: 8], 1'b0, INIT[   6*8 +: 8], 1'b0, INIT[   3*8 +: 8], 1'b0, INIT[   2*8 +: 8], 
          1'b0, INIT[2045*8 +: 8], 1'b0, INIT[2044*8 +: 8], 1'b0, INIT[2041*8 +: 8], 1'b0, INIT[2040*8 +: 8], 
          1'b0, INIT[2037*8 +: 8], 1'b0, INIT[2036*8 +: 8], 1'b0, INIT[2033*8 +: 8], 1'b0, INIT[2032*8 +: 8], 
          1'b0, INIT[2029*8 +: 8], 1'b0, INIT[2028*8 +: 8], 1'b0, INIT[2025*8 +: 8], 1'b0, INIT[2024*8 +: 8], 
          1'b0, INIT[2021*8 +: 8], 1'b0, INIT[2020*8 +: 8], 1'b0, INIT[2017*8 +: 8], 1'b0, INIT[2016*8 +: 8], 
          1'b0, INIT[2013*8 +: 8], 1'b0, INIT[2012*8 +: 8], 1'b0, INIT[2009*8 +: 8], 1'b0, INIT[2008*8 +: 8], 
          1'b0, INIT[2005*8 +: 8], 1'b0, INIT[2004*8 +: 8], 1'b0, INIT[2001*8 +: 8], 1'b0, INIT[2000*8 +: 8], 
          1'b0, INIT[1997*8 +: 8], 1'b0, INIT[1996*8 +: 8], 1'b0, INIT[1993*8 +: 8], 1'b0, INIT[1992*8 +: 8], 
          1'b0, INIT[1989*8 +: 8], 1'b0, INIT[1988*8 +: 8], 1'b0, INIT[1985*8 +: 8], 1'b0, INIT[1984*8 +: 8], 
          1'b0, INIT[1981*8 +: 8], 1'b0, INIT[1980*8 +: 8], 1'b0, INIT[1977*8 +: 8], 1'b0, INIT[1976*8 +: 8], 
          1'b0, INIT[1973*8 +: 8], 1'b0, INIT[1972*8 +: 8], 1'b0, INIT[1969*8 +: 8], 1'b0, INIT[1968*8 +: 8], 
          1'b0, INIT[1965*8 +: 8], 1'b0, INIT[1964*8 +: 8], 1'b0, INIT[1961*8 +: 8], 1'b0, INIT[1960*8 +: 8], 
          1'b0, INIT[1957*8 +: 8], 1'b0, INIT[1956*8 +: 8], 1'b0, INIT[1953*8 +: 8], 1'b0, INIT[1952*8 +: 8], 
          1'b0, INIT[1949*8 +: 8], 1'b0, INIT[1948*8 +: 8], 1'b0, INIT[1945*8 +: 8], 1'b0, INIT[1944*8 +: 8], 
          1'b0, INIT[1941*8 +: 8], 1'b0, INIT[1940*8 +: 8], 1'b0, INIT[1937*8 +: 8], 1'b0, INIT[1936*8 +: 8], 
          1'b0, INIT[1933*8 +: 8], 1'b0, INIT[1932*8 +: 8], 1'b0, INIT[1929*8 +: 8], 1'b0, INIT[1928*8 +: 8], 
          1'b0, INIT[1925*8 +: 8], 1'b0, INIT[1924*8 +: 8], 1'b0, INIT[1921*8 +: 8], 1'b0, INIT[1920*8 +: 8], 
          1'b0, INIT[1917*8 +: 8], 1'b0, INIT[1916*8 +: 8], 1'b0, INIT[1913*8 +: 8], 1'b0, INIT[1912*8 +: 8], 
          1'b0, INIT[1909*8 +: 8], 1'b0, INIT[1908*8 +: 8], 1'b0, INIT[1905*8 +: 8], 1'b0, INIT[1904*8 +: 8], 
          1'b0, INIT[1901*8 +: 8], 1'b0, INIT[1900*8 +: 8], 1'b0, INIT[1897*8 +: 8], 1'b0, INIT[1896*8 +: 8], 
          1'b0, INIT[1893*8 +: 8], 1'b0, INIT[1892*8 +: 8], 1'b0, INIT[1889*8 +: 8], 1'b0, INIT[1888*8 +: 8], 
          1'b0, INIT[1885*8 +: 8], 1'b0, INIT[1884*8 +: 8], 1'b0, INIT[1881*8 +: 8], 1'b0, INIT[1880*8 +: 8], 
          1'b0, INIT[1877*8 +: 8], 1'b0, INIT[1876*8 +: 8], 1'b0, INIT[1873*8 +: 8], 1'b0, INIT[1872*8 +: 8], 
          1'b0, INIT[1869*8 +: 8], 1'b0, INIT[1868*8 +: 8], 1'b0, INIT[1865*8 +: 8], 1'b0, INIT[1864*8 +: 8], 
          1'b0, INIT[1861*8 +: 8], 1'b0, INIT[1860*8 +: 8], 1'b0, INIT[1857*8 +: 8], 1'b0, INIT[1856*8 +: 8], 
          1'b0, INIT[1853*8 +: 8], 1'b0, INIT[1852*8 +: 8], 1'b0, INIT[1849*8 +: 8], 1'b0, INIT[1848*8 +: 8], 
          1'b0, INIT[1845*8 +: 8], 1'b0, INIT[1844*8 +: 8], 1'b0, INIT[1841*8 +: 8], 1'b0, INIT[1840*8 +: 8], 
          1'b0, INIT[1837*8 +: 8], 1'b0, INIT[1836*8 +: 8], 1'b0, INIT[1833*8 +: 8], 1'b0, INIT[1832*8 +: 8], 
          1'b0, INIT[1829*8 +: 8], 1'b0, INIT[1828*8 +: 8], 1'b0, INIT[1825*8 +: 8], 1'b0, INIT[1824*8 +: 8], 
          1'b0, INIT[1821*8 +: 8], 1'b0, INIT[1820*8 +: 8], 1'b0, INIT[1817*8 +: 8], 1'b0, INIT[1816*8 +: 8], 
          1'b0, INIT[1813*8 +: 8], 1'b0, INIT[1812*8 +: 8], 1'b0, INIT[1809*8 +: 8], 1'b0, INIT[1808*8 +: 8], 
          1'b0, INIT[1805*8 +: 8], 1'b0, INIT[1804*8 +: 8], 1'b0, INIT[1801*8 +: 8], 1'b0, INIT[1800*8 +: 8], 
          1'b0, INIT[1797*8 +: 8], 1'b0, INIT[1796*8 +: 8], 1'b0, INIT[1793*8 +: 8], 1'b0, INIT[1792*8 +: 8], 
          1'b0, INIT[1789*8 +: 8], 1'b0, INIT[1788*8 +: 8], 1'b0, INIT[1785*8 +: 8], 1'b0, INIT[1784*8 +: 8], 
          1'b0, INIT[1781*8 +: 8], 1'b0, INIT[1780*8 +: 8], 1'b0, INIT[1777*8 +: 8], 1'b0, INIT[1776*8 +: 8], 
          1'b0, INIT[1773*8 +: 8], 1'b0, INIT[1772*8 +: 8], 1'b0, INIT[1769*8 +: 8], 1'b0, INIT[1768*8 +: 8], 
          1'b0, INIT[1765*8 +: 8], 1'b0, INIT[1764*8 +: 8], 1'b0, INIT[1761*8 +: 8], 1'b0, INIT[1760*8 +: 8], 
          1'b0, INIT[1757*8 +: 8], 1'b0, INIT[1756*8 +: 8], 1'b0, INIT[1753*8 +: 8], 1'b0, INIT[1752*8 +: 8], 
          1'b0, INIT[1749*8 +: 8], 1'b0, INIT[1748*8 +: 8], 1'b0, INIT[1745*8 +: 8], 1'b0, INIT[1744*8 +: 8], 
          1'b0, INIT[1741*8 +: 8], 1'b0, INIT[1740*8 +: 8], 1'b0, INIT[1737*8 +: 8], 1'b0, INIT[1736*8 +: 8], 
          1'b0, INIT[1733*8 +: 8], 1'b0, INIT[1732*8 +: 8], 1'b0, INIT[1729*8 +: 8], 1'b0, INIT[1728*8 +: 8], 
          1'b0, INIT[1725*8 +: 8], 1'b0, INIT[1724*8 +: 8], 1'b0, INIT[1721*8 +: 8], 1'b0, INIT[1720*8 +: 8], 
          1'b0, INIT[1717*8 +: 8], 1'b0, INIT[1716*8 +: 8], 1'b0, INIT[1713*8 +: 8], 1'b0, INIT[1712*8 +: 8], 
          1'b0, INIT[1709*8 +: 8], 1'b0, INIT[1708*8 +: 8], 1'b0, INIT[1705*8 +: 8], 1'b0, INIT[1704*8 +: 8], 
          1'b0, INIT[1701*8 +: 8], 1'b0, INIT[1700*8 +: 8], 1'b0, INIT[1697*8 +: 8], 1'b0, INIT[1696*8 +: 8], 
          1'b0, INIT[1693*8 +: 8], 1'b0, INIT[1692*8 +: 8], 1'b0, INIT[1689*8 +: 8], 1'b0, INIT[1688*8 +: 8], 
          1'b0, INIT[1685*8 +: 8], 1'b0, INIT[1684*8 +: 8], 1'b0, INIT[1681*8 +: 8], 1'b0, INIT[1680*8 +: 8], 
          1'b0, INIT[1677*8 +: 8], 1'b0, INIT[1676*8 +: 8], 1'b0, INIT[1673*8 +: 8], 1'b0, INIT[1672*8 +: 8], 
          1'b0, INIT[1669*8 +: 8], 1'b0, INIT[1668*8 +: 8], 1'b0, INIT[1665*8 +: 8], 1'b0, INIT[1664*8 +: 8], 
          1'b0, INIT[1661*8 +: 8], 1'b0, INIT[1660*8 +: 8], 1'b0, INIT[1657*8 +: 8], 1'b0, INIT[1656*8 +: 8], 
          1'b0, INIT[1653*8 +: 8], 1'b0, INIT[1652*8 +: 8], 1'b0, INIT[1649*8 +: 8], 1'b0, INIT[1648*8 +: 8], 
          1'b0, INIT[1645*8 +: 8], 1'b0, INIT[1644*8 +: 8], 1'b0, INIT[1641*8 +: 8], 1'b0, INIT[1640*8 +: 8], 
          1'b0, INIT[1637*8 +: 8], 1'b0, INIT[1636*8 +: 8], 1'b0, INIT[1633*8 +: 8], 1'b0, INIT[1632*8 +: 8], 
          1'b0, INIT[1629*8 +: 8], 1'b0, INIT[1628*8 +: 8], 1'b0, INIT[1625*8 +: 8], 1'b0, INIT[1624*8 +: 8], 
          1'b0, INIT[1621*8 +: 8], 1'b0, INIT[1620*8 +: 8], 1'b0, INIT[1617*8 +: 8], 1'b0, INIT[1616*8 +: 8], 
          1'b0, INIT[1613*8 +: 8], 1'b0, INIT[1612*8 +: 8], 1'b0, INIT[1609*8 +: 8], 1'b0, INIT[1608*8 +: 8], 
          1'b0, INIT[1605*8 +: 8], 1'b0, INIT[1604*8 +: 8], 1'b0, INIT[1601*8 +: 8], 1'b0, INIT[1600*8 +: 8], 
          1'b0, INIT[1597*8 +: 8], 1'b0, INIT[1596*8 +: 8], 1'b0, INIT[1593*8 +: 8], 1'b0, INIT[1592*8 +: 8], 
          1'b0, INIT[1589*8 +: 8], 1'b0, INIT[1588*8 +: 8], 1'b0, INIT[1585*8 +: 8], 1'b0, INIT[1584*8 +: 8], 
          1'b0, INIT[1581*8 +: 8], 1'b0, INIT[1580*8 +: 8], 1'b0, INIT[1577*8 +: 8], 1'b0, INIT[1576*8 +: 8], 
          1'b0, INIT[1573*8 +: 8], 1'b0, INIT[1572*8 +: 8], 1'b0, INIT[1569*8 +: 8], 1'b0, INIT[1568*8 +: 8], 
          1'b0, INIT[1565*8 +: 8], 1'b0, INIT[1564*8 +: 8], 1'b0, INIT[1561*8 +: 8], 1'b0, INIT[1560*8 +: 8], 
          1'b0, INIT[1557*8 +: 8], 1'b0, INIT[1556*8 +: 8], 1'b0, INIT[1553*8 +: 8], 1'b0, INIT[1552*8 +: 8], 
          1'b0, INIT[1549*8 +: 8], 1'b0, INIT[1548*8 +: 8], 1'b0, INIT[1545*8 +: 8], 1'b0, INIT[1544*8 +: 8], 
          1'b0, INIT[1541*8 +: 8], 1'b0, INIT[1540*8 +: 8], 1'b0, INIT[1537*8 +: 8], 1'b0, INIT[1536*8 +: 8], 
          1'b0, INIT[1533*8 +: 8], 1'b0, INIT[1532*8 +: 8], 1'b0, INIT[1529*8 +: 8], 1'b0, INIT[1528*8 +: 8], 
          1'b0, INIT[1525*8 +: 8], 1'b0, INIT[1524*8 +: 8], 1'b0, INIT[1521*8 +: 8], 1'b0, INIT[1520*8 +: 8], 
          1'b0, INIT[1517*8 +: 8], 1'b0, INIT[1516*8 +: 8], 1'b0, INIT[1513*8 +: 8], 1'b0, INIT[1512*8 +: 8], 
          1'b0, INIT[1509*8 +: 8], 1'b0, INIT[1508*8 +: 8], 1'b0, INIT[1505*8 +: 8], 1'b0, INIT[1504*8 +: 8], 
          1'b0, INIT[1501*8 +: 8], 1'b0, INIT[1500*8 +: 8], 1'b0, INIT[1497*8 +: 8], 1'b0, INIT[1496*8 +: 8], 
          1'b0, INIT[1493*8 +: 8], 1'b0, INIT[1492*8 +: 8], 1'b0, INIT[1489*8 +: 8], 1'b0, INIT[1488*8 +: 8], 
          1'b0, INIT[1485*8 +: 8], 1'b0, INIT[1484*8 +: 8], 1'b0, INIT[1481*8 +: 8], 1'b0, INIT[1480*8 +: 8], 
          1'b0, INIT[1477*8 +: 8], 1'b0, INIT[1476*8 +: 8], 1'b0, INIT[1473*8 +: 8], 1'b0, INIT[1472*8 +: 8], 
          1'b0, INIT[1469*8 +: 8], 1'b0, INIT[1468*8 +: 8], 1'b0, INIT[1465*8 +: 8], 1'b0, INIT[1464*8 +: 8], 
          1'b0, INIT[1461*8 +: 8], 1'b0, INIT[1460*8 +: 8], 1'b0, INIT[1457*8 +: 8], 1'b0, INIT[1456*8 +: 8], 
          1'b0, INIT[1453*8 +: 8], 1'b0, INIT[1452*8 +: 8], 1'b0, INIT[1449*8 +: 8], 1'b0, INIT[1448*8 +: 8], 
          1'b0, INIT[1445*8 +: 8], 1'b0, INIT[1444*8 +: 8], 1'b0, INIT[1441*8 +: 8], 1'b0, INIT[1440*8 +: 8], 
          1'b0, INIT[1437*8 +: 8], 1'b0, INIT[1436*8 +: 8], 1'b0, INIT[1433*8 +: 8], 1'b0, INIT[1432*8 +: 8], 
          1'b0, INIT[1429*8 +: 8], 1'b0, INIT[1428*8 +: 8], 1'b0, INIT[1425*8 +: 8], 1'b0, INIT[1424*8 +: 8], 
          1'b0, INIT[1421*8 +: 8], 1'b0, INIT[1420*8 +: 8], 1'b0, INIT[1417*8 +: 8], 1'b0, INIT[1416*8 +: 8], 
          1'b0, INIT[1413*8 +: 8], 1'b0, INIT[1412*8 +: 8], 1'b0, INIT[1409*8 +: 8], 1'b0, INIT[1408*8 +: 8], 
          1'b0, INIT[1405*8 +: 8], 1'b0, INIT[1404*8 +: 8], 1'b0, INIT[1401*8 +: 8], 1'b0, INIT[1400*8 +: 8], 
          1'b0, INIT[1397*8 +: 8], 1'b0, INIT[1396*8 +: 8], 1'b0, INIT[1393*8 +: 8], 1'b0, INIT[1392*8 +: 8], 
          1'b0, INIT[1389*8 +: 8], 1'b0, INIT[1388*8 +: 8], 1'b0, INIT[1385*8 +: 8], 1'b0, INIT[1384*8 +: 8], 
          1'b0, INIT[1381*8 +: 8], 1'b0, INIT[1380*8 +: 8], 1'b0, INIT[1377*8 +: 8], 1'b0, INIT[1376*8 +: 8], 
          1'b0, INIT[1373*8 +: 8], 1'b0, INIT[1372*8 +: 8], 1'b0, INIT[1369*8 +: 8], 1'b0, INIT[1368*8 +: 8], 
          1'b0, INIT[1365*8 +: 8], 1'b0, INIT[1364*8 +: 8], 1'b0, INIT[1361*8 +: 8], 1'b0, INIT[1360*8 +: 8], 
          1'b0, INIT[1357*8 +: 8], 1'b0, INIT[1356*8 +: 8], 1'b0, INIT[1353*8 +: 8], 1'b0, INIT[1352*8 +: 8], 
          1'b0, INIT[1349*8 +: 8], 1'b0, INIT[1348*8 +: 8], 1'b0, INIT[1345*8 +: 8], 1'b0, INIT[1344*8 +: 8], 
          1'b0, INIT[1341*8 +: 8], 1'b0, INIT[1340*8 +: 8], 1'b0, INIT[1337*8 +: 8], 1'b0, INIT[1336*8 +: 8], 
          1'b0, INIT[1333*8 +: 8], 1'b0, INIT[1332*8 +: 8], 1'b0, INIT[1329*8 +: 8], 1'b0, INIT[1328*8 +: 8], 
          1'b0, INIT[1325*8 +: 8], 1'b0, INIT[1324*8 +: 8], 1'b0, INIT[1321*8 +: 8], 1'b0, INIT[1320*8 +: 8], 
          1'b0, INIT[1317*8 +: 8], 1'b0, INIT[1316*8 +: 8], 1'b0, INIT[1313*8 +: 8], 1'b0, INIT[1312*8 +: 8], 
          1'b0, INIT[1309*8 +: 8], 1'b0, INIT[1308*8 +: 8], 1'b0, INIT[1305*8 +: 8], 1'b0, INIT[1304*8 +: 8], 
          1'b0, INIT[1301*8 +: 8], 1'b0, INIT[1300*8 +: 8], 1'b0, INIT[1297*8 +: 8], 1'b0, INIT[1296*8 +: 8], 
          1'b0, INIT[1293*8 +: 8], 1'b0, INIT[1292*8 +: 8], 1'b0, INIT[1289*8 +: 8], 1'b0, INIT[1288*8 +: 8], 
          1'b0, INIT[1285*8 +: 8], 1'b0, INIT[1284*8 +: 8], 1'b0, INIT[1281*8 +: 8], 1'b0, INIT[1280*8 +: 8], 
          1'b0, INIT[1277*8 +: 8], 1'b0, INIT[1276*8 +: 8], 1'b0, INIT[1273*8 +: 8], 1'b0, INIT[1272*8 +: 8], 
          1'b0, INIT[1269*8 +: 8], 1'b0, INIT[1268*8 +: 8], 1'b0, INIT[1265*8 +: 8], 1'b0, INIT[1264*8 +: 8], 
          1'b0, INIT[1261*8 +: 8], 1'b0, INIT[1260*8 +: 8], 1'b0, INIT[1257*8 +: 8], 1'b0, INIT[1256*8 +: 8], 
          1'b0, INIT[1253*8 +: 8], 1'b0, INIT[1252*8 +: 8], 1'b0, INIT[1249*8 +: 8], 1'b0, INIT[1248*8 +: 8], 
          1'b0, INIT[1245*8 +: 8], 1'b0, INIT[1244*8 +: 8], 1'b0, INIT[1241*8 +: 8], 1'b0, INIT[1240*8 +: 8], 
          1'b0, INIT[1237*8 +: 8], 1'b0, INIT[1236*8 +: 8], 1'b0, INIT[1233*8 +: 8], 1'b0, INIT[1232*8 +: 8], 
          1'b0, INIT[1229*8 +: 8], 1'b0, INIT[1228*8 +: 8], 1'b0, INIT[1225*8 +: 8], 1'b0, INIT[1224*8 +: 8], 
          1'b0, INIT[1221*8 +: 8], 1'b0, INIT[1220*8 +: 8], 1'b0, INIT[1217*8 +: 8], 1'b0, INIT[1216*8 +: 8], 
          1'b0, INIT[1213*8 +: 8], 1'b0, INIT[1212*8 +: 8], 1'b0, INIT[1209*8 +: 8], 1'b0, INIT[1208*8 +: 8], 
          1'b0, INIT[1205*8 +: 8], 1'b0, INIT[1204*8 +: 8], 1'b0, INIT[1201*8 +: 8], 1'b0, INIT[1200*8 +: 8], 
          1'b0, INIT[1197*8 +: 8], 1'b0, INIT[1196*8 +: 8], 1'b0, INIT[1193*8 +: 8], 1'b0, INIT[1192*8 +: 8], 
          1'b0, INIT[1189*8 +: 8], 1'b0, INIT[1188*8 +: 8], 1'b0, INIT[1185*8 +: 8], 1'b0, INIT[1184*8 +: 8], 
          1'b0, INIT[1181*8 +: 8], 1'b0, INIT[1180*8 +: 8], 1'b0, INIT[1177*8 +: 8], 1'b0, INIT[1176*8 +: 8], 
          1'b0, INIT[1173*8 +: 8], 1'b0, INIT[1172*8 +: 8], 1'b0, INIT[1169*8 +: 8], 1'b0, INIT[1168*8 +: 8], 
          1'b0, INIT[1165*8 +: 8], 1'b0, INIT[1164*8 +: 8], 1'b0, INIT[1161*8 +: 8], 1'b0, INIT[1160*8 +: 8], 
          1'b0, INIT[1157*8 +: 8], 1'b0, INIT[1156*8 +: 8], 1'b0, INIT[1153*8 +: 8], 1'b0, INIT[1152*8 +: 8], 
          1'b0, INIT[1149*8 +: 8], 1'b0, INIT[1148*8 +: 8], 1'b0, INIT[1145*8 +: 8], 1'b0, INIT[1144*8 +: 8], 
          1'b0, INIT[1141*8 +: 8], 1'b0, INIT[1140*8 +: 8], 1'b0, INIT[1137*8 +: 8], 1'b0, INIT[1136*8 +: 8], 
          1'b0, INIT[1133*8 +: 8], 1'b0, INIT[1132*8 +: 8], 1'b0, INIT[1129*8 +: 8], 1'b0, INIT[1128*8 +: 8], 
          1'b0, INIT[1125*8 +: 8], 1'b0, INIT[1124*8 +: 8], 1'b0, INIT[1121*8 +: 8], 1'b0, INIT[1120*8 +: 8], 
          1'b0, INIT[1117*8 +: 8], 1'b0, INIT[1116*8 +: 8], 1'b0, INIT[1113*8 +: 8], 1'b0, INIT[1112*8 +: 8], 
          1'b0, INIT[1109*8 +: 8], 1'b0, INIT[1108*8 +: 8], 1'b0, INIT[1105*8 +: 8], 1'b0, INIT[1104*8 +: 8], 
          1'b0, INIT[1101*8 +: 8], 1'b0, INIT[1100*8 +: 8], 1'b0, INIT[1097*8 +: 8], 1'b0, INIT[1096*8 +: 8], 
          1'b0, INIT[1093*8 +: 8], 1'b0, INIT[1092*8 +: 8], 1'b0, INIT[1089*8 +: 8], 1'b0, INIT[1088*8 +: 8], 
          1'b0, INIT[1085*8 +: 8], 1'b0, INIT[1084*8 +: 8], 1'b0, INIT[1081*8 +: 8], 1'b0, INIT[1080*8 +: 8], 
          1'b0, INIT[1077*8 +: 8], 1'b0, INIT[1076*8 +: 8], 1'b0, INIT[1073*8 +: 8], 1'b0, INIT[1072*8 +: 8], 
          1'b0, INIT[1069*8 +: 8], 1'b0, INIT[1068*8 +: 8], 1'b0, INIT[1065*8 +: 8], 1'b0, INIT[1064*8 +: 8], 
          1'b0, INIT[1061*8 +: 8], 1'b0, INIT[1060*8 +: 8], 1'b0, INIT[1057*8 +: 8], 1'b0, INIT[1056*8 +: 8], 
          1'b0, INIT[1053*8 +: 8], 1'b0, INIT[1052*8 +: 8], 1'b0, INIT[1049*8 +: 8], 1'b0, INIT[1048*8 +: 8], 
          1'b0, INIT[1045*8 +: 8], 1'b0, INIT[1044*8 +: 8], 1'b0, INIT[1041*8 +: 8], 1'b0, INIT[1040*8 +: 8], 
          1'b0, INIT[1037*8 +: 8], 1'b0, INIT[1036*8 +: 8], 1'b0, INIT[1033*8 +: 8], 1'b0, INIT[1032*8 +: 8], 
          1'b0, INIT[1029*8 +: 8], 1'b0, INIT[1028*8 +: 8], 1'b0, INIT[1025*8 +: 8], 1'b0, INIT[1024*8 +: 8], 
          1'b0, INIT[1021*8 +: 8], 1'b0, INIT[1020*8 +: 8], 1'b0, INIT[1017*8 +: 8], 1'b0, INIT[1016*8 +: 8], 
          1'b0, INIT[1013*8 +: 8], 1'b0, INIT[1012*8 +: 8], 1'b0, INIT[1009*8 +: 8], 1'b0, INIT[1008*8 +: 8], 
          1'b0, INIT[1005*8 +: 8], 1'b0, INIT[1004*8 +: 8], 1'b0, INIT[1001*8 +: 8], 1'b0, INIT[1000*8 +: 8], 
          1'b0, INIT[ 997*8 +: 8], 1'b0, INIT[ 996*8 +: 8], 1'b0, INIT[ 993*8 +: 8], 1'b0, INIT[ 992*8 +: 8], 
          1'b0, INIT[ 989*8 +: 8], 1'b0, INIT[ 988*8 +: 8], 1'b0, INIT[ 985*8 +: 8], 1'b0, INIT[ 984*8 +: 8], 
          1'b0, INIT[ 981*8 +: 8], 1'b0, INIT[ 980*8 +: 8], 1'b0, INIT[ 977*8 +: 8], 1'b0, INIT[ 976*8 +: 8], 
          1'b0, INIT[ 973*8 +: 8], 1'b0, INIT[ 972*8 +: 8], 1'b0, INIT[ 969*8 +: 8], 1'b0, INIT[ 968*8 +: 8], 
          1'b0, INIT[ 965*8 +: 8], 1'b0, INIT[ 964*8 +: 8], 1'b0, INIT[ 961*8 +: 8], 1'b0, INIT[ 960*8 +: 8], 
          1'b0, INIT[ 957*8 +: 8], 1'b0, INIT[ 956*8 +: 8], 1'b0, INIT[ 953*8 +: 8], 1'b0, INIT[ 952*8 +: 8], 
          1'b0, INIT[ 949*8 +: 8], 1'b0, INIT[ 948*8 +: 8], 1'b0, INIT[ 945*8 +: 8], 1'b0, INIT[ 944*8 +: 8], 
          1'b0, INIT[ 941*8 +: 8], 1'b0, INIT[ 940*8 +: 8], 1'b0, INIT[ 937*8 +: 8], 1'b0, INIT[ 936*8 +: 8], 
          1'b0, INIT[ 933*8 +: 8], 1'b0, INIT[ 932*8 +: 8], 1'b0, INIT[ 929*8 +: 8], 1'b0, INIT[ 928*8 +: 8], 
          1'b0, INIT[ 925*8 +: 8], 1'b0, INIT[ 924*8 +: 8], 1'b0, INIT[ 921*8 +: 8], 1'b0, INIT[ 920*8 +: 8], 
          1'b0, INIT[ 917*8 +: 8], 1'b0, INIT[ 916*8 +: 8], 1'b0, INIT[ 913*8 +: 8], 1'b0, INIT[ 912*8 +: 8], 
          1'b0, INIT[ 909*8 +: 8], 1'b0, INIT[ 908*8 +: 8], 1'b0, INIT[ 905*8 +: 8], 1'b0, INIT[ 904*8 +: 8], 
          1'b0, INIT[ 901*8 +: 8], 1'b0, INIT[ 900*8 +: 8], 1'b0, INIT[ 897*8 +: 8], 1'b0, INIT[ 896*8 +: 8], 
          1'b0, INIT[ 893*8 +: 8], 1'b0, INIT[ 892*8 +: 8], 1'b0, INIT[ 889*8 +: 8], 1'b0, INIT[ 888*8 +: 8], 
          1'b0, INIT[ 885*8 +: 8], 1'b0, INIT[ 884*8 +: 8], 1'b0, INIT[ 881*8 +: 8], 1'b0, INIT[ 880*8 +: 8], 
          1'b0, INIT[ 877*8 +: 8], 1'b0, INIT[ 876*8 +: 8], 1'b0, INIT[ 873*8 +: 8], 1'b0, INIT[ 872*8 +: 8], 
          1'b0, INIT[ 869*8 +: 8], 1'b0, INIT[ 868*8 +: 8], 1'b0, INIT[ 865*8 +: 8], 1'b0, INIT[ 864*8 +: 8], 
          1'b0, INIT[ 861*8 +: 8], 1'b0, INIT[ 860*8 +: 8], 1'b0, INIT[ 857*8 +: 8], 1'b0, INIT[ 856*8 +: 8], 
          1'b0, INIT[ 853*8 +: 8], 1'b0, INIT[ 852*8 +: 8], 1'b0, INIT[ 849*8 +: 8], 1'b0, INIT[ 848*8 +: 8], 
          1'b0, INIT[ 845*8 +: 8], 1'b0, INIT[ 844*8 +: 8], 1'b0, INIT[ 841*8 +: 8], 1'b0, INIT[ 840*8 +: 8], 
          1'b0, INIT[ 837*8 +: 8], 1'b0, INIT[ 836*8 +: 8], 1'b0, INIT[ 833*8 +: 8], 1'b0, INIT[ 832*8 +: 8], 
          1'b0, INIT[ 829*8 +: 8], 1'b0, INIT[ 828*8 +: 8], 1'b0, INIT[ 825*8 +: 8], 1'b0, INIT[ 824*8 +: 8], 
          1'b0, INIT[ 821*8 +: 8], 1'b0, INIT[ 820*8 +: 8], 1'b0, INIT[ 817*8 +: 8], 1'b0, INIT[ 816*8 +: 8], 
          1'b0, INIT[ 813*8 +: 8], 1'b0, INIT[ 812*8 +: 8], 1'b0, INIT[ 809*8 +: 8], 1'b0, INIT[ 808*8 +: 8], 
          1'b0, INIT[ 805*8 +: 8], 1'b0, INIT[ 804*8 +: 8], 1'b0, INIT[ 801*8 +: 8], 1'b0, INIT[ 800*8 +: 8], 
          1'b0, INIT[ 797*8 +: 8], 1'b0, INIT[ 796*8 +: 8], 1'b0, INIT[ 793*8 +: 8], 1'b0, INIT[ 792*8 +: 8], 
          1'b0, INIT[ 789*8 +: 8], 1'b0, INIT[ 788*8 +: 8], 1'b0, INIT[ 785*8 +: 8], 1'b0, INIT[ 784*8 +: 8], 
          1'b0, INIT[ 781*8 +: 8], 1'b0, INIT[ 780*8 +: 8], 1'b0, INIT[ 777*8 +: 8], 1'b0, INIT[ 776*8 +: 8], 
          1'b0, INIT[ 773*8 +: 8], 1'b0, INIT[ 772*8 +: 8], 1'b0, INIT[ 769*8 +: 8], 1'b0, INIT[ 768*8 +: 8], 
          1'b0, INIT[ 765*8 +: 8], 1'b0, INIT[ 764*8 +: 8], 1'b0, INIT[ 761*8 +: 8], 1'b0, INIT[ 760*8 +: 8], 
          1'b0, INIT[ 757*8 +: 8], 1'b0, INIT[ 756*8 +: 8], 1'b0, INIT[ 753*8 +: 8], 1'b0, INIT[ 752*8 +: 8], 
          1'b0, INIT[ 749*8 +: 8], 1'b0, INIT[ 748*8 +: 8], 1'b0, INIT[ 745*8 +: 8], 1'b0, INIT[ 744*8 +: 8], 
          1'b0, INIT[ 741*8 +: 8], 1'b0, INIT[ 740*8 +: 8], 1'b0, INIT[ 737*8 +: 8], 1'b0, INIT[ 736*8 +: 8], 
          1'b0, INIT[ 733*8 +: 8], 1'b0, INIT[ 732*8 +: 8], 1'b0, INIT[ 729*8 +: 8], 1'b0, INIT[ 728*8 +: 8], 
          1'b0, INIT[ 725*8 +: 8], 1'b0, INIT[ 724*8 +: 8], 1'b0, INIT[ 721*8 +: 8], 1'b0, INIT[ 720*8 +: 8], 
          1'b0, INIT[ 717*8 +: 8], 1'b0, INIT[ 716*8 +: 8], 1'b0, INIT[ 713*8 +: 8], 1'b0, INIT[ 712*8 +: 8], 
          1'b0, INIT[ 709*8 +: 8], 1'b0, INIT[ 708*8 +: 8], 1'b0, INIT[ 705*8 +: 8], 1'b0, INIT[ 704*8 +: 8], 
          1'b0, INIT[ 701*8 +: 8], 1'b0, INIT[ 700*8 +: 8], 1'b0, INIT[ 697*8 +: 8], 1'b0, INIT[ 696*8 +: 8], 
          1'b0, INIT[ 693*8 +: 8], 1'b0, INIT[ 692*8 +: 8], 1'b0, INIT[ 689*8 +: 8], 1'b0, INIT[ 688*8 +: 8], 
          1'b0, INIT[ 685*8 +: 8], 1'b0, INIT[ 684*8 +: 8], 1'b0, INIT[ 681*8 +: 8], 1'b0, INIT[ 680*8 +: 8], 
          1'b0, INIT[ 677*8 +: 8], 1'b0, INIT[ 676*8 +: 8], 1'b0, INIT[ 673*8 +: 8], 1'b0, INIT[ 672*8 +: 8], 
          1'b0, INIT[ 669*8 +: 8], 1'b0, INIT[ 668*8 +: 8], 1'b0, INIT[ 665*8 +: 8], 1'b0, INIT[ 664*8 +: 8], 
          1'b0, INIT[ 661*8 +: 8], 1'b0, INIT[ 660*8 +: 8], 1'b0, INIT[ 657*8 +: 8], 1'b0, INIT[ 656*8 +: 8], 
          1'b0, INIT[ 653*8 +: 8], 1'b0, INIT[ 652*8 +: 8], 1'b0, INIT[ 649*8 +: 8], 1'b0, INIT[ 648*8 +: 8], 
          1'b0, INIT[ 645*8 +: 8], 1'b0, INIT[ 644*8 +: 8], 1'b0, INIT[ 641*8 +: 8], 1'b0, INIT[ 640*8 +: 8], 
          1'b0, INIT[ 637*8 +: 8], 1'b0, INIT[ 636*8 +: 8], 1'b0, INIT[ 633*8 +: 8], 1'b0, INIT[ 632*8 +: 8], 
          1'b0, INIT[ 629*8 +: 8], 1'b0, INIT[ 628*8 +: 8], 1'b0, INIT[ 625*8 +: 8], 1'b0, INIT[ 624*8 +: 8], 
          1'b0, INIT[ 621*8 +: 8], 1'b0, INIT[ 620*8 +: 8], 1'b0, INIT[ 617*8 +: 8], 1'b0, INIT[ 616*8 +: 8], 
          1'b0, INIT[ 613*8 +: 8], 1'b0, INIT[ 612*8 +: 8], 1'b0, INIT[ 609*8 +: 8], 1'b0, INIT[ 608*8 +: 8], 
          1'b0, INIT[ 605*8 +: 8], 1'b0, INIT[ 604*8 +: 8], 1'b0, INIT[ 601*8 +: 8], 1'b0, INIT[ 600*8 +: 8], 
          1'b0, INIT[ 597*8 +: 8], 1'b0, INIT[ 596*8 +: 8], 1'b0, INIT[ 593*8 +: 8], 1'b0, INIT[ 592*8 +: 8], 
          1'b0, INIT[ 589*8 +: 8], 1'b0, INIT[ 588*8 +: 8], 1'b0, INIT[ 585*8 +: 8], 1'b0, INIT[ 584*8 +: 8], 
          1'b0, INIT[ 581*8 +: 8], 1'b0, INIT[ 580*8 +: 8], 1'b0, INIT[ 577*8 +: 8], 1'b0, INIT[ 576*8 +: 8], 
          1'b0, INIT[ 573*8 +: 8], 1'b0, INIT[ 572*8 +: 8], 1'b0, INIT[ 569*8 +: 8], 1'b0, INIT[ 568*8 +: 8], 
          1'b0, INIT[ 565*8 +: 8], 1'b0, INIT[ 564*8 +: 8], 1'b0, INIT[ 561*8 +: 8], 1'b0, INIT[ 560*8 +: 8], 
          1'b0, INIT[ 557*8 +: 8], 1'b0, INIT[ 556*8 +: 8], 1'b0, INIT[ 553*8 +: 8], 1'b0, INIT[ 552*8 +: 8], 
          1'b0, INIT[ 549*8 +: 8], 1'b0, INIT[ 548*8 +: 8], 1'b0, INIT[ 545*8 +: 8], 1'b0, INIT[ 544*8 +: 8], 
          1'b0, INIT[ 541*8 +: 8], 1'b0, INIT[ 540*8 +: 8], 1'b0, INIT[ 537*8 +: 8], 1'b0, INIT[ 536*8 +: 8], 
          1'b0, INIT[ 533*8 +: 8], 1'b0, INIT[ 532*8 +: 8], 1'b0, INIT[ 529*8 +: 8], 1'b0, INIT[ 528*8 +: 8], 
          1'b0, INIT[ 525*8 +: 8], 1'b0, INIT[ 524*8 +: 8], 1'b0, INIT[ 521*8 +: 8], 1'b0, INIT[ 520*8 +: 8], 
          1'b0, INIT[ 517*8 +: 8], 1'b0, INIT[ 516*8 +: 8], 1'b0, INIT[ 513*8 +: 8], 1'b0, INIT[ 512*8 +: 8], 
          1'b0, INIT[ 509*8 +: 8], 1'b0, INIT[ 508*8 +: 8], 1'b0, INIT[ 505*8 +: 8], 1'b0, INIT[ 504*8 +: 8], 
          1'b0, INIT[ 501*8 +: 8], 1'b0, INIT[ 500*8 +: 8], 1'b0, INIT[ 497*8 +: 8], 1'b0, INIT[ 496*8 +: 8], 
          1'b0, INIT[ 493*8 +: 8], 1'b0, INIT[ 492*8 +: 8], 1'b0, INIT[ 489*8 +: 8], 1'b0, INIT[ 488*8 +: 8], 
          1'b0, INIT[ 485*8 +: 8], 1'b0, INIT[ 484*8 +: 8], 1'b0, INIT[ 481*8 +: 8], 1'b0, INIT[ 480*8 +: 8], 
          1'b0, INIT[ 477*8 +: 8], 1'b0, INIT[ 476*8 +: 8], 1'b0, INIT[ 473*8 +: 8], 1'b0, INIT[ 472*8 +: 8], 
          1'b0, INIT[ 469*8 +: 8], 1'b0, INIT[ 468*8 +: 8], 1'b0, INIT[ 465*8 +: 8], 1'b0, INIT[ 464*8 +: 8], 
          1'b0, INIT[ 461*8 +: 8], 1'b0, INIT[ 460*8 +: 8], 1'b0, INIT[ 457*8 +: 8], 1'b0, INIT[ 456*8 +: 8], 
          1'b0, INIT[ 453*8 +: 8], 1'b0, INIT[ 452*8 +: 8], 1'b0, INIT[ 449*8 +: 8], 1'b0, INIT[ 448*8 +: 8], 
          1'b0, INIT[ 445*8 +: 8], 1'b0, INIT[ 444*8 +: 8], 1'b0, INIT[ 441*8 +: 8], 1'b0, INIT[ 440*8 +: 8], 
          1'b0, INIT[ 437*8 +: 8], 1'b0, INIT[ 436*8 +: 8], 1'b0, INIT[ 433*8 +: 8], 1'b0, INIT[ 432*8 +: 8], 
          1'b0, INIT[ 429*8 +: 8], 1'b0, INIT[ 428*8 +: 8], 1'b0, INIT[ 425*8 +: 8], 1'b0, INIT[ 424*8 +: 8], 
          1'b0, INIT[ 421*8 +: 8], 1'b0, INIT[ 420*8 +: 8], 1'b0, INIT[ 417*8 +: 8], 1'b0, INIT[ 416*8 +: 8], 
          1'b0, INIT[ 413*8 +: 8], 1'b0, INIT[ 412*8 +: 8], 1'b0, INIT[ 409*8 +: 8], 1'b0, INIT[ 408*8 +: 8], 
          1'b0, INIT[ 405*8 +: 8], 1'b0, INIT[ 404*8 +: 8], 1'b0, INIT[ 401*8 +: 8], 1'b0, INIT[ 400*8 +: 8], 
          1'b0, INIT[ 397*8 +: 8], 1'b0, INIT[ 396*8 +: 8], 1'b0, INIT[ 393*8 +: 8], 1'b0, INIT[ 392*8 +: 8], 
          1'b0, INIT[ 389*8 +: 8], 1'b0, INIT[ 388*8 +: 8], 1'b0, INIT[ 385*8 +: 8], 1'b0, INIT[ 384*8 +: 8], 
          1'b0, INIT[ 381*8 +: 8], 1'b0, INIT[ 380*8 +: 8], 1'b0, INIT[ 377*8 +: 8], 1'b0, INIT[ 376*8 +: 8], 
          1'b0, INIT[ 373*8 +: 8], 1'b0, INIT[ 372*8 +: 8], 1'b0, INIT[ 369*8 +: 8], 1'b0, INIT[ 368*8 +: 8], 
          1'b0, INIT[ 365*8 +: 8], 1'b0, INIT[ 364*8 +: 8], 1'b0, INIT[ 361*8 +: 8], 1'b0, INIT[ 360*8 +: 8], 
          1'b0, INIT[ 357*8 +: 8], 1'b0, INIT[ 356*8 +: 8], 1'b0, INIT[ 353*8 +: 8], 1'b0, INIT[ 352*8 +: 8], 
          1'b0, INIT[ 349*8 +: 8], 1'b0, INIT[ 348*8 +: 8], 1'b0, INIT[ 345*8 +: 8], 1'b0, INIT[ 344*8 +: 8], 
          1'b0, INIT[ 341*8 +: 8], 1'b0, INIT[ 340*8 +: 8], 1'b0, INIT[ 337*8 +: 8], 1'b0, INIT[ 336*8 +: 8], 
          1'b0, INIT[ 333*8 +: 8], 1'b0, INIT[ 332*8 +: 8], 1'b0, INIT[ 329*8 +: 8], 1'b0, INIT[ 328*8 +: 8], 
          1'b0, INIT[ 325*8 +: 8], 1'b0, INIT[ 324*8 +: 8], 1'b0, INIT[ 321*8 +: 8], 1'b0, INIT[ 320*8 +: 8], 
          1'b0, INIT[ 317*8 +: 8], 1'b0, INIT[ 316*8 +: 8], 1'b0, INIT[ 313*8 +: 8], 1'b0, INIT[ 312*8 +: 8], 
          1'b0, INIT[ 309*8 +: 8], 1'b0, INIT[ 308*8 +: 8], 1'b0, INIT[ 305*8 +: 8], 1'b0, INIT[ 304*8 +: 8], 
          1'b0, INIT[ 301*8 +: 8], 1'b0, INIT[ 300*8 +: 8], 1'b0, INIT[ 297*8 +: 8], 1'b0, INIT[ 296*8 +: 8], 
          1'b0, INIT[ 293*8 +: 8], 1'b0, INIT[ 292*8 +: 8], 1'b0, INIT[ 289*8 +: 8], 1'b0, INIT[ 288*8 +: 8], 
          1'b0, INIT[ 285*8 +: 8], 1'b0, INIT[ 284*8 +: 8], 1'b0, INIT[ 281*8 +: 8], 1'b0, INIT[ 280*8 +: 8], 
          1'b0, INIT[ 277*8 +: 8], 1'b0, INIT[ 276*8 +: 8], 1'b0, INIT[ 273*8 +: 8], 1'b0, INIT[ 272*8 +: 8], 
          1'b0, INIT[ 269*8 +: 8], 1'b0, INIT[ 268*8 +: 8], 1'b0, INIT[ 265*8 +: 8], 1'b0, INIT[ 264*8 +: 8], 
          1'b0, INIT[ 261*8 +: 8], 1'b0, INIT[ 260*8 +: 8], 1'b0, INIT[ 257*8 +: 8], 1'b0, INIT[ 256*8 +: 8], 
          1'b0, INIT[ 253*8 +: 8], 1'b0, INIT[ 252*8 +: 8], 1'b0, INIT[ 249*8 +: 8], 1'b0, INIT[ 248*8 +: 8], 
          1'b0, INIT[ 245*8 +: 8], 1'b0, INIT[ 244*8 +: 8], 1'b0, INIT[ 241*8 +: 8], 1'b0, INIT[ 240*8 +: 8], 
          1'b0, INIT[ 237*8 +: 8], 1'b0, INIT[ 236*8 +: 8], 1'b0, INIT[ 233*8 +: 8], 1'b0, INIT[ 232*8 +: 8], 
          1'b0, INIT[ 229*8 +: 8], 1'b0, INIT[ 228*8 +: 8], 1'b0, INIT[ 225*8 +: 8], 1'b0, INIT[ 224*8 +: 8], 
          1'b0, INIT[ 221*8 +: 8], 1'b0, INIT[ 220*8 +: 8], 1'b0, INIT[ 217*8 +: 8], 1'b0, INIT[ 216*8 +: 8], 
          1'b0, INIT[ 213*8 +: 8], 1'b0, INIT[ 212*8 +: 8], 1'b0, INIT[ 209*8 +: 8], 1'b0, INIT[ 208*8 +: 8], 
          1'b0, INIT[ 205*8 +: 8], 1'b0, INIT[ 204*8 +: 8], 1'b0, INIT[ 201*8 +: 8], 1'b0, INIT[ 200*8 +: 8], 
          1'b0, INIT[ 197*8 +: 8], 1'b0, INIT[ 196*8 +: 8], 1'b0, INIT[ 193*8 +: 8], 1'b0, INIT[ 192*8 +: 8], 
          1'b0, INIT[ 189*8 +: 8], 1'b0, INIT[ 188*8 +: 8], 1'b0, INIT[ 185*8 +: 8], 1'b0, INIT[ 184*8 +: 8], 
          1'b0, INIT[ 181*8 +: 8], 1'b0, INIT[ 180*8 +: 8], 1'b0, INIT[ 177*8 +: 8], 1'b0, INIT[ 176*8 +: 8], 
          1'b0, INIT[ 173*8 +: 8], 1'b0, INIT[ 172*8 +: 8], 1'b0, INIT[ 169*8 +: 8], 1'b0, INIT[ 168*8 +: 8], 
          1'b0, INIT[ 165*8 +: 8], 1'b0, INIT[ 164*8 +: 8], 1'b0, INIT[ 161*8 +: 8], 1'b0, INIT[ 160*8 +: 8], 
          1'b0, INIT[ 157*8 +: 8], 1'b0, INIT[ 156*8 +: 8], 1'b0, INIT[ 153*8 +: 8], 1'b0, INIT[ 152*8 +: 8], 
          1'b0, INIT[ 149*8 +: 8], 1'b0, INIT[ 148*8 +: 8], 1'b0, INIT[ 145*8 +: 8], 1'b0, INIT[ 144*8 +: 8], 
          1'b0, INIT[ 141*8 +: 8], 1'b0, INIT[ 140*8 +: 8], 1'b0, INIT[ 137*8 +: 8], 1'b0, INIT[ 136*8 +: 8], 
          1'b0, INIT[ 133*8 +: 8], 1'b0, INIT[ 132*8 +: 8], 1'b0, INIT[ 129*8 +: 8], 1'b0, INIT[ 128*8 +: 8], 
          1'b0, INIT[ 125*8 +: 8], 1'b0, INIT[ 124*8 +: 8], 1'b0, INIT[ 121*8 +: 8], 1'b0, INIT[ 120*8 +: 8], 
          1'b0, INIT[ 117*8 +: 8], 1'b0, INIT[ 116*8 +: 8], 1'b0, INIT[ 113*8 +: 8], 1'b0, INIT[ 112*8 +: 8], 
          1'b0, INIT[ 109*8 +: 8], 1'b0, INIT[ 108*8 +: 8], 1'b0, INIT[ 105*8 +: 8], 1'b0, INIT[ 104*8 +: 8], 
          1'b0, INIT[ 101*8 +: 8], 1'b0, INIT[ 100*8 +: 8], 1'b0, INIT[  97*8 +: 8], 1'b0, INIT[  96*8 +: 8], 
          1'b0, INIT[  93*8 +: 8], 1'b0, INIT[  92*8 +: 8], 1'b0, INIT[  89*8 +: 8], 1'b0, INIT[  88*8 +: 8], 
          1'b0, INIT[  85*8 +: 8], 1'b0, INIT[  84*8 +: 8], 1'b0, INIT[  81*8 +: 8], 1'b0, INIT[  80*8 +: 8], 
          1'b0, INIT[  77*8 +: 8], 1'b0, INIT[  76*8 +: 8], 1'b0, INIT[  73*8 +: 8], 1'b0, INIT[  72*8 +: 8], 
          1'b0, INIT[  69*8 +: 8], 1'b0, INIT[  68*8 +: 8], 1'b0, INIT[  65*8 +: 8], 1'b0, INIT[  64*8 +: 8], 
          1'b0, INIT[  61*8 +: 8], 1'b0, INIT[  60*8 +: 8], 1'b0, INIT[  57*8 +: 8], 1'b0, INIT[  56*8 +: 8], 
          1'b0, INIT[  53*8 +: 8], 1'b0, INIT[  52*8 +: 8], 1'b0, INIT[  49*8 +: 8], 1'b0, INIT[  48*8 +: 8], 
          1'b0, INIT[  45*8 +: 8], 1'b0, INIT[  44*8 +: 8], 1'b0, INIT[  41*8 +: 8], 1'b0, INIT[  40*8 +: 8], 
          1'b0, INIT[  37*8 +: 8], 1'b0, INIT[  36*8 +: 8], 1'b0, INIT[  33*8 +: 8], 1'b0, INIT[  32*8 +: 8], 
          1'b0, INIT[  29*8 +: 8], 1'b0, INIT[  28*8 +: 8], 1'b0, INIT[  25*8 +: 8], 1'b0, INIT[  24*8 +: 8], 
          1'b0, INIT[  21*8 +: 8], 1'b0, INIT[  20*8 +: 8], 1'b0, INIT[  17*8 +: 8], 1'b0, INIT[  16*8 +: 8], 
          1'b0, INIT[  13*8 +: 8], 1'b0, INIT[  12*8 +: 8], 1'b0, INIT[   9*8 +: 8], 1'b0, INIT[   8*8 +: 8], 
          1'b0, INIT[  11*8 +: 8], 1'b0, INIT[   4*8 +: 8], 1'b0, INIT[   1*8 +: 8], 1'b0, INIT[   5*8 +: 8]
          })