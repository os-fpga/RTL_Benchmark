//------------------------------------------------------------------------
// Filename     : atcapbbrg100_config.vh
// Description  : specify APB bridge configurations
//------------------------------------------------------------------------
`ifdef ATCAPBBRG100_CONFIG
`else
`define ATCAPBBRG100_CONFIG

`define ATCAPBBRG100_FLOP_OUT

// Specify APB slave according to SoC configuration
`include "ae350_config.vh"
`include "ae350_const.vh"

`define ATCAPBBRG100_SLV_1

`ifdef AE350_UART1_SUPPORT
`define ATCAPBBRG100_SLV_2
`endif

`ifdef AE350_UART2_SUPPORT
`define ATCAPBBRG100_SLV_3
`endif

`ifdef AE350_PIT_SUPPORT
`define ATCAPBBRG100_SLV_4
`endif

`ifdef AE350_WDT_SUPPORT
`define ATCAPBBRG100_SLV_5
`endif

`ifdef AE350_RTC_SUPPORT
`define ATCAPBBRG100_SLV_6
`endif

`ifdef AE350_GPIO_SUPPORT
`define ATCAPBBRG100_SLV_7
`endif

`ifdef AE350_I2C_SUPPORT
`define ATCAPBBRG100_SLV_8
`endif

`ifdef AE350_SPI1_SUPPORT
`define ATCAPBBRG100_SLV_9
`endif

`ifdef AE350_SPI2_SUPPORT
`define ATCAPBBRG100_SLV_10
`endif

`ifdef AE350_SDC_SUPPORT
`define ATCAPBBRG100_SLV_11
`endif

`ifdef AE350_DMA_SUPPORT
`define ATCAPBBRG100_SLV_12
`endif

`ifdef AE350_SSP_SUPPORT
`define ATCAPBBRG100_SLV_13
`endif

`ifdef AE350_DTROM_SUPPORT
`define ATCAPBBRG100_SLV_14
`endif

`ifdef NDS_TRACE_TILELINK
`define ATCAPBBRG100_SLV_15
`endif 

`ifdef ATCAPBBRG100_ADDR_WIDTH_24
// NA
`else //~ATCAPBBRG100_ADDR_WIDTH_24
	`define	ATCAPBBRG100_ADDR_DECODE_WIDTH	28
	`define	ATCAPBBRG100_SLV1_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0100000
	`define	ATCAPBBRG100_SLV2_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0200000
	`define	ATCAPBBRG100_SLV3_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0300000
	`define	ATCAPBBRG100_SLV4_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0400000
	`define	ATCAPBBRG100_SLV5_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0500000
	`define	ATCAPBBRG100_SLV6_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0600000
	`define	ATCAPBBRG100_SLV7_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0700000
	`define	ATCAPBBRG100_SLV8_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0A00000
	`define	ATCAPBBRG100_SLV9_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0B00000
	`define	ATCAPBBRG100_SLV10_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0F00000
	`define	ATCAPBBRG100_SLV11_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0e00000
	`define	ATCAPBBRG100_SLV12_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0C00000
	`define	ATCAPBBRG100_SLV13_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0d00000
	`define	ATCAPBBRG100_SLV14_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h2000000	// DTROM
	`define	ATCAPBBRG100_SLV15_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0800000	// Signal Dump

	`define	ATCAPBBRG100_SLV1_SIZE		1
	`define	ATCAPBBRG100_SLV2_SIZE		1
	`define	ATCAPBBRG100_SLV3_SIZE		1
	`define	ATCAPBBRG100_SLV4_SIZE		1
	`define	ATCAPBBRG100_SLV5_SIZE		1
	`define	ATCAPBBRG100_SLV6_SIZE		1
	`define	ATCAPBBRG100_SLV7_SIZE		1
	`define	ATCAPBBRG100_SLV8_SIZE		1
	`define	ATCAPBBRG100_SLV9_SIZE		1
	`define	ATCAPBBRG100_SLV10_SIZE		1
	`define	ATCAPBBRG100_SLV11_SIZE		1
	`define	ATCAPBBRG100_SLV12_SIZE		1
	`define	ATCAPBBRG100_SLV13_SIZE		1
	`define	ATCAPBBRG100_SLV14_SIZE		1
	`define	ATCAPBBRG100_SLV15_SIZE		1
`endif //ATCAPBBRG100_ADDR_WIDTH_24

`endif //ATCAPBBRG100_CONFIG
