// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: data_output_monitor.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Sat Apr 27 13:59:59 2019
//=============================================================================
// Description: Monitor for data_output
//=============================================================================

`ifndef DATA_OUTPUT_MONITOR_SV
`define DATA_OUTPUT_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file data_output.tpl

class data_output_monitor extends uvm_monitor;

  `uvm_component_utils(data_output_monitor)

  virtual data_output_if vif;

  uvm_analysis_port #(output_tx) analysis_port;

  output_tx m_trans;

  extern function new(string name, uvm_component parent);

  // Methods build_phase, run_phase, and do_mon generated by setting monitor_inc in file data_output.tpl
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file data_output.tpl

endclass : data_output_monitor 


function data_output_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


function void data_output_monitor::build_phase(uvm_phase phase);
endfunction : build_phase


task data_output_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = output_tx::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/data_output_do_mon.sv
task data_output_monitor::do_mon;
  forever @(posedge vif.clk)
  begin
    wait (vif.reset == 1);
    if (vif.valid && vif.ready)
    begin
      m_trans.data = vif.data;
      analysis_port.write(m_trans);
      `uvm_info(get_type_name(), $sformatf("Output data = %0d",m_trans.data), UVM_HIGH)
    end
  end
endtask
// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file data_output.tpl

`endif // DATA_OUTPUT_MONITOR_SV

