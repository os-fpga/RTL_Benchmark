--
-- crc32_fast1024_tab.vhd: A 32-bit CRC (IEEE) table for processing fixed 1024 bits in parallel
-- Copyright (C) 2011 CESNET
-- Author(s): Lukas Kekely <xkekel00@stud.fit.vutbr.cz>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;
use WORK.math_pack.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity crc32_fast1024_tab is
   port(
      DI    : in  std_logic_vector(1024-1 downto 0);
      DO    : out std_logic_vector(31 downto 0)
   );
end entity crc32_fast1024_tab;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture arch of crc32_fast1024_tab is
begin
-- 32-bit CRC equations processing 1024 bits in parallel (VHDL code)
-- Generator polynomial: 0x104C11DB7
   DO(0) <= DI(576) XOR DI(269) XOR DI(1000) XOR DI(42) XOR DI(748) XOR DI(354) XOR DI(587) XOR DI(769) XOR DI(776) XOR DI(906) XOR DI(86) XOR DI(46) XOR DI(280) XOR DI(868) XOR DI(707) XOR DI(588) XOR DI(446) XOR DI(302) XOR DI(89) XOR DI(380) XOR DI(337) XOR DI(834) XOR DI(995) XOR DI(330) XOR DI(45) XOR DI(797) XOR DI(309) XOR DI(185) XOR DI(855) XOR DI(572) XOR DI(979) XOR DI(559) XOR DI(53) XOR DI(90) XOR DI(940) XOR DI(50) XOR DI(171) XOR DI(91) XOR DI(925) XOR DI(355) XOR DI(689) XOR DI(873) XOR DI(93) XOR DI(575) XOR DI(796) XOR DI(926) XOR DI(838) XOR DI(69) XOR DI(333) XOR DI(417) XOR DI(976) XOR DI(765) XOR DI(734) XOR DI(612) XOR DI(49) XOR DI(106) XOR DI(192) XOR DI(301) XOR DI(841) XOR DI(468) XOR DI(996) XOR DI(858) XOR DI(562) XOR DI(969) XOR DI(966) XOR DI(755) XOR DI(182) XOR DI(831) XOR DI(552) XOR DI(959) XOR DI(956) XOR DI(439) XOR DI(153) XOR DI(638) XOR DI(358) XOR DI(580) XOR DI(704) XOR DI(123) XOR DI(449) XOR DI(163) XOR DI(221) XOR DI(737) XOR DI(605) XOR DI(648) XOR DI(240) XOR DI(495) XOR DI(66) XOR DI(702) XOR DI(633) XOR DI(5) XOR DI(187) XOR DI(910) XOR DI(980) XOR DI(842) XOR DI(107) XOR DI(686) XOR DI(368) XOR DI(482) XOR DI(913) XOR DI(998) XOR DI(421) XOR DI(798) XOR DI(531) XOR DI(384) XOR DI(174) XOR DI(927) XOR DI(498) XOR DI(590) XOR DI(800) XOR DI(261) XOR DI(226) XOR DI(636) XOR DI(304) XOR DI(8) XOR DI(977) XOR DI(714) XOR DI(266) XOR DI(104) XOR DI(544) XOR DI(941) XOR DI(356) XOR DI(189) XOR DI(929) XOR DI(133) XOR DI(675) XOR DI(1014) XOR DI(760) XOR DI(767) XOR DI(897) XOR DI(437) XOR DI(371) XOR DI(300) XOR DI(563) XOR DI(787) XOR DI(756) XOR DI(725) XOR DI(292) XOR DI(459) XOR DI(173) XOR DI(822) XOR DI(543) XOR DI(231) XOR DI(57) XOR DI(624) XOR DI(833) XOR DI(359) XOR DI(522) XOR DI(375) XOR DI(918) XOR DI(217) XOR DI(705) XOR DI(257) XOR DI(124) XOR DI(666) XOR DI(751) XOR DI(888) XOR DI(428) XOR DI(747) XOR DI(283) XOR DI(450) XOR DI(534) XOR DI(222) XOR DI(615) XOR DI(513) XOR DI(248) XOR DI(738) XOR DI(441) XOR DI(213) XOR DI(239) XOR DI(729) XOR DI(880) XOR DI(485) XOR DI(814) XOR DI(889) XOR DI(727) XOR DI(404) XOR DI(634) XOR DI(887) XOR DI(658) XOR DI(16) XOR DI(250) XOR DI(608) XOR DI(326) XOR DI(420) XOR DI(505) XOR DI(466) XOR DI(494) XOR DI(71) XOR DI(853) XOR DI(322) XOR DI(30) XOR DI(156) XOR DI(76) XOR DI(911) XOR DI(823) XOR DI(961) XOR DI(547) XOR DI(424) XOR DI(138) XOR DI(148) XOR DI(687) XOR DI(898) XOR DI(999) XOR DI(772) XOR DI(109) XOR DI(736) XOR DI(413) XOR DI(224) XOR DI(470) XOR DI(712) XOR DI(643) XOR DI(15) XOR DI(896) XOR DI(175) XOR DI(928) XOR DI(667) XOR DI(25) XOR DI(259) XOR DI(288) XOR DI(32) XOR DI(591) XOR DI(617) XOR DI(400) XOR DI(335) XOR DI(812) XOR DI(429) XOR DI(866) XOR DI(305) XOR DI(284) XOR DI(545) XOR DI(662) XOR DI(942) XOR DI(126) XOR DI(357) XOR DI(146) XOR DI(190) XOR DI(197) XOR DI(616) XOR DI(943) XOR DI(854) XOR DI(514) XOR DI(533) XOR DI(930) XOR DI(134) XOR DI(475) XOR DI(682) XOR DI(503) XOR DI(1015) XOR DI(994) XOR DI(763) XOR DI(80) XOR DI(40) XOR DI(274) XOR DI(862) XOR DI(83) XOR DI(331) XOR DI(324) XOR DI(39) XOR DI(303) XOR DI(566) XOR DI(47) XOR DI(44) XOR DI(165) XOR DI(85) XOR DI(349) XOR DI(683) XOR DI(790) XOR DI(920) XOR DI(832) XOR DI(411) XOR DI(970) XOR DI(759) XOR DI(728) XOR DI(606) XOR DI(43) XOR DI(295) XOR DI(990) XOR DI(852) XOR DI(556) XOR DI(963) XOR DI(176) XOR DI(825) XOR DI(433) XOR DI(147) XOR DI(632) XOR DI(352) XOR DI(574) XOR DI(117) XOR DI(157) XOR DI(215) XOR DI(489) XOR DI(696) XOR DI(974) XOR DI(836) XOR DI(680) XOR DI(907) XOR DI(992) XOR DI(415) XOR DI(378) XOR DI(921) XOR DI(492) XOR DI(794) XOR DI(255) XOR DI(220) XOR DI(971) XOR DI(538) XOR DI(350) XOR DI(923) XOR DI(127) XOR DI(1008) XOR DI(431) XOR DI(781) XOR DI(750) XOR DI(719) XOR DI(453) XOR DI(167) XOR DI(816) XOR DI(827) XOR DI(516) XOR DI(369) XOR DI(211) XOR DI(118) XOR DI(745) XOR DI(422) XOR DI(741) XOR DI(277) XOR DI(444) XOR DI(216) XOR DI(242) XOR DI(732) XOR DI(233) XOR DI(479) XOR DI(808) XOR DI(721) XOR DI(398) XOR DI(628) XOR DI(881) XOR DI(652) XOR DI(244) XOR DI(602) XOR DI(320) XOR DI(414) XOR DI(499) XOR DI(65) XOR DI(316) XOR DI(24) XOR DI(150) XOR DI(70) XOR DI(905) XOR DI(817) XOR DI(541) XOR DI(418) XOR DI(892) XOR DI(993) XOR DI(730) XOR DI(407) XOR DI(218) XOR DI(464) XOR DI(706) XOR DI(637) XOR DI(9) XOR DI(890) XOR DI(661) XOR DI(19) XOR DI(282) XOR DI(26) XOR DI(394) XOR DI(329) XOR DI(299) XOR DI(656) XOR DI(120) XOR DI(351) XOR DI(184) XOR DI(610) XOR DI(937) XOR DI(508) XOR DI(128) XOR DI(469) XOR DI(676) XOR DI(74) XOR DI(34) XOR DI(268) XOR DI(297) XOR DI(560) XOR DI(41) XOR DI(677) XOR DI(914) XOR DI(826) XOR DI(405) XOR DI(964) XOR DI(722) XOR DI(600) XOR DI(957) XOR DI(170) XOR DI(141) XOR DI(626) XOR DI(151) XOR DI(209) XOR DI(690) XOR DI(830) XOR DI(901) XOR DI(409) XOR DI(372) XOR DI(214) XOR DI(532) XOR DI(344) XOR DI(121) XOR DI(425) XOR DI(161) XOR DI(810) XOR DI(821) XOR DI(510) XOR DI(205) XOR DI(271) XOR DI(438) XOR DI(210) XOR DI(236) XOR DI(726) XOR DI(473) XOR DI(715) XOR DI(392) XOR DI(875) XOR DI(646) XOR DI(238) XOR DI(314) XOR DI(493) XOR DI(18) XOR DI(64) XOR DI(899) XOR DI(535) XOR DI(412) XOR DI(987) XOR DI(724) XOR DI(401) XOR DI(212) XOR DI(631) XOR DI(3) XOR DI(655) XOR DI(13) XOR DI(276) XOR DI(20) XOR DI(388) XOR DI(323) XOR DI(293) XOR DI(650) XOR DI(114) XOR DI(178) XOR DI(502) XOR DI(122) XOR DI(463) XOR DI(28) XOR DI(262) XOR DI(554) XOR DI(671) XOR DI(908) XOR DI(958) XOR DI(951) XOR DI(164) XOR DI(135) XOR DI(620) XOR DI(145) XOR DI(366) XOR DI(208) XOR DI(338) XOR DI(155) XOR DI(815) XOR DI(199) XOR DI(432) XOR DI(467) XOR DI(709) XOR DI(869) XOR DI(12) XOR DI(529) XOR DI(395) XOR DI(206) XOR DI(625) XOR DI(382) XOR DI(317) XOR DI(496) XOR DI(457) XOR DI(548) XOR DI(665) XOR DI(952) XOR DI(945) XOR DI(149) XOR DI(461) XOR DI(703) XOR DI(863) XOR DI(6) XOR DI(523) XOR DI(200) XOR DI(619) XOR DI(376) XOR DI(490) XOR DI(451) XOR DI(542) XOR DI(939) XOR DI(143) XOR DI(697) XOR DI(857) XOR DI(0) XOR DI(517) XOR DI(484) XOR DI(536) XOR DI(137) XOR DI(691) XOR DI(530) XOR DI(131) XOR DI(685) XOR DI(524) XOR DI(125) XOR DI(679) XOR DI(518) XOR DI(512) XOR DI(506) XOR DI(1012) XOR DI(1018);
   DO(1) <= DI(577) XOR DI(270) XOR DI(1001) XOR DI(43) XOR DI(749) XOR DI(355) XOR DI(588) XOR DI(770) XOR DI(777) XOR DI(907) XOR DI(87) XOR DI(47) XOR DI(281) XOR DI(869) XOR DI(708) XOR DI(589) XOR DI(447) XOR DI(303) XOR DI(90) XOR DI(381) XOR DI(338) XOR DI(835) XOR DI(996) XOR DI(331) XOR DI(46) XOR DI(798) XOR DI(310) XOR DI(186) XOR DI(856) XOR DI(573) XOR DI(980) XOR DI(560) XOR DI(54) XOR DI(91) XOR DI(941) XOR DI(51) XOR DI(172) XOR DI(92) XOR DI(926) XOR DI(356) XOR DI(690) XOR DI(874) XOR DI(94) XOR DI(576) XOR DI(797) XOR DI(927) XOR DI(839) XOR DI(70) XOR DI(334) XOR DI(418) XOR DI(977) XOR DI(766) XOR DI(735) XOR DI(613) XOR DI(50) XOR DI(107) XOR DI(193) XOR DI(302) XOR DI(842) XOR DI(469) XOR DI(997) XOR DI(859) XOR DI(563) XOR DI(970) XOR DI(967) XOR DI(756) XOR DI(183) XOR DI(832) XOR DI(553) XOR DI(960) XOR DI(957) XOR DI(440) XOR DI(154) XOR DI(639) XOR DI(359) XOR DI(581) XOR DI(705) XOR DI(124) XOR DI(450) XOR DI(164) XOR DI(222) XOR DI(738) XOR DI(606) XOR DI(649) XOR DI(241) XOR DI(496) XOR DI(67) XOR DI(703) XOR DI(634) XOR DI(6) XOR DI(188) XOR DI(911) XOR DI(981) XOR DI(843) XOR DI(108) XOR DI(687) XOR DI(369) XOR DI(483) XOR DI(914) XOR DI(999) XOR DI(422) XOR DI(799) XOR DI(532) XOR DI(385) XOR DI(175) XOR DI(928) XOR DI(499) XOR DI(591) XOR DI(801) XOR DI(262) XOR DI(227) XOR DI(637) XOR DI(305) XOR DI(9) XOR DI(978) XOR DI(715) XOR DI(267) XOR DI(105) XOR DI(545) XOR DI(942) XOR DI(357) XOR DI(190) XOR DI(930) XOR DI(134) XOR DI(676) XOR DI(1015) XOR DI(761) XOR DI(768) XOR DI(898) XOR DI(438) XOR DI(372) XOR DI(301) XOR DI(564) XOR DI(788) XOR DI(757) XOR DI(726) XOR DI(293) XOR DI(460) XOR DI(174) XOR DI(823) XOR DI(544) XOR DI(232) XOR DI(58) XOR DI(625) XOR DI(834) XOR DI(360) XOR DI(523) XOR DI(376) XOR DI(919) XOR DI(218) XOR DI(706) XOR DI(258) XOR DI(125) XOR DI(667) XOR DI(752) XOR DI(889) XOR DI(429) XOR DI(748) XOR DI(284) XOR DI(451) XOR DI(535) XOR DI(223) XOR DI(616) XOR DI(514) XOR DI(249) XOR DI(739) XOR DI(442) XOR DI(214) XOR DI(240) XOR DI(730) XOR DI(881) XOR DI(486) XOR DI(815) XOR DI(890) XOR DI(728) XOR DI(405) XOR DI(635) XOR DI(888) XOR DI(659) XOR DI(17) XOR DI(251) XOR DI(609) XOR DI(327) XOR DI(421) XOR DI(506) XOR DI(467) XOR DI(495) XOR DI(72) XOR DI(854) XOR DI(323) XOR DI(31) XOR DI(157) XOR DI(77) XOR DI(912) XOR DI(824) XOR DI(962) XOR DI(548) XOR DI(425) XOR DI(139) XOR DI(149) XOR DI(688) XOR DI(899) XOR DI(1000) XOR DI(773) XOR DI(110) XOR DI(737) XOR DI(414) XOR DI(225) XOR DI(471) XOR DI(713) XOR DI(644) XOR DI(16) XOR DI(897) XOR DI(176) XOR DI(929) XOR DI(668) XOR DI(26) XOR DI(260) XOR DI(289) XOR DI(33) XOR DI(592) XOR DI(618) XOR DI(401) XOR DI(336) XOR DI(813) XOR DI(430) XOR DI(867) XOR DI(306) XOR DI(285) XOR DI(546) XOR DI(663) XOR DI(943) XOR DI(127) XOR DI(358) XOR DI(147) XOR DI(191) XOR DI(198) XOR DI(617) XOR DI(944) XOR DI(855) XOR DI(515) XOR DI(534) XOR DI(931) XOR DI(135) XOR DI(476) XOR DI(683) XOR DI(504) XOR DI(1016) XOR DI(995) XOR DI(764) XOR DI(81) XOR DI(41) XOR DI(275) XOR DI(863) XOR DI(84) XOR DI(332) XOR DI(325) XOR DI(40) XOR DI(304) XOR DI(567) XOR DI(48) XOR DI(45) XOR DI(166) XOR DI(86) XOR DI(350) XOR DI(684) XOR DI(791) XOR DI(921) XOR DI(833) XOR DI(412) XOR DI(971) XOR DI(760) XOR DI(729) XOR DI(607) XOR DI(44) XOR DI(296) XOR DI(991) XOR DI(853) XOR DI(557) XOR DI(964) XOR DI(177) XOR DI(826) XOR DI(434) XOR DI(148) XOR DI(633) XOR DI(353) XOR DI(575) XOR DI(118) XOR DI(158) XOR DI(216) XOR DI(490) XOR DI(697) XOR DI(0) XOR DI(975) XOR DI(837) XOR DI(681) XOR DI(908) XOR DI(993) XOR DI(416) XOR DI(379) XOR DI(922) XOR DI(493) XOR DI(795) XOR DI(256) XOR DI(221) XOR DI(972) XOR DI(539) XOR DI(351) XOR DI(924) XOR DI(128) XOR DI(1009) XOR DI(432) XOR DI(782) XOR DI(751) XOR DI(720) XOR DI(454) XOR DI(168) XOR DI(817) XOR DI(828) XOR DI(517) XOR DI(370) XOR DI(212) XOR DI(119) XOR DI(746) XOR DI(423) XOR DI(742) XOR DI(278) XOR DI(445) XOR DI(217) XOR DI(243) XOR DI(733) XOR DI(234) XOR DI(480) XOR DI(809) XOR DI(722) XOR DI(399) XOR DI(629) XOR DI(882) XOR DI(653) XOR DI(245) XOR DI(603) XOR DI(321) XOR DI(415) XOR DI(500) XOR DI(66) XOR DI(317) XOR DI(25) XOR DI(151) XOR DI(71) XOR DI(906) XOR DI(818) XOR DI(542) XOR DI(419) XOR DI(893) XOR DI(994) XOR DI(731) XOR DI(408) XOR DI(219) XOR DI(465) XOR DI(707) XOR DI(638) XOR DI(10) XOR DI(891) XOR DI(662) XOR DI(20) XOR DI(283) XOR DI(27) XOR DI(395) XOR DI(330) XOR DI(300) XOR DI(657) XOR DI(121) XOR DI(352) XOR DI(185) XOR DI(611) XOR DI(938) XOR DI(509) XOR DI(129) XOR DI(470) XOR DI(677) XOR DI(75) XOR DI(35) XOR DI(269) XOR DI(298) XOR DI(561) XOR DI(42) XOR DI(678) XOR DI(915) XOR DI(827) XOR DI(406) XOR DI(965) XOR DI(723) XOR DI(601) XOR DI(958) XOR DI(171) XOR DI(142) XOR DI(627) XOR DI(152) XOR DI(210) XOR DI(691) XOR DI(831) XOR DI(902) XOR DI(410) XOR DI(373) XOR DI(215) XOR DI(533) XOR DI(345) XOR DI(122) XOR DI(426) XOR DI(162) XOR DI(811) XOR DI(822) XOR DI(511) XOR DI(206) XOR DI(272) XOR DI(439) XOR DI(211) XOR DI(237) XOR DI(727) XOR DI(474) XOR DI(716) XOR DI(393) XOR DI(876) XOR DI(647) XOR DI(239) XOR DI(315) XOR DI(494) XOR DI(19) XOR DI(65) XOR DI(900) XOR DI(536) XOR DI(413) XOR DI(988) XOR DI(725) XOR DI(402) XOR DI(213) XOR DI(632) XOR DI(4) XOR DI(656) XOR DI(14) XOR DI(277) XOR DI(21) XOR DI(389) XOR DI(324) XOR DI(294) XOR DI(651) XOR DI(115) XOR DI(179) XOR DI(503) XOR DI(123) XOR DI(464) XOR DI(29) XOR DI(263) XOR DI(555) XOR DI(672) XOR DI(909) XOR DI(959) XOR DI(952) XOR DI(165) XOR DI(136) XOR DI(621) XOR DI(146) XOR DI(367) XOR DI(209) XOR DI(339) XOR DI(156) XOR DI(816) XOR DI(200) XOR DI(433) XOR DI(468) XOR DI(710) XOR DI(870) XOR DI(13) XOR DI(530) XOR DI(396) XOR DI(207) XOR DI(626) XOR DI(383) XOR DI(318) XOR DI(497) XOR DI(458) XOR DI(549) XOR DI(666) XOR DI(953) XOR DI(946) XOR DI(150) XOR DI(462) XOR DI(704) XOR DI(864) XOR DI(7) XOR DI(524) XOR DI(201) XOR DI(620) XOR DI(377) XOR DI(491) XOR DI(452) XOR DI(543) XOR DI(940) XOR DI(144) XOR DI(698) XOR DI(858) XOR DI(1) XOR DI(518) XOR DI(485) XOR DI(537) XOR DI(138) XOR DI(692) XOR DI(531) XOR DI(132) XOR DI(686) XOR DI(525) XOR DI(126) XOR DI(680) XOR DI(519) XOR DI(513) XOR DI(507) XOR DI(1013) XOR DI(1019);
   DO(2) <= DI(578) XOR DI(271) XOR DI(1002) XOR DI(44) XOR DI(750) XOR DI(356) XOR DI(589) XOR DI(771) XOR DI(778) XOR DI(908) XOR DI(88) XOR DI(48) XOR DI(282) XOR DI(870) XOR DI(709) XOR DI(590) XOR DI(448) XOR DI(304) XOR DI(91) XOR DI(382) XOR DI(339) XOR DI(836) XOR DI(997) XOR DI(332) XOR DI(47) XOR DI(799) XOR DI(311) XOR DI(187) XOR DI(857) XOR DI(574) XOR DI(981) XOR DI(561) XOR DI(55) XOR DI(92) XOR DI(942) XOR DI(52) XOR DI(173) XOR DI(93) XOR DI(927) XOR DI(357) XOR DI(691) XOR DI(875) XOR DI(95) XOR DI(577) XOR DI(798) XOR DI(928) XOR DI(840) XOR DI(71) XOR DI(335) XOR DI(419) XOR DI(978) XOR DI(767) XOR DI(736) XOR DI(614) XOR DI(51) XOR DI(108) XOR DI(194) XOR DI(303) XOR DI(843) XOR DI(470) XOR DI(998) XOR DI(860) XOR DI(564) XOR DI(971) XOR DI(968) XOR DI(757) XOR DI(184) XOR DI(833) XOR DI(554) XOR DI(961) XOR DI(958) XOR DI(441) XOR DI(155) XOR DI(640) XOR DI(360) XOR DI(582) XOR DI(706) XOR DI(125) XOR DI(451) XOR DI(165) XOR DI(223) XOR DI(739) XOR DI(607) XOR DI(650) XOR DI(242) XOR DI(497) XOR DI(68) XOR DI(704) XOR DI(635) XOR DI(7) XOR DI(189) XOR DI(912) XOR DI(982) XOR DI(844) XOR DI(109) XOR DI(688) XOR DI(370) XOR DI(484) XOR DI(915) XOR DI(1000) XOR DI(423) XOR DI(800) XOR DI(533) XOR DI(386) XOR DI(176) XOR DI(929) XOR DI(500) XOR DI(592) XOR DI(802) XOR DI(263) XOR DI(228) XOR DI(638) XOR DI(306) XOR DI(10) XOR DI(979) XOR DI(716) XOR DI(268) XOR DI(106) XOR DI(546) XOR DI(943) XOR DI(358) XOR DI(191) XOR DI(931) XOR DI(135) XOR DI(677) XOR DI(1016) XOR DI(762) XOR DI(769) XOR DI(899) XOR DI(439) XOR DI(373) XOR DI(302) XOR DI(565) XOR DI(789) XOR DI(758) XOR DI(727) XOR DI(294) XOR DI(461) XOR DI(175) XOR DI(824) XOR DI(545) XOR DI(233) XOR DI(59) XOR DI(626) XOR DI(835) XOR DI(361) XOR DI(524) XOR DI(377) XOR DI(920) XOR DI(219) XOR DI(707) XOR DI(259) XOR DI(126) XOR DI(668) XOR DI(753) XOR DI(890) XOR DI(430) XOR DI(749) XOR DI(285) XOR DI(452) XOR DI(536) XOR DI(224) XOR DI(617) XOR DI(515) XOR DI(250) XOR DI(740) XOR DI(443) XOR DI(215) XOR DI(241) XOR DI(731) XOR DI(882) XOR DI(487) XOR DI(816) XOR DI(891) XOR DI(729) XOR DI(406) XOR DI(636) XOR DI(889) XOR DI(660) XOR DI(18) XOR DI(252) XOR DI(610) XOR DI(328) XOR DI(422) XOR DI(507) XOR DI(468) XOR DI(496) XOR DI(73) XOR DI(855) XOR DI(324) XOR DI(32) XOR DI(158) XOR DI(78) XOR DI(913) XOR DI(825) XOR DI(963) XOR DI(549) XOR DI(426) XOR DI(140) XOR DI(150) XOR DI(689) XOR DI(900) XOR DI(1001) XOR DI(774) XOR DI(111) XOR DI(738) XOR DI(415) XOR DI(226) XOR DI(472) XOR DI(714) XOR DI(645) XOR DI(17) XOR DI(898) XOR DI(177) XOR DI(930) XOR DI(669) XOR DI(27) XOR DI(261) XOR DI(290) XOR DI(34) XOR DI(593) XOR DI(619) XOR DI(402) XOR DI(337) XOR DI(814) XOR DI(431) XOR DI(868) XOR DI(307) XOR DI(286) XOR DI(547) XOR DI(664) XOR DI(944) XOR DI(128) XOR DI(359) XOR DI(148) XOR DI(192) XOR DI(199) XOR DI(618) XOR DI(945) XOR DI(856) XOR DI(516) XOR DI(535) XOR DI(932) XOR DI(136) XOR DI(477) XOR DI(684) XOR DI(505) XOR DI(1017) XOR DI(996) XOR DI(765) XOR DI(82) XOR DI(42) XOR DI(276) XOR DI(864) XOR DI(85) XOR DI(333) XOR DI(326) XOR DI(41) XOR DI(305) XOR DI(568) XOR DI(49) XOR DI(46) XOR DI(167) XOR DI(87) XOR DI(351) XOR DI(685) XOR DI(792) XOR DI(922) XOR DI(834) XOR DI(413) XOR DI(972) XOR DI(761) XOR DI(730) XOR DI(608) XOR DI(45) XOR DI(297) XOR DI(992) XOR DI(854) XOR DI(558) XOR DI(965) XOR DI(178) XOR DI(827) XOR DI(435) XOR DI(149) XOR DI(634) XOR DI(354) XOR DI(576) XOR DI(119) XOR DI(159) XOR DI(217) XOR DI(491) XOR DI(698) XOR DI(1) XOR DI(976) XOR DI(838) XOR DI(682) XOR DI(909) XOR DI(994) XOR DI(417) XOR DI(380) XOR DI(923) XOR DI(494) XOR DI(796) XOR DI(257) XOR DI(222) XOR DI(973) XOR DI(540) XOR DI(352) XOR DI(925) XOR DI(129) XOR DI(1010) XOR DI(433) XOR DI(783) XOR DI(752) XOR DI(721) XOR DI(455) XOR DI(169) XOR DI(818) XOR DI(829) XOR DI(518) XOR DI(371) XOR DI(213) XOR DI(120) XOR DI(747) XOR DI(424) XOR DI(743) XOR DI(279) XOR DI(446) XOR DI(218) XOR DI(244) XOR DI(734) XOR DI(235) XOR DI(481) XOR DI(810) XOR DI(723) XOR DI(400) XOR DI(630) XOR DI(883) XOR DI(654) XOR DI(246) XOR DI(604) XOR DI(322) XOR DI(416) XOR DI(501) XOR DI(67) XOR DI(318) XOR DI(26) XOR DI(152) XOR DI(72) XOR DI(907) XOR DI(819) XOR DI(543) XOR DI(420) XOR DI(894) XOR DI(995) XOR DI(732) XOR DI(409) XOR DI(220) XOR DI(466) XOR DI(708) XOR DI(639) XOR DI(11) XOR DI(892) XOR DI(663) XOR DI(21) XOR DI(284) XOR DI(28) XOR DI(396) XOR DI(331) XOR DI(301) XOR DI(658) XOR DI(122) XOR DI(353) XOR DI(186) XOR DI(612) XOR DI(939) XOR DI(510) XOR DI(130) XOR DI(471) XOR DI(678) XOR DI(76) XOR DI(36) XOR DI(270) XOR DI(299) XOR DI(562) XOR DI(43) XOR DI(679) XOR DI(916) XOR DI(828) XOR DI(407) XOR DI(966) XOR DI(724) XOR DI(602) XOR DI(959) XOR DI(172) XOR DI(143) XOR DI(628) XOR DI(153) XOR DI(211) XOR DI(692) XOR DI(832) XOR DI(903) XOR DI(411) XOR DI(374) XOR DI(216) XOR DI(534) XOR DI(346) XOR DI(123) XOR DI(427) XOR DI(163) XOR DI(812) XOR DI(823) XOR DI(512) XOR DI(207) XOR DI(273) XOR DI(440) XOR DI(212) XOR DI(238) XOR DI(728) XOR DI(475) XOR DI(717) XOR DI(394) XOR DI(877) XOR DI(648) XOR DI(240) XOR DI(316) XOR DI(495) XOR DI(20) XOR DI(66) XOR DI(901) XOR DI(537) XOR DI(414) XOR DI(989) XOR DI(726) XOR DI(403) XOR DI(214) XOR DI(633) XOR DI(5) XOR DI(657) XOR DI(15) XOR DI(278) XOR DI(22) XOR DI(390) XOR DI(325) XOR DI(295) XOR DI(652) XOR DI(116) XOR DI(180) XOR DI(504) XOR DI(124) XOR DI(465) XOR DI(30) XOR DI(264) XOR DI(556) XOR DI(673) XOR DI(910) XOR DI(960) XOR DI(953) XOR DI(166) XOR DI(137) XOR DI(622) XOR DI(147) XOR DI(368) XOR DI(210) XOR DI(340) XOR DI(157) XOR DI(817) XOR DI(201) XOR DI(434) XOR DI(469) XOR DI(711) XOR DI(871) XOR DI(14) XOR DI(531) XOR DI(397) XOR DI(208) XOR DI(627) XOR DI(384) XOR DI(319) XOR DI(498) XOR DI(459) XOR DI(550) XOR DI(667) XOR DI(954) XOR DI(947) XOR DI(151) XOR DI(463) XOR DI(705) XOR DI(865) XOR DI(8) XOR DI(525) XOR DI(202) XOR DI(621) XOR DI(378) XOR DI(492) XOR DI(453) XOR DI(544) XOR DI(941) XOR DI(145) XOR DI(699) XOR DI(859) XOR DI(2) XOR DI(519) XOR DI(486) XOR DI(538) XOR DI(139) XOR DI(693) XOR DI(532) XOR DI(133) XOR DI(687) XOR DI(526) XOR DI(127) XOR DI(681) XOR DI(520) XOR DI(514) XOR DI(508) XOR DI(1014) XOR DI(1020);
   DO(3) <= DI(579) XOR DI(272) XOR DI(1003) XOR DI(45) XOR DI(751) XOR DI(357) XOR DI(590) XOR DI(772) XOR DI(779) XOR DI(909) XOR DI(89) XOR DI(49) XOR DI(283) XOR DI(871) XOR DI(710) XOR DI(591) XOR DI(449) XOR DI(305) XOR DI(92) XOR DI(383) XOR DI(340) XOR DI(837) XOR DI(998) XOR DI(333) XOR DI(48) XOR DI(800) XOR DI(312) XOR DI(188) XOR DI(858) XOR DI(575) XOR DI(982) XOR DI(562) XOR DI(56) XOR DI(93) XOR DI(943) XOR DI(53) XOR DI(174) XOR DI(94) XOR DI(928) XOR DI(358) XOR DI(692) XOR DI(876) XOR DI(96) XOR DI(578) XOR DI(799) XOR DI(929) XOR DI(841) XOR DI(72) XOR DI(336) XOR DI(420) XOR DI(979) XOR DI(768) XOR DI(737) XOR DI(615) XOR DI(52) XOR DI(109) XOR DI(195) XOR DI(304) XOR DI(844) XOR DI(471) XOR DI(999) XOR DI(861) XOR DI(565) XOR DI(972) XOR DI(969) XOR DI(758) XOR DI(185) XOR DI(834) XOR DI(555) XOR DI(962) XOR DI(959) XOR DI(442) XOR DI(156) XOR DI(641) XOR DI(361) XOR DI(583) XOR DI(707) XOR DI(126) XOR DI(452) XOR DI(166) XOR DI(224) XOR DI(740) XOR DI(608) XOR DI(651) XOR DI(243) XOR DI(498) XOR DI(69) XOR DI(705) XOR DI(636) XOR DI(8) XOR DI(190) XOR DI(913) XOR DI(983) XOR DI(845) XOR DI(110) XOR DI(689) XOR DI(371) XOR DI(485) XOR DI(916) XOR DI(1001) XOR DI(424) XOR DI(801) XOR DI(534) XOR DI(387) XOR DI(177) XOR DI(930) XOR DI(501) XOR DI(593) XOR DI(803) XOR DI(264) XOR DI(229) XOR DI(639) XOR DI(307) XOR DI(11) XOR DI(980) XOR DI(717) XOR DI(269) XOR DI(107) XOR DI(547) XOR DI(944) XOR DI(359) XOR DI(192) XOR DI(932) XOR DI(136) XOR DI(678) XOR DI(1017) XOR DI(763) XOR DI(770) XOR DI(900) XOR DI(440) XOR DI(374) XOR DI(303) XOR DI(566) XOR DI(790) XOR DI(759) XOR DI(728) XOR DI(295) XOR DI(462) XOR DI(176) XOR DI(825) XOR DI(546) XOR DI(234) XOR DI(60) XOR DI(627) XOR DI(836) XOR DI(362) XOR DI(525) XOR DI(378) XOR DI(921) XOR DI(220) XOR DI(708) XOR DI(260) XOR DI(127) XOR DI(669) XOR DI(754) XOR DI(891) XOR DI(431) XOR DI(750) XOR DI(286) XOR DI(453) XOR DI(537) XOR DI(225) XOR DI(618) XOR DI(516) XOR DI(251) XOR DI(741) XOR DI(444) XOR DI(216) XOR DI(242) XOR DI(732) XOR DI(883) XOR DI(488) XOR DI(817) XOR DI(892) XOR DI(730) XOR DI(407) XOR DI(637) XOR DI(890) XOR DI(661) XOR DI(19) XOR DI(253) XOR DI(611) XOR DI(329) XOR DI(423) XOR DI(508) XOR DI(469) XOR DI(497) XOR DI(74) XOR DI(856) XOR DI(325) XOR DI(33) XOR DI(159) XOR DI(79) XOR DI(914) XOR DI(826) XOR DI(964) XOR DI(550) XOR DI(427) XOR DI(141) XOR DI(151) XOR DI(690) XOR DI(901) XOR DI(1002) XOR DI(775) XOR DI(112) XOR DI(739) XOR DI(416) XOR DI(227) XOR DI(473) XOR DI(715) XOR DI(646) XOR DI(18) XOR DI(899) XOR DI(178) XOR DI(931) XOR DI(670) XOR DI(28) XOR DI(262) XOR DI(291) XOR DI(35) XOR DI(594) XOR DI(620) XOR DI(403) XOR DI(338) XOR DI(815) XOR DI(432) XOR DI(869) XOR DI(308) XOR DI(287) XOR DI(548) XOR DI(665) XOR DI(945) XOR DI(129) XOR DI(360) XOR DI(149) XOR DI(193) XOR DI(200) XOR DI(619) XOR DI(946) XOR DI(857) XOR DI(517) XOR DI(536) XOR DI(933) XOR DI(137) XOR DI(478) XOR DI(685) XOR DI(506) XOR DI(1018) XOR DI(997) XOR DI(766) XOR DI(83) XOR DI(43) XOR DI(277) XOR DI(865) XOR DI(86) XOR DI(334) XOR DI(327) XOR DI(42) XOR DI(306) XOR DI(569) XOR DI(50) XOR DI(47) XOR DI(168) XOR DI(88) XOR DI(352) XOR DI(686) XOR DI(793) XOR DI(923) XOR DI(835) XOR DI(414) XOR DI(973) XOR DI(762) XOR DI(731) XOR DI(609) XOR DI(46) XOR DI(298) XOR DI(993) XOR DI(855) XOR DI(559) XOR DI(966) XOR DI(179) XOR DI(828) XOR DI(436) XOR DI(150) XOR DI(635) XOR DI(355) XOR DI(577) XOR DI(120) XOR DI(160) XOR DI(218) XOR DI(492) XOR DI(699) XOR DI(2) XOR DI(977) XOR DI(839) XOR DI(683) XOR DI(910) XOR DI(995) XOR DI(418) XOR DI(381) XOR DI(924) XOR DI(495) XOR DI(797) XOR DI(258) XOR DI(223) XOR DI(974) XOR DI(541) XOR DI(353) XOR DI(926) XOR DI(130) XOR DI(1011) XOR DI(434) XOR DI(784) XOR DI(753) XOR DI(722) XOR DI(456) XOR DI(170) XOR DI(819) XOR DI(830) XOR DI(519) XOR DI(372) XOR DI(214) XOR DI(121) XOR DI(748) XOR DI(425) XOR DI(744) XOR DI(280) XOR DI(447) XOR DI(219) XOR DI(245) XOR DI(735) XOR DI(236) XOR DI(482) XOR DI(811) XOR DI(724) XOR DI(401) XOR DI(631) XOR DI(884) XOR DI(655) XOR DI(247) XOR DI(605) XOR DI(323) XOR DI(417) XOR DI(502) XOR DI(68) XOR DI(319) XOR DI(27) XOR DI(153) XOR DI(73) XOR DI(908) XOR DI(820) XOR DI(544) XOR DI(421) XOR DI(895) XOR DI(996) XOR DI(733) XOR DI(410) XOR DI(221) XOR DI(467) XOR DI(709) XOR DI(640) XOR DI(12) XOR DI(893) XOR DI(664) XOR DI(22) XOR DI(285) XOR DI(29) XOR DI(397) XOR DI(332) XOR DI(302) XOR DI(659) XOR DI(123) XOR DI(354) XOR DI(187) XOR DI(613) XOR DI(940) XOR DI(511) XOR DI(131) XOR DI(472) XOR DI(679) XOR DI(77) XOR DI(37) XOR DI(271) XOR DI(300) XOR DI(563) XOR DI(44) XOR DI(680) XOR DI(917) XOR DI(829) XOR DI(408) XOR DI(967) XOR DI(725) XOR DI(603) XOR DI(960) XOR DI(173) XOR DI(144) XOR DI(629) XOR DI(154) XOR DI(212) XOR DI(693) XOR DI(833) XOR DI(904) XOR DI(412) XOR DI(375) XOR DI(217) XOR DI(535) XOR DI(347) XOR DI(124) XOR DI(428) XOR DI(164) XOR DI(813) XOR DI(824) XOR DI(513) XOR DI(208) XOR DI(274) XOR DI(441) XOR DI(213) XOR DI(239) XOR DI(729) XOR DI(476) XOR DI(718) XOR DI(395) XOR DI(878) XOR DI(649) XOR DI(241) XOR DI(317) XOR DI(496) XOR DI(21) XOR DI(67) XOR DI(902) XOR DI(538) XOR DI(415) XOR DI(990) XOR DI(727) XOR DI(404) XOR DI(215) XOR DI(634) XOR DI(6) XOR DI(658) XOR DI(16) XOR DI(279) XOR DI(23) XOR DI(391) XOR DI(326) XOR DI(296) XOR DI(653) XOR DI(117) XOR DI(181) XOR DI(505) XOR DI(125) XOR DI(466) XOR DI(31) XOR DI(265) XOR DI(557) XOR DI(674) XOR DI(911) XOR DI(961) XOR DI(954) XOR DI(167) XOR DI(138) XOR DI(623) XOR DI(148) XOR DI(369) XOR DI(211) XOR DI(341) XOR DI(158) XOR DI(818) XOR DI(202) XOR DI(435) XOR DI(470) XOR DI(712) XOR DI(872) XOR DI(15) XOR DI(532) XOR DI(398) XOR DI(209) XOR DI(628) XOR DI(385) XOR DI(320) XOR DI(499) XOR DI(460) XOR DI(551) XOR DI(668) XOR DI(955) XOR DI(948) XOR DI(152) XOR DI(464) XOR DI(706) XOR DI(866) XOR DI(9) XOR DI(526) XOR DI(203) XOR DI(622) XOR DI(379) XOR DI(493) XOR DI(454) XOR DI(545) XOR DI(942) XOR DI(146) XOR DI(700) XOR DI(860) XOR DI(3) XOR DI(520) XOR DI(487) XOR DI(539) XOR DI(140) XOR DI(694) XOR DI(533) XOR DI(134) XOR DI(688) XOR DI(527) XOR DI(128) XOR DI(682) XOR DI(521) XOR DI(515) XOR DI(509) XOR DI(1015) XOR DI(1021);
   DO(4) <= DI(580) XOR DI(273) XOR DI(1004) XOR DI(46) XOR DI(752) XOR DI(358) XOR DI(591) XOR DI(773) XOR DI(780) XOR DI(910) XOR DI(90) XOR DI(50) XOR DI(284) XOR DI(872) XOR DI(711) XOR DI(592) XOR DI(450) XOR DI(306) XOR DI(93) XOR DI(384) XOR DI(341) XOR DI(838) XOR DI(999) XOR DI(334) XOR DI(49) XOR DI(801) XOR DI(313) XOR DI(189) XOR DI(859) XOR DI(576) XOR DI(983) XOR DI(563) XOR DI(57) XOR DI(94) XOR DI(944) XOR DI(54) XOR DI(175) XOR DI(95) XOR DI(929) XOR DI(359) XOR DI(693) XOR DI(877) XOR DI(97) XOR DI(579) XOR DI(800) XOR DI(930) XOR DI(842) XOR DI(73) XOR DI(337) XOR DI(421) XOR DI(980) XOR DI(769) XOR DI(738) XOR DI(616) XOR DI(53) XOR DI(110) XOR DI(196) XOR DI(305) XOR DI(845) XOR DI(472) XOR DI(1000) XOR DI(862) XOR DI(566) XOR DI(973) XOR DI(970) XOR DI(759) XOR DI(186) XOR DI(835) XOR DI(556) XOR DI(963) XOR DI(960) XOR DI(443) XOR DI(157) XOR DI(642) XOR DI(362) XOR DI(584) XOR DI(708) XOR DI(127) XOR DI(453) XOR DI(167) XOR DI(225) XOR DI(741) XOR DI(609) XOR DI(652) XOR DI(244) XOR DI(499) XOR DI(70) XOR DI(706) XOR DI(637) XOR DI(9) XOR DI(191) XOR DI(914) XOR DI(984) XOR DI(846) XOR DI(111) XOR DI(690) XOR DI(372) XOR DI(486) XOR DI(917) XOR DI(1002) XOR DI(425) XOR DI(802) XOR DI(535) XOR DI(388) XOR DI(178) XOR DI(931) XOR DI(502) XOR DI(594) XOR DI(804) XOR DI(265) XOR DI(230) XOR DI(640) XOR DI(308) XOR DI(12) XOR DI(981) XOR DI(718) XOR DI(270) XOR DI(108) XOR DI(548) XOR DI(945) XOR DI(360) XOR DI(193) XOR DI(933) XOR DI(137) XOR DI(679) XOR DI(1018) XOR DI(764) XOR DI(771) XOR DI(901) XOR DI(441) XOR DI(375) XOR DI(304) XOR DI(567) XOR DI(791) XOR DI(760) XOR DI(729) XOR DI(296) XOR DI(463) XOR DI(177) XOR DI(826) XOR DI(547) XOR DI(235) XOR DI(61) XOR DI(628) XOR DI(0) XOR DI(837) XOR DI(363) XOR DI(526) XOR DI(379) XOR DI(922) XOR DI(221) XOR DI(709) XOR DI(261) XOR DI(128) XOR DI(670) XOR DI(755) XOR DI(892) XOR DI(432) XOR DI(751) XOR DI(287) XOR DI(454) XOR DI(538) XOR DI(226) XOR DI(619) XOR DI(517) XOR DI(252) XOR DI(742) XOR DI(445) XOR DI(217) XOR DI(243) XOR DI(733) XOR DI(884) XOR DI(489) XOR DI(818) XOR DI(893) XOR DI(731) XOR DI(408) XOR DI(638) XOR DI(891) XOR DI(662) XOR DI(20) XOR DI(254) XOR DI(612) XOR DI(330) XOR DI(424) XOR DI(509) XOR DI(470) XOR DI(498) XOR DI(75) XOR DI(857) XOR DI(326) XOR DI(34) XOR DI(160) XOR DI(80) XOR DI(915) XOR DI(827) XOR DI(965) XOR DI(551) XOR DI(428) XOR DI(142) XOR DI(152) XOR DI(691) XOR DI(902) XOR DI(1003) XOR DI(776) XOR DI(113) XOR DI(740) XOR DI(417) XOR DI(228) XOR DI(474) XOR DI(716) XOR DI(647) XOR DI(19) XOR DI(900) XOR DI(179) XOR DI(932) XOR DI(671) XOR DI(29) XOR DI(263) XOR DI(292) XOR DI(36) XOR DI(595) XOR DI(621) XOR DI(404) XOR DI(339) XOR DI(816) XOR DI(433) XOR DI(870) XOR DI(309) XOR DI(288) XOR DI(549) XOR DI(666) XOR DI(946) XOR DI(130) XOR DI(361) XOR DI(150) XOR DI(194) XOR DI(201) XOR DI(620) XOR DI(947) XOR DI(858) XOR DI(518) XOR DI(537) XOR DI(934) XOR DI(138) XOR DI(479) XOR DI(686) XOR DI(507) XOR DI(1019) XOR DI(998) XOR DI(767) XOR DI(84) XOR DI(44) XOR DI(278) XOR DI(866) XOR DI(87) XOR DI(335) XOR DI(328) XOR DI(43) XOR DI(307) XOR DI(570) XOR DI(51) XOR DI(48) XOR DI(169) XOR DI(89) XOR DI(353) XOR DI(687) XOR DI(794) XOR DI(924) XOR DI(836) XOR DI(415) XOR DI(974) XOR DI(763) XOR DI(732) XOR DI(610) XOR DI(47) XOR DI(299) XOR DI(994) XOR DI(856) XOR DI(560) XOR DI(967) XOR DI(180) XOR DI(829) XOR DI(437) XOR DI(151) XOR DI(636) XOR DI(356) XOR DI(578) XOR DI(121) XOR DI(161) XOR DI(219) XOR DI(493) XOR DI(700) XOR DI(3) XOR DI(978) XOR DI(840) XOR DI(684) XOR DI(911) XOR DI(996) XOR DI(419) XOR DI(382) XOR DI(925) XOR DI(496) XOR DI(798) XOR DI(259) XOR DI(224) XOR DI(975) XOR DI(542) XOR DI(354) XOR DI(927) XOR DI(131) XOR DI(1012) XOR DI(435) XOR DI(785) XOR DI(754) XOR DI(723) XOR DI(457) XOR DI(171) XOR DI(820) XOR DI(831) XOR DI(520) XOR DI(373) XOR DI(215) XOR DI(122) XOR DI(749) XOR DI(426) XOR DI(745) XOR DI(281) XOR DI(448) XOR DI(220) XOR DI(246) XOR DI(736) XOR DI(237) XOR DI(483) XOR DI(812) XOR DI(725) XOR DI(402) XOR DI(632) XOR DI(885) XOR DI(656) XOR DI(248) XOR DI(606) XOR DI(324) XOR DI(418) XOR DI(503) XOR DI(69) XOR DI(320) XOR DI(28) XOR DI(154) XOR DI(74) XOR DI(909) XOR DI(821) XOR DI(545) XOR DI(422) XOR DI(896) XOR DI(997) XOR DI(734) XOR DI(411) XOR DI(222) XOR DI(468) XOR DI(710) XOR DI(641) XOR DI(13) XOR DI(894) XOR DI(665) XOR DI(23) XOR DI(286) XOR DI(30) XOR DI(398) XOR DI(333) XOR DI(303) XOR DI(660) XOR DI(124) XOR DI(355) XOR DI(188) XOR DI(614) XOR DI(941) XOR DI(512) XOR DI(132) XOR DI(473) XOR DI(680) XOR DI(78) XOR DI(38) XOR DI(272) XOR DI(301) XOR DI(564) XOR DI(45) XOR DI(681) XOR DI(918) XOR DI(830) XOR DI(409) XOR DI(968) XOR DI(726) XOR DI(604) XOR DI(961) XOR DI(174) XOR DI(145) XOR DI(630) XOR DI(155) XOR DI(213) XOR DI(694) XOR DI(834) XOR DI(905) XOR DI(413) XOR DI(376) XOR DI(218) XOR DI(536) XOR DI(348) XOR DI(125) XOR DI(429) XOR DI(165) XOR DI(814) XOR DI(825) XOR DI(514) XOR DI(209) XOR DI(275) XOR DI(442) XOR DI(214) XOR DI(240) XOR DI(730) XOR DI(477) XOR DI(719) XOR DI(396) XOR DI(879) XOR DI(650) XOR DI(242) XOR DI(318) XOR DI(497) XOR DI(22) XOR DI(68) XOR DI(903) XOR DI(539) XOR DI(416) XOR DI(991) XOR DI(728) XOR DI(405) XOR DI(216) XOR DI(635) XOR DI(7) XOR DI(659) XOR DI(17) XOR DI(280) XOR DI(24) XOR DI(392) XOR DI(327) XOR DI(297) XOR DI(654) XOR DI(118) XOR DI(182) XOR DI(506) XOR DI(126) XOR DI(467) XOR DI(32) XOR DI(266) XOR DI(558) XOR DI(675) XOR DI(912) XOR DI(962) XOR DI(955) XOR DI(168) XOR DI(139) XOR DI(624) XOR DI(149) XOR DI(370) XOR DI(212) XOR DI(342) XOR DI(159) XOR DI(819) XOR DI(203) XOR DI(436) XOR DI(471) XOR DI(713) XOR DI(873) XOR DI(16) XOR DI(533) XOR DI(399) XOR DI(210) XOR DI(629) XOR DI(386) XOR DI(321) XOR DI(500) XOR DI(461) XOR DI(552) XOR DI(669) XOR DI(956) XOR DI(949) XOR DI(153) XOR DI(465) XOR DI(707) XOR DI(867) XOR DI(10) XOR DI(527) XOR DI(204) XOR DI(623) XOR DI(380) XOR DI(494) XOR DI(455) XOR DI(546) XOR DI(943) XOR DI(147) XOR DI(701) XOR DI(861) XOR DI(4) XOR DI(521) XOR DI(488) XOR DI(540) XOR DI(141) XOR DI(695) XOR DI(534) XOR DI(135) XOR DI(689) XOR DI(528) XOR DI(129) XOR DI(683) XOR DI(522) XOR DI(516) XOR DI(510) XOR DI(1016) XOR DI(1022);
   DO(5) <= DI(581) XOR DI(274) XOR DI(1005) XOR DI(47) XOR DI(753) XOR DI(359) XOR DI(592) XOR DI(774) XOR DI(781) XOR DI(911) XOR DI(91) XOR DI(51) XOR DI(285) XOR DI(873) XOR DI(712) XOR DI(593) XOR DI(451) XOR DI(307) XOR DI(94) XOR DI(385) XOR DI(342) XOR DI(839) XOR DI(1000) XOR DI(335) XOR DI(50) XOR DI(802) XOR DI(314) XOR DI(190) XOR DI(860) XOR DI(577) XOR DI(984) XOR DI(564) XOR DI(58) XOR DI(95) XOR DI(945) XOR DI(55) XOR DI(176) XOR DI(96) XOR DI(930) XOR DI(360) XOR DI(694) XOR DI(878) XOR DI(98) XOR DI(580) XOR DI(801) XOR DI(931) XOR DI(843) XOR DI(74) XOR DI(338) XOR DI(422) XOR DI(981) XOR DI(770) XOR DI(739) XOR DI(617) XOR DI(54) XOR DI(111) XOR DI(197) XOR DI(306) XOR DI(846) XOR DI(473) XOR DI(1001) XOR DI(863) XOR DI(567) XOR DI(974) XOR DI(971) XOR DI(760) XOR DI(187) XOR DI(836) XOR DI(557) XOR DI(964) XOR DI(961) XOR DI(444) XOR DI(158) XOR DI(643) XOR DI(0) XOR DI(363) XOR DI(585) XOR DI(709) XOR DI(128) XOR DI(454) XOR DI(168) XOR DI(226) XOR DI(742) XOR DI(610) XOR DI(653) XOR DI(245) XOR DI(500) XOR DI(71) XOR DI(707) XOR DI(638) XOR DI(10) XOR DI(192) XOR DI(915) XOR DI(985) XOR DI(847) XOR DI(112) XOR DI(691) XOR DI(373) XOR DI(487) XOR DI(918) XOR DI(1003) XOR DI(426) XOR DI(803) XOR DI(536) XOR DI(389) XOR DI(179) XOR DI(932) XOR DI(503) XOR DI(595) XOR DI(805) XOR DI(266) XOR DI(231) XOR DI(641) XOR DI(309) XOR DI(13) XOR DI(982) XOR DI(719) XOR DI(271) XOR DI(109) XOR DI(549) XOR DI(946) XOR DI(361) XOR DI(194) XOR DI(934) XOR DI(138) XOR DI(680) XOR DI(1019) XOR DI(765) XOR DI(772) XOR DI(902) XOR DI(442) XOR DI(376) XOR DI(305) XOR DI(568) XOR DI(792) XOR DI(761) XOR DI(730) XOR DI(297) XOR DI(464) XOR DI(178) XOR DI(827) XOR DI(548) XOR DI(236) XOR DI(62) XOR DI(629) XOR DI(1) XOR DI(838) XOR DI(364) XOR DI(527) XOR DI(380) XOR DI(923) XOR DI(222) XOR DI(710) XOR DI(262) XOR DI(129) XOR DI(671) XOR DI(756) XOR DI(893) XOR DI(433) XOR DI(752) XOR DI(288) XOR DI(455) XOR DI(539) XOR DI(227) XOR DI(620) XOR DI(518) XOR DI(253) XOR DI(743) XOR DI(446) XOR DI(218) XOR DI(244) XOR DI(734) XOR DI(885) XOR DI(490) XOR DI(819) XOR DI(894) XOR DI(732) XOR DI(409) XOR DI(639) XOR DI(892) XOR DI(663) XOR DI(21) XOR DI(255) XOR DI(613) XOR DI(331) XOR DI(425) XOR DI(510) XOR DI(471) XOR DI(499) XOR DI(76) XOR DI(858) XOR DI(327) XOR DI(35) XOR DI(161) XOR DI(81) XOR DI(916) XOR DI(828) XOR DI(966) XOR DI(552) XOR DI(429) XOR DI(143) XOR DI(153) XOR DI(692) XOR DI(903) XOR DI(1004) XOR DI(777) XOR DI(114) XOR DI(741) XOR DI(418) XOR DI(229) XOR DI(475) XOR DI(717) XOR DI(648) XOR DI(20) XOR DI(901) XOR DI(180) XOR DI(933) XOR DI(672) XOR DI(30) XOR DI(264) XOR DI(293) XOR DI(37) XOR DI(596) XOR DI(622) XOR DI(405) XOR DI(340) XOR DI(817) XOR DI(434) XOR DI(871) XOR DI(310) XOR DI(289) XOR DI(550) XOR DI(667) XOR DI(947) XOR DI(131) XOR DI(362) XOR DI(151) XOR DI(195) XOR DI(202) XOR DI(621) XOR DI(948) XOR DI(859) XOR DI(519) XOR DI(538) XOR DI(935) XOR DI(139) XOR DI(480) XOR DI(687) XOR DI(508) XOR DI(1020) XOR DI(999) XOR DI(768) XOR DI(85) XOR DI(45) XOR DI(279) XOR DI(867) XOR DI(88) XOR DI(336) XOR DI(329) XOR DI(44) XOR DI(308) XOR DI(571) XOR DI(52) XOR DI(49) XOR DI(170) XOR DI(90) XOR DI(354) XOR DI(688) XOR DI(795) XOR DI(925) XOR DI(837) XOR DI(416) XOR DI(975) XOR DI(764) XOR DI(733) XOR DI(611) XOR DI(48) XOR DI(300) XOR DI(995) XOR DI(857) XOR DI(561) XOR DI(968) XOR DI(181) XOR DI(830) XOR DI(438) XOR DI(152) XOR DI(637) XOR DI(357) XOR DI(579) XOR DI(122) XOR DI(162) XOR DI(220) XOR DI(494) XOR DI(701) XOR DI(4) XOR DI(979) XOR DI(841) XOR DI(685) XOR DI(912) XOR DI(997) XOR DI(420) XOR DI(383) XOR DI(926) XOR DI(497) XOR DI(799) XOR DI(260) XOR DI(225) XOR DI(976) XOR DI(543) XOR DI(355) XOR DI(928) XOR DI(132) XOR DI(1013) XOR DI(436) XOR DI(786) XOR DI(755) XOR DI(724) XOR DI(458) XOR DI(172) XOR DI(821) XOR DI(832) XOR DI(521) XOR DI(374) XOR DI(216) XOR DI(123) XOR DI(750) XOR DI(427) XOR DI(746) XOR DI(282) XOR DI(449) XOR DI(221) XOR DI(247) XOR DI(737) XOR DI(238) XOR DI(484) XOR DI(813) XOR DI(726) XOR DI(403) XOR DI(633) XOR DI(886) XOR DI(657) XOR DI(249) XOR DI(607) XOR DI(325) XOR DI(419) XOR DI(504) XOR DI(70) XOR DI(321) XOR DI(29) XOR DI(155) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(546) XOR DI(423) XOR DI(897) XOR DI(998) XOR DI(735) XOR DI(412) XOR DI(223) XOR DI(469) XOR DI(711) XOR DI(642) XOR DI(14) XOR DI(895) XOR DI(666) XOR DI(24) XOR DI(287) XOR DI(31) XOR DI(399) XOR DI(334) XOR DI(304) XOR DI(661) XOR DI(125) XOR DI(356) XOR DI(189) XOR DI(615) XOR DI(942) XOR DI(513) XOR DI(133) XOR DI(474) XOR DI(681) XOR DI(79) XOR DI(39) XOR DI(273) XOR DI(302) XOR DI(565) XOR DI(46) XOR DI(682) XOR DI(919) XOR DI(831) XOR DI(410) XOR DI(969) XOR DI(727) XOR DI(605) XOR DI(962) XOR DI(175) XOR DI(146) XOR DI(631) XOR DI(156) XOR DI(214) XOR DI(695) XOR DI(835) XOR DI(906) XOR DI(414) XOR DI(377) XOR DI(219) XOR DI(537) XOR DI(349) XOR DI(126) XOR DI(430) XOR DI(166) XOR DI(815) XOR DI(826) XOR DI(515) XOR DI(210) XOR DI(276) XOR DI(443) XOR DI(215) XOR DI(241) XOR DI(731) XOR DI(478) XOR DI(720) XOR DI(397) XOR DI(880) XOR DI(651) XOR DI(243) XOR DI(319) XOR DI(498) XOR DI(23) XOR DI(69) XOR DI(904) XOR DI(540) XOR DI(417) XOR DI(992) XOR DI(729) XOR DI(406) XOR DI(217) XOR DI(636) XOR DI(8) XOR DI(660) XOR DI(18) XOR DI(281) XOR DI(25) XOR DI(393) XOR DI(328) XOR DI(298) XOR DI(655) XOR DI(119) XOR DI(183) XOR DI(507) XOR DI(127) XOR DI(468) XOR DI(33) XOR DI(267) XOR DI(559) XOR DI(676) XOR DI(913) XOR DI(963) XOR DI(956) XOR DI(169) XOR DI(140) XOR DI(625) XOR DI(150) XOR DI(371) XOR DI(213) XOR DI(343) XOR DI(160) XOR DI(820) XOR DI(204) XOR DI(437) XOR DI(472) XOR DI(714) XOR DI(874) XOR DI(17) XOR DI(534) XOR DI(400) XOR DI(211) XOR DI(630) XOR DI(387) XOR DI(322) XOR DI(501) XOR DI(462) XOR DI(553) XOR DI(670) XOR DI(957) XOR DI(950) XOR DI(154) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(11) XOR DI(528) XOR DI(205) XOR DI(624) XOR DI(381) XOR DI(495) XOR DI(456) XOR DI(547) XOR DI(944) XOR DI(148) XOR DI(702) XOR DI(862) XOR DI(5) XOR DI(522) XOR DI(489) XOR DI(541) XOR DI(142) XOR DI(696) XOR DI(535) XOR DI(136) XOR DI(690) XOR DI(529) XOR DI(130) XOR DI(684) XOR DI(523) XOR DI(517) XOR DI(511) XOR DI(1017) XOR DI(1023);
   DO(6) <= DI(231) XOR DI(582) XOR DI(275) XOR DI(1006) XOR DI(857) XOR DI(825) XOR DI(48) XOR DI(754) XOR DI(74) XOR DI(781) XOR DI(575) XOR DI(360) XOR DI(593) XOR DI(775) XOR DI(890) XOR DI(650) XOR DI(574) XOR DI(432) XOR DI(841) XOR DI(782) XOR DI(912) XOR DI(92) XOR DI(690) XOR DI(109) XOR DI(591) XOR DI(52) XOR DI(619) XOR DI(93) XOR DI(468) XOR DI(899) XOR DI(517) XOR DI(286) XOR DI(874) XOR DI(269) XOR DI(713) XOR DI(873) XOR DI(594) XOR DI(452) XOR DI(57) XOR DI(308) XOR DI(95) XOR DI(386) XOR DI(928) XOR DI(343) XOR DI(840) XOR DI(1001) XOR DI(69) XOR DI(776) XOR DI(338) XOR DI(336) XOR DI(767) XOR DI(707) XOR DI(51) XOR DI(803) XOR DI(979) XOR DI(315) XOR DI(191) XOR DI(861) XOR DI(324) XOR DI(192) XOR DI(578) XOR DI(985) XOR DI(930) XOR DI(565) XOR DI(59) XOR DI(96) XOR DI(946) XOR DI(56) XOR DI(177) XOR DI(97) XOR DI(931) XOR DI(665) XOR DI(750) XOR DI(361) XOR DI(695) XOR DI(879) XOR DI(484) XOR DI(99) XOR DI(165) XOR DI(581) XOR DI(802) XOR DI(932) XOR DI(844) XOR DI(75) XOR DI(339) XOR DI(815) XOR DI(423) XOR DI(107) XOR DI(982) XOR DI(771) XOR DI(740) XOR DI(359) XOR DI(798) XOR DI(618) XOR DI(55) XOR DI(880) XOR DI(600) XOR DI(666) XOR DI(64) XOR DI(590) XOR DI(199) XOR DI(200) XOR DI(636) XOR DI(304) XOR DI(714) XOR DI(112) XOR DI(610) XOR DI(198) XOR DI(307) XOR DI(451) XOR DI(847) XOR DI(474) XOR DI(1002) XOR DI(772) XOR DI(276) XOR DI(864) XOR DI(85) XOR DI(376) XOR DI(333) XOR DI(568) XOR DI(975) XOR DI(921) XOR DI(834) XOR DI(65) XOR DI(972) XOR DI(761) XOR DI(188) XOR DI(837) XOR DI(558) XOR DI(965) XOR DI(962) XOR DI(178) XOR DI(952) XOR DI(576) XOR DI(445) XOR DI(159) XOR DI(644) XOR DI(1) XOR DI(906) XOR DI(364) XOR DI(994) XOR DI(380) XOR DI(494) XOR DI(586) XOR DI(257) XOR DI(710) XOR DI(262) XOR DI(185) XOR DI(129) XOR DI(763) XOR DI(433) XOR DI(455) XOR DI(169) XOR DI(227) XOR DI(620) XOR DI(371) XOR DI(743) XOR DI(611) XOR DI(810) XOR DI(654) XOR DI(246) XOR DI(501) XOR DI(72) XOR DI(543) XOR DI(708) XOR DI(639) XOR DI(11) XOR DI(892) XOR DI(255) XOR DI(284) XOR DI(28) XOR DI(331) XOR DI(808) XOR DI(862) XOR DI(193) XOR DI(759) XOR DI(916) XOR DI(755) XOR DI(986) XOR DI(848) XOR DI(552) XOR DI(959) XOR DI(113) XOR DI(692) XOR DI(374) XOR DI(488) XOR DI(790) XOR DI(534) XOR DI(919) XOR DI(1004) XOR DI(427) XOR DI(449) XOR DI(741) XOR DI(737) XOR DI(238) XOR DI(804) XOR DI(624) XOR DI(648) XOR DI(240) XOR DI(316) XOR DI(20) XOR DI(901) XOR DI(537) XOR DI(888) XOR DI(390) XOR DI(295) XOR DI(180) XOR DI(933) XOR DI(504) XOR DI(293) XOR DI(596) XOR DI(826) XOR DI(897) XOR DI(405) XOR DI(806) XOR DI(817) XOR DI(506) XOR DI(267) XOR DI(232) XOR DI(642) XOR DI(310) XOR DI(14) XOR DI(983) XOR DI(720) XOR DI(272) XOR DI(646) XOR DI(110) XOR DI(174) XOR DI(550) XOR DI(947) XOR DI(362) XOR DI(195) XOR DI(705) XOR DI(8) XOR DI(453) XOR DI(941) XOR DI(615) XOR DI(935) XOR DI(139) XOR DI(853) XOR DI(681) XOR DI(675) XOR DI(1008) XOR DI(1020) XOR DI(266) XOR DI(39) XOR DI(745) XOR DI(351) XOR DI(766) XOR DI(773) XOR DI(903) XOR DI(83) XOR DI(43) XOR DI(704) XOR DI(443) XOR DI(377) XOR DI(992) XOR DI(42) XOR DI(794) XOR DI(306) XOR DI(852) XOR DI(569) XOR DI(556) XOR DI(937) XOR DI(352) XOR DI(90) XOR DI(793) XOR DI(923) XOR DI(66) XOR DI(414) XOR DI(762) XOR DI(731) XOR DI(189) XOR DI(298) XOR DI(465) XOR DI(855) XOR DI(559) XOR DI(966) XOR DI(179) XOR DI(828) XOR DI(549) XOR DI(956) XOR DI(150) XOR DI(446) XOR DI(602) XOR DI(237) XOR DI(492) XOR DI(63) XOR DI(630) XOR DI(2) XOR DI(839) XOR DI(104) XOR DI(365) XOR DI(910) XOR DI(995) XOR DI(528) XOR DI(381) XOR DI(924) XOR DI(587) XOR DI(797) XOR DI(223) XOR DI(633) XOR DI(974) XOR DI(711) XOR DI(263) XOR DI(130) XOR DI(672) XOR DI(757) XOR DI(894) XOR DI(434) XOR DI(368) XOR DI(297) XOR DI(753) XOR DI(722) XOR DI(289) XOR DI(456) XOR DI(540) XOR DI(228) XOR DI(621) XOR DI(830) XOR DI(519) XOR DI(254) XOR DI(121) XOR DI(748) XOR DI(425) XOR DI(744) XOR DI(447) XOR DI(531) XOR DI(219) XOR DI(510) XOR DI(245) XOR DI(735) XOR DI(210) XOR DI(236) XOR DI(726) XOR DI(482) XOR DI(886) XOR DI(724) XOR DI(655) XOR DI(13) XOR DI(605) XOR DI(491) XOR DI(908) XOR DI(820) XOR DI(135) XOR DI(145) XOR DI(895) XOR DI(106) XOR DI(733) XOR DI(410) XOR DI(640) XOR DI(893) XOR DI(925) XOR DI(664) XOR DI(22) XOR DI(256) XOR DI(588) XOR DI(614) XOR DI(332) XOR DI(426) XOR DI(302) XOR DI(939) XOR DI(354) XOR DI(187) XOR DI(940) XOR DI(511) XOR DI(472) XOR DI(679) XOR DI(500) XOR DI(1012) XOR DI(760) XOR DI(77) XOR DI(271) XOR DI(859) XOR DI(328) XOR DI(36) XOR DI(300) XOR DI(563) XOR DI(44) XOR DI(41) XOR DI(162) XOR DI(82) XOR DI(680) XOR DI(917) XOR DI(829) XOR DI(967) XOR DI(292) XOR DI(987) XOR DI(553) XOR DI(430) XOR DI(144) XOR DI(349) XOR DI(114) XOR DI(154) XOR DI(693) XOR DI(971) XOR DI(904) XOR DI(412) XOR DI(918) XOR DI(489) XOR DI(1005) XOR DI(778) XOR DI(164) XOR DI(513) XOR DI(366) XOR DI(208) XOR DI(115) XOR DI(742) XOR DI(419) XOR DI(441) XOR DI(213) XOR DI(729) XOR DI(230) XOR DI(476) XOR DI(718) XOR DI(395) XOR DI(649) XOR DI(317) XOR DI(21) XOR DI(902) XOR DI(889) XOR DI(990) XOR DI(461) XOR DI(16) XOR DI(117) XOR DI(181) XOR DI(934) XOR DI(125) XOR DI(466) XOR DI(673) XOR DI(31) XOR DI(265) XOR DI(294) XOR DI(38) XOR DI(961) XOR DI(719) XOR DI(597) XOR DI(138) XOR DI(623) XOR DI(148) XOR DI(687) XOR DI(406) XOR DI(369) XOR DI(341) XOR DI(118) XOR DI(422) XOR DI(818) XOR DI(435) XOR DI(233) XOR DI(872) XOR DI(311) XOR DI(532) XOR DI(409) XOR DI(209) XOR DI(628) XOR DI(290) XOR DI(175) XOR DI(259) XOR DI(551) XOR DI(668) XOR DI(948) XOR DI(132) XOR DI(617) XOR DI(363) XOR DI(152) XOR DI(812) XOR DI(196) XOR DI(429) XOR DI(464) XOR DI(706) XOR DI(866) XOR DI(392) XOR DI(203) XOR DI(622) XOR DI(314) XOR DI(493) XOR DI(545) XOR DI(949) XOR DI(942) XOR DI(146) XOR DI(860) XOR DI(3) XOR DI(520) XOR DI(197) XOR DI(539) XOR DI(936) XOR DI(140) XOR DI(854) XOR DI(481) XOR DI(533) XOR DI(688) XOR DI(122) XOR DI(676) XOR DI(509) XOR DI(503) XOR DI(1015) XOR DI(1021);
   DO(7) <= DI(232) XOR DI(583) XOR DI(276) XOR DI(1007) XOR DI(858) XOR DI(826) XOR DI(49) XOR DI(755) XOR DI(75) XOR DI(782) XOR DI(576) XOR DI(361) XOR DI(594) XOR DI(776) XOR DI(891) XOR DI(651) XOR DI(575) XOR DI(433) XOR DI(842) XOR DI(783) XOR DI(913) XOR DI(93) XOR DI(691) XOR DI(110) XOR DI(592) XOR DI(53) XOR DI(620) XOR DI(94) XOR DI(469) XOR DI(900) XOR DI(518) XOR DI(287) XOR DI(875) XOR DI(270) XOR DI(714) XOR DI(874) XOR DI(595) XOR DI(453) XOR DI(58) XOR DI(309) XOR DI(96) XOR DI(387) XOR DI(929) XOR DI(344) XOR DI(841) XOR DI(1002) XOR DI(70) XOR DI(777) XOR DI(339) XOR DI(337) XOR DI(768) XOR DI(708) XOR DI(52) XOR DI(804) XOR DI(980) XOR DI(316) XOR DI(192) XOR DI(862) XOR DI(325) XOR DI(193) XOR DI(579) XOR DI(986) XOR DI(931) XOR DI(566) XOR DI(60) XOR DI(97) XOR DI(947) XOR DI(57) XOR DI(178) XOR DI(98) XOR DI(932) XOR DI(666) XOR DI(751) XOR DI(362) XOR DI(696) XOR DI(880) XOR DI(485) XOR DI(100) XOR DI(166) XOR DI(582) XOR DI(803) XOR DI(933) XOR DI(845) XOR DI(76) XOR DI(340) XOR DI(816) XOR DI(424) XOR DI(108) XOR DI(983) XOR DI(772) XOR DI(741) XOR DI(360) XOR DI(799) XOR DI(619) XOR DI(56) XOR DI(881) XOR DI(601) XOR DI(667) XOR DI(65) XOR DI(591) XOR DI(200) XOR DI(201) XOR DI(637) XOR DI(305) XOR DI(715) XOR DI(113) XOR DI(611) XOR DI(199) XOR DI(308) XOR DI(452) XOR DI(848) XOR DI(475) XOR DI(1003) XOR DI(773) XOR DI(277) XOR DI(865) XOR DI(86) XOR DI(377) XOR DI(334) XOR DI(569) XOR DI(976) XOR DI(922) XOR DI(835) XOR DI(66) XOR DI(973) XOR DI(762) XOR DI(189) XOR DI(838) XOR DI(559) XOR DI(966) XOR DI(963) XOR DI(179) XOR DI(953) XOR DI(577) XOR DI(446) XOR DI(160) XOR DI(645) XOR DI(2) XOR DI(907) XOR DI(365) XOR DI(995) XOR DI(381) XOR DI(495) XOR DI(587) XOR DI(258) XOR DI(711) XOR DI(263) XOR DI(186) XOR DI(130) XOR DI(764) XOR DI(434) XOR DI(456) XOR DI(170) XOR DI(228) XOR DI(621) XOR DI(372) XOR DI(744) XOR DI(612) XOR DI(811) XOR DI(655) XOR DI(247) XOR DI(502) XOR DI(73) XOR DI(544) XOR DI(709) XOR DI(640) XOR DI(12) XOR DI(893) XOR DI(256) XOR DI(285) XOR DI(29) XOR DI(332) XOR DI(809) XOR DI(863) XOR DI(194) XOR DI(760) XOR DI(917) XOR DI(756) XOR DI(987) XOR DI(849) XOR DI(553) XOR DI(960) XOR DI(114) XOR DI(693) XOR DI(375) XOR DI(489) XOR DI(791) XOR DI(535) XOR DI(920) XOR DI(1005) XOR DI(428) XOR DI(450) XOR DI(742) XOR DI(738) XOR DI(239) XOR DI(805) XOR DI(625) XOR DI(649) XOR DI(241) XOR DI(317) XOR DI(21) XOR DI(902) XOR DI(538) XOR DI(889) XOR DI(391) XOR DI(296) XOR DI(181) XOR DI(934) XOR DI(505) XOR DI(294) XOR DI(597) XOR DI(827) XOR DI(898) XOR DI(406) XOR DI(807) XOR DI(818) XOR DI(507) XOR DI(268) XOR DI(233) XOR DI(643) XOR DI(311) XOR DI(15) XOR DI(984) XOR DI(721) XOR DI(273) XOR DI(647) XOR DI(111) XOR DI(175) XOR DI(551) XOR DI(948) XOR DI(363) XOR DI(196) XOR DI(706) XOR DI(9) XOR DI(454) XOR DI(942) XOR DI(616) XOR DI(936) XOR DI(140) XOR DI(854) XOR DI(682) XOR DI(676) XOR DI(1009) XOR DI(1021) XOR DI(267) XOR DI(40) XOR DI(746) XOR DI(352) XOR DI(767) XOR DI(774) XOR DI(904) XOR DI(84) XOR DI(44) XOR DI(705) XOR DI(444) XOR DI(378) XOR DI(993) XOR DI(43) XOR DI(795) XOR DI(307) XOR DI(853) XOR DI(570) XOR DI(557) XOR DI(938) XOR DI(353) XOR DI(91) XOR DI(794) XOR DI(924) XOR DI(67) XOR DI(415) XOR DI(763) XOR DI(732) XOR DI(190) XOR DI(299) XOR DI(466) XOR DI(856) XOR DI(560) XOR DI(967) XOR DI(180) XOR DI(829) XOR DI(550) XOR DI(957) XOR DI(151) XOR DI(447) XOR DI(603) XOR DI(238) XOR DI(493) XOR DI(64) XOR DI(631) XOR DI(3) XOR DI(840) XOR DI(105) XOR DI(366) XOR DI(911) XOR DI(996) XOR DI(529) XOR DI(382) XOR DI(925) XOR DI(588) XOR DI(798) XOR DI(224) XOR DI(634) XOR DI(975) XOR DI(712) XOR DI(264) XOR DI(131) XOR DI(673) XOR DI(758) XOR DI(895) XOR DI(435) XOR DI(369) XOR DI(298) XOR DI(754) XOR DI(723) XOR DI(290) XOR DI(457) XOR DI(541) XOR DI(229) XOR DI(622) XOR DI(831) XOR DI(520) XOR DI(255) XOR DI(122) XOR DI(749) XOR DI(426) XOR DI(745) XOR DI(448) XOR DI(532) XOR DI(220) XOR DI(511) XOR DI(246) XOR DI(736) XOR DI(211) XOR DI(237) XOR DI(727) XOR DI(483) XOR DI(887) XOR DI(725) XOR DI(656) XOR DI(14) XOR DI(606) XOR DI(492) XOR DI(909) XOR DI(821) XOR DI(136) XOR DI(146) XOR DI(896) XOR DI(107) XOR DI(734) XOR DI(411) XOR DI(641) XOR DI(894) XOR DI(926) XOR DI(665) XOR DI(23) XOR DI(257) XOR DI(589) XOR DI(615) XOR DI(333) XOR DI(427) XOR DI(303) XOR DI(940) XOR DI(355) XOR DI(188) XOR DI(941) XOR DI(512) XOR DI(473) XOR DI(680) XOR DI(501) XOR DI(1013) XOR DI(761) XOR DI(78) XOR DI(272) XOR DI(860) XOR DI(329) XOR DI(37) XOR DI(301) XOR DI(564) XOR DI(45) XOR DI(42) XOR DI(163) XOR DI(83) XOR DI(681) XOR DI(918) XOR DI(830) XOR DI(968) XOR DI(293) XOR DI(988) XOR DI(554) XOR DI(431) XOR DI(145) XOR DI(350) XOR DI(115) XOR DI(155) XOR DI(694) XOR DI(972) XOR DI(905) XOR DI(413) XOR DI(919) XOR DI(490) XOR DI(1006) XOR DI(779) XOR DI(165) XOR DI(514) XOR DI(367) XOR DI(209) XOR DI(116) XOR DI(743) XOR DI(420) XOR DI(442) XOR DI(214) XOR DI(730) XOR DI(231) XOR DI(477) XOR DI(719) XOR DI(396) XOR DI(650) XOR DI(318) XOR DI(22) XOR DI(903) XOR DI(890) XOR DI(991) XOR DI(462) XOR DI(17) XOR DI(118) XOR DI(182) XOR DI(935) XOR DI(126) XOR DI(467) XOR DI(674) XOR DI(32) XOR DI(266) XOR DI(295) XOR DI(39) XOR DI(962) XOR DI(720) XOR DI(598) XOR DI(139) XOR DI(624) XOR DI(149) XOR DI(688) XOR DI(407) XOR DI(370) XOR DI(342) XOR DI(119) XOR DI(423) XOR DI(819) XOR DI(436) XOR DI(234) XOR DI(873) XOR DI(312) XOR DI(533) XOR DI(410) XOR DI(210) XOR DI(629) XOR DI(291) XOR DI(176) XOR DI(260) XOR DI(552) XOR DI(669) XOR DI(949) XOR DI(133) XOR DI(618) XOR DI(364) XOR DI(153) XOR DI(813) XOR DI(197) XOR DI(430) XOR DI(465) XOR DI(707) XOR DI(867) XOR DI(393) XOR DI(204) XOR DI(623) XOR DI(315) XOR DI(494) XOR DI(546) XOR DI(950) XOR DI(943) XOR DI(147) XOR DI(861) XOR DI(4) XOR DI(521) XOR DI(198) XOR DI(540) XOR DI(937) XOR DI(141) XOR DI(855) XOR DI(482) XOR DI(534) XOR DI(689) XOR DI(123) XOR DI(677) XOR DI(510) XOR DI(504) XOR DI(1016) XOR DI(1022);
   DO(8) <= DI(233) XOR DI(584) XOR DI(277) XOR DI(1008) XOR DI(859) XOR DI(827) XOR DI(50) XOR DI(756) XOR DI(76) XOR DI(783) XOR DI(577) XOR DI(362) XOR DI(595) XOR DI(777) XOR DI(892) XOR DI(652) XOR DI(576) XOR DI(434) XOR DI(843) XOR DI(784) XOR DI(914) XOR DI(94) XOR DI(692) XOR DI(111) XOR DI(593) XOR DI(54) XOR DI(621) XOR DI(95) XOR DI(470) XOR DI(901) XOR DI(519) XOR DI(288) XOR DI(876) XOR DI(271) XOR DI(715) XOR DI(875) XOR DI(596) XOR DI(454) XOR DI(59) XOR DI(310) XOR DI(97) XOR DI(388) XOR DI(930) XOR DI(345) XOR DI(842) XOR DI(1003) XOR DI(71) XOR DI(778) XOR DI(340) XOR DI(338) XOR DI(769) XOR DI(709) XOR DI(53) XOR DI(805) XOR DI(981) XOR DI(317) XOR DI(193) XOR DI(863) XOR DI(326) XOR DI(194) XOR DI(580) XOR DI(987) XOR DI(932) XOR DI(567) XOR DI(61) XOR DI(98) XOR DI(948) XOR DI(58) XOR DI(179) XOR DI(99) XOR DI(0) XOR DI(933) XOR DI(667) XOR DI(752) XOR DI(363) XOR DI(697) XOR DI(881) XOR DI(486) XOR DI(101) XOR DI(167) XOR DI(583) XOR DI(804) XOR DI(934) XOR DI(846) XOR DI(77) XOR DI(341) XOR DI(817) XOR DI(425) XOR DI(109) XOR DI(984) XOR DI(773) XOR DI(742) XOR DI(361) XOR DI(800) XOR DI(620) XOR DI(57) XOR DI(882) XOR DI(602) XOR DI(668) XOR DI(66) XOR DI(592) XOR DI(201) XOR DI(202) XOR DI(638) XOR DI(306) XOR DI(716) XOR DI(114) XOR DI(612) XOR DI(200) XOR DI(309) XOR DI(453) XOR DI(849) XOR DI(476) XOR DI(1004) XOR DI(774) XOR DI(278) XOR DI(866) XOR DI(87) XOR DI(378) XOR DI(335) XOR DI(570) XOR DI(977) XOR DI(923) XOR DI(836) XOR DI(67) XOR DI(974) XOR DI(763) XOR DI(190) XOR DI(839) XOR DI(560) XOR DI(967) XOR DI(964) XOR DI(180) XOR DI(954) XOR DI(578) XOR DI(447) XOR DI(161) XOR DI(646) XOR DI(3) XOR DI(908) XOR DI(366) XOR DI(996) XOR DI(382) XOR DI(496) XOR DI(588) XOR DI(259) XOR DI(712) XOR DI(264) XOR DI(187) XOR DI(131) XOR DI(765) XOR DI(435) XOR DI(457) XOR DI(171) XOR DI(229) XOR DI(622) XOR DI(373) XOR DI(745) XOR DI(613) XOR DI(812) XOR DI(656) XOR DI(248) XOR DI(503) XOR DI(74) XOR DI(545) XOR DI(710) XOR DI(641) XOR DI(13) XOR DI(894) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(333) XOR DI(810) XOR DI(864) XOR DI(195) XOR DI(761) XOR DI(918) XOR DI(757) XOR DI(988) XOR DI(850) XOR DI(554) XOR DI(961) XOR DI(115) XOR DI(694) XOR DI(376) XOR DI(490) XOR DI(792) XOR DI(536) XOR DI(921) XOR DI(1006) XOR DI(429) XOR DI(451) XOR DI(743) XOR DI(739) XOR DI(240) XOR DI(806) XOR DI(626) XOR DI(650) XOR DI(242) XOR DI(318) XOR DI(22) XOR DI(903) XOR DI(539) XOR DI(890) XOR DI(392) XOR DI(297) XOR DI(182) XOR DI(935) XOR DI(506) XOR DI(295) XOR DI(598) XOR DI(828) XOR DI(899) XOR DI(407) XOR DI(808) XOR DI(819) XOR DI(508) XOR DI(269) XOR DI(234) XOR DI(644) XOR DI(312) XOR DI(16) XOR DI(985) XOR DI(722) XOR DI(274) XOR DI(648) XOR DI(112) XOR DI(176) XOR DI(552) XOR DI(949) XOR DI(364) XOR DI(197) XOR DI(707) XOR DI(10) XOR DI(455) XOR DI(943) XOR DI(617) XOR DI(937) XOR DI(141) XOR DI(855) XOR DI(683) XOR DI(677) XOR DI(1010) XOR DI(1022) XOR DI(268) XOR DI(41) XOR DI(747) XOR DI(353) XOR DI(768) XOR DI(775) XOR DI(905) XOR DI(85) XOR DI(45) XOR DI(706) XOR DI(445) XOR DI(379) XOR DI(994) XOR DI(44) XOR DI(796) XOR DI(308) XOR DI(854) XOR DI(571) XOR DI(558) XOR DI(939) XOR DI(354) XOR DI(92) XOR DI(795) XOR DI(925) XOR DI(68) XOR DI(416) XOR DI(764) XOR DI(733) XOR DI(191) XOR DI(300) XOR DI(467) XOR DI(857) XOR DI(561) XOR DI(968) XOR DI(181) XOR DI(830) XOR DI(551) XOR DI(958) XOR DI(152) XOR DI(448) XOR DI(604) XOR DI(239) XOR DI(494) XOR DI(65) XOR DI(632) XOR DI(4) XOR DI(841) XOR DI(106) XOR DI(367) XOR DI(912) XOR DI(997) XOR DI(530) XOR DI(383) XOR DI(926) XOR DI(589) XOR DI(799) XOR DI(225) XOR DI(635) XOR DI(976) XOR DI(713) XOR DI(265) XOR DI(132) XOR DI(674) XOR DI(759) XOR DI(896) XOR DI(436) XOR DI(370) XOR DI(299) XOR DI(755) XOR DI(724) XOR DI(291) XOR DI(458) XOR DI(542) XOR DI(230) XOR DI(623) XOR DI(832) XOR DI(521) XOR DI(256) XOR DI(123) XOR DI(750) XOR DI(427) XOR DI(746) XOR DI(449) XOR DI(533) XOR DI(221) XOR DI(512) XOR DI(247) XOR DI(737) XOR DI(212) XOR DI(238) XOR DI(728) XOR DI(484) XOR DI(888) XOR DI(726) XOR DI(657) XOR DI(15) XOR DI(607) XOR DI(493) XOR DI(910) XOR DI(822) XOR DI(137) XOR DI(147) XOR DI(897) XOR DI(108) XOR DI(735) XOR DI(412) XOR DI(642) XOR DI(895) XOR DI(927) XOR DI(666) XOR DI(24) XOR DI(258) XOR DI(590) XOR DI(616) XOR DI(334) XOR DI(428) XOR DI(304) XOR DI(941) XOR DI(356) XOR DI(189) XOR DI(942) XOR DI(513) XOR DI(474) XOR DI(681) XOR DI(502) XOR DI(1014) XOR DI(762) XOR DI(79) XOR DI(273) XOR DI(861) XOR DI(330) XOR DI(38) XOR DI(302) XOR DI(565) XOR DI(46) XOR DI(43) XOR DI(164) XOR DI(84) XOR DI(682) XOR DI(919) XOR DI(831) XOR DI(969) XOR DI(294) XOR DI(989) XOR DI(555) XOR DI(432) XOR DI(146) XOR DI(351) XOR DI(116) XOR DI(156) XOR DI(695) XOR DI(973) XOR DI(906) XOR DI(414) XOR DI(920) XOR DI(491) XOR DI(1007) XOR DI(780) XOR DI(166) XOR DI(515) XOR DI(368) XOR DI(210) XOR DI(117) XOR DI(744) XOR DI(421) XOR DI(443) XOR DI(215) XOR DI(731) XOR DI(232) XOR DI(478) XOR DI(720) XOR DI(397) XOR DI(651) XOR DI(319) XOR DI(23) XOR DI(904) XOR DI(891) XOR DI(992) XOR DI(463) XOR DI(18) XOR DI(119) XOR DI(183) XOR DI(936) XOR DI(127) XOR DI(468) XOR DI(675) XOR DI(33) XOR DI(267) XOR DI(296) XOR DI(40) XOR DI(963) XOR DI(721) XOR DI(599) XOR DI(140) XOR DI(625) XOR DI(150) XOR DI(689) XOR DI(408) XOR DI(371) XOR DI(343) XOR DI(120) XOR DI(424) XOR DI(820) XOR DI(437) XOR DI(235) XOR DI(874) XOR DI(313) XOR DI(534) XOR DI(411) XOR DI(211) XOR DI(630) XOR DI(292) XOR DI(177) XOR DI(261) XOR DI(553) XOR DI(670) XOR DI(950) XOR DI(134) XOR DI(619) XOR DI(365) XOR DI(154) XOR DI(814) XOR DI(198) XOR DI(431) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(394) XOR DI(205) XOR DI(624) XOR DI(316) XOR DI(495) XOR DI(547) XOR DI(951) XOR DI(944) XOR DI(148) XOR DI(862) XOR DI(5) XOR DI(522) XOR DI(199) XOR DI(541) XOR DI(938) XOR DI(142) XOR DI(856) XOR DI(483) XOR DI(535) XOR DI(690) XOR DI(124) XOR DI(678) XOR DI(511) XOR DI(505) XOR DI(1017) XOR DI(1023);
   DO(9) <= DI(767) XOR DI(234) XOR DI(836) XOR DI(378) XOR DI(794) XOR DI(971) XOR DI(687) XOR DI(772) XOR DI(838) XOR DI(628) XOR DI(585) XOR DI(278) XOR DI(508) XOR DI(1009) XOR DI(860) XOR DI(828) XOR DI(91) XOR DI(662) XOR DI(218) XOR DI(602) XOR DI(26) XOR DI(104) XOR DI(961) XOR DI(242) XOR DI(817) XOR DI(51) XOR DI(757) XOR DI(77) XOR DI(560) XOR DI(677) XOR DI(784) XOR DI(470) XOR DI(578) XOR DI(280) XOR DI(161) XOR DI(363) XOR DI(392) XOR DI(646) XOR DI(596) XOR DI(3) XOR DI(20) XOR DI(71) XOR DI(778) XOR DI(908) XOR DI(996) XOR DI(441) XOR DI(893) XOR DI(382) XOR DI(588) XOR DI(798) XOR DI(634) XOR DI(376) XOR DI(638) XOR DI(490) XOR DI(451) XOR DI(187) XOR DI(653) XOR DI(1000) XOR DI(1012) XOR DI(576) XOR DI(577) XOR DI(435) XOR DI(844) XOR DI(785) XOR DI(915) XOR DI(95) XOR DI(693) XOR DI(112) XOR DI(594) XOR DI(55) XOR DI(622) XOR DI(176) XOR DI(96) XOR DI(471) XOR DI(902) XOR DI(520) XOR DI(966) XOR DI(289) XOR DI(877) XOR DI(272) XOR DI(716) XOR DI(876) XOR DI(597) XOR DI(455) XOR DI(60) XOR DI(311) XOR DI(812) XOR DI(98) XOR DI(656) XOR DI(606) XOR DI(389) XOR DI(931) XOR DI(346) XOR DI(843) XOR DI(1004) XOR DI(72) XOR DI(28) XOR DI(74) XOR DI(338) XOR DI(779) XOR DI(284) XOR DI(341) XOR DI(563) XOR DI(244) XOR DI(339) XOR DI(770) XOR DI(710) XOR DI(54) XOR DI(806) XOR DI(982) XOR DI(453) XOR DI(650) XOR DI(271) XOR DI(318) XOR DI(30) XOR DI(333) XOR DI(194) XOR DI(864) XOR DI(53) XOR DI(401) XOR DI(197) XOR DI(327) XOR DI(518) XOR DI(195) XOR DI(473) XOR DI(741) XOR DI(580) XOR DI(899) XOR DI(581) XOR DI(439) XOR DI(827) XOR DI(988) XOR DI(790) XOR DI(83) XOR DI(933) XOR DI(918) XOR DI(866) XOR DI(568) XOR DI(62) XOR DI(326) XOR DI(99) XOR DI(185) XOR DI(834) XOR DI(461) XOR DI(545) XOR DI(949) XOR DI(697) XOR DI(730) XOR DI(59) XOR DI(180) XOR DI(100) XOR DI(524) XOR DI(1) XOR DI(934) XOR DI(668) XOR DI(753) XOR DI(890) XOR DI(364) XOR DI(224) XOR DI(50) XOR DI(698) XOR DI(250) XOR DI(881) XOR DI(873) XOR DI(882) XOR DI(9) XOR DI(487) XOR DI(131) XOR DI(680) XOR DI(102) XOR DI(168) XOR DI(584) XOR DI(610) XOR DI(805) XOR DI(277) XOR DI(538) XOR DI(935) XOR DI(847) XOR DI(923) XOR DI(987) XOR DI(76) XOR DI(324) XOR DI(32) XOR DI(78) XOR DI(342) XOR DI(288) XOR DI(818) XOR DI(426) XOR DI(110) XOR DI(482) XOR DI(985) XOR DI(914) XOR DI(787) XOR DI(774) XOR DI(743) XOR DI(712) XOR DI(362) XOR DI(801) XOR DI(621) XOR DI(407) XOR DI(58) XOR DI(810) XOR DI(457) XOR DI(883) XOR DI(603) XOR DI(930) XOR DI(669) XOR DI(67) XOR DI(715) XOR DI(593) XOR DI(202) XOR DI(114) XOR DI(418) XOR DI(203) XOR DI(719) XOR DI(639) XOR DI(307) XOR DI(57) XOR DI(405) XOR DI(980) XOR DI(717) XOR DI(648) XOR DI(13) XOR DI(171) XOR DI(115) XOR DI(255) XOR DI(901) XOR DI(613) XOR DI(359) XOR DI(201) XOR DI(808) XOR DI(388) XOR DI(310) XOR DI(454) XOR DI(612) XOR DI(850) XOR DI(510) XOR DI(477) XOR DI(499) XOR DI(1005) XOR DI(575) XOR DI(999) XOR DI(775) XOR DI(279) XOR DI(867) XOR DI(706) XOR DI(587) XOR DI(88) XOR DI(379) XOR DI(336) XOR DI(994) XOR DI(329) XOR DI(854) XOR DI(571) XOR DI(978) XOR DI(89) XOR DI(49) XOR DI(170) XOR DI(90) XOR DI(924) XOR DI(574) XOR DI(925) XOR DI(837) XOR DI(68) XOR DI(975) XOR DI(764) XOR DI(191) XOR DI(840) XOR DI(561) XOR DI(968) XOR DI(965) XOR DI(181) XOR DI(830) XOR DI(958) XOR DI(955) XOR DI(637) XOR DI(579) XOR DI(703) XOR DI(122) XOR DI(448) XOR DI(162) XOR DI(220) XOR DI(647) XOR DI(65) XOR DI(632) XOR DI(4) XOR DI(909) XOR DI(979) XOR DI(841) XOR DI(106) XOR DI(685) XOR DI(367) XOR DI(997) XOR DI(420) XOR DI(530) XOR DI(383) XOR DI(173) XOR DI(497) XOR DI(589) XOR DI(260) XOR DI(976) XOR DI(713) XOR DI(265) XOR DI(188) XOR DI(132) XOR DI(759) XOR DI(766) XOR DI(436) XOR DI(299) XOR DI(755) XOR DI(724) XOR DI(458) XOR DI(172) XOR DI(230) XOR DI(623) XOR DI(358) XOR DI(374) XOR DI(704) XOR DI(123) XOR DI(665) XOR DI(750) XOR DI(887) XOR DI(746) XOR DI(282) XOR DI(533) XOR DI(221) XOR DI(614) XOR DI(737) XOR DI(238) XOR DI(728) XOR DI(813) XOR DI(888) XOR DI(726) XOR DI(657) XOR DI(15) XOR DI(249) XOR DI(504) XOR DI(493) XOR DI(70) XOR DI(852) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(546) XOR DI(137) XOR DI(686) XOR DI(711) XOR DI(642) XOR DI(14) XOR DI(895) XOR DI(174) XOR DI(666) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(616) XOR DI(334) XOR DI(811) XOR DI(865) XOR DI(304) XOR DI(283) XOR DI(544) XOR DI(661) XOR DI(941) XOR DI(356) XOR DI(145) XOR DI(189) XOR DI(196) XOR DI(615) XOR DI(853) XOR DI(532) XOR DI(929) XOR DI(502) XOR DI(1014) XOR DI(762) XOR DI(330) XOR DI(323) XOR DI(302) XOR DI(43) XOR DI(164) XOR DI(919) XOR DI(758) XOR DI(989) XOR DI(851) XOR DI(555) XOR DI(962) XOR DI(175) XOR DI(146) XOR DI(351) XOR DI(116) XOR DI(156) XOR DI(214) XOR DI(695) XOR DI(414) XOR DI(377) XOR DI(491) XOR DI(793) XOR DI(537) XOR DI(349) XOR DI(922) XOR DI(126) XOR DI(1007) XOR DI(430) XOR DI(452) XOR DI(826) XOR DI(210) XOR DI(744) XOR DI(421) XOR DI(740) XOR DI(276) XOR DI(215) XOR DI(241) XOR DI(807) XOR DI(627) XOR DI(880) XOR DI(651) XOR DI(243) XOR DI(319) XOR DI(498) XOR DI(64) XOR DI(23) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(891) XOR DI(992) XOR DI(217) XOR DI(463) XOR DI(705) XOR DI(8) XOR DI(18) XOR DI(393) XOR DI(298) XOR DI(655) XOR DI(350) XOR DI(183) XOR DI(936) XOR DI(507) XOR DI(127) XOR DI(296) XOR DI(40) XOR DI(825) XOR DI(404) XOR DI(963) XOR DI(599) XOR DI(956) XOR DI(150) XOR DI(208) XOR DI(689) XOR DI(829) XOR DI(900) XOR DI(408) XOR DI(424) XOR DI(809) XOR DI(820) XOR DI(509) XOR DI(270) XOR DI(209) XOR DI(235) XOR DI(645) XOR DI(313) XOR DI(17) XOR DI(411) XOR DI(986) XOR DI(723) XOR DI(400) XOR DI(12) XOR DI(275) XOR DI(322) XOR DI(649) XOR DI(113) XOR DI(177) XOR DI(261) XOR DI(553) XOR DI(957) XOR DI(950) XOR DI(163) XOR DI(134) XOR DI(619) XOR DI(365) XOR DI(337) XOR DI(814) XOR DI(198) XOR DI(431) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(11) XOR DI(394) XOR DI(205) XOR DI(316) XOR DI(456) XOR DI(547) XOR DI(944) XOR DI(702) XOR DI(618) XOR DI(375) XOR DI(489) XOR DI(541) XOR DI(938) XOR DI(142) XOR DI(856) XOR DI(529) XOR DI(684) XOR DI(678) XOR DI(517) XOR DI(505) XOR DI(1011) XOR DI(1023);
   DO(10) <= DI(768) XOR DI(833) XOR DI(86) XOR DI(834) XOR DI(466) XOR DI(148) XOR DI(999) XOR DI(772) XOR DI(235) XOR DI(837) XOR DI(559) XOR DI(587) XOR DI(301) XOR DI(379) XOR DI(795) XOR DI(49) XOR DI(972) XOR DI(688) XOR DI(773) XOR DI(217) XOR DI(873) XOR DI(839) XOR DI(629) XOR DI(25) XOR DI(682) XOR DI(586) XOR DI(943) XOR DI(424) XOR DI(279) XOR DI(689) XOR DI(509) XOR DI(1010) XOR DI(861) XOR DI(57) XOR DI(829) XOR DI(470) XOR DI(92) XOR DI(663) XOR DI(219) XOR DI(45) XOR DI(612) XOR DI(906) XOR DI(603) XOR DI(185) XOR DI(27) XOR DI(105) XOR DI(962) XOR DI(243) XOR DI(996) XOR DI(769) XOR DI(796) XOR DI(818) XOR DI(224) XOR DI(634) XOR DI(302) XOR DI(52) XOR DI(354) XOR DI(758) XOR DI(269) XOR DI(78) XOR DI(326) XOR DI(561) XOR DI(42) XOR DI(678) XOR DI(785) XOR DI(322) XOR DI(471) XOR DI(579) XOR DI(93) XOR DI(281) XOR DI(162) XOR DI(46) XOR DI(364) XOR DI(417) XOR DI(736) XOR DI(393) XOR DI(647) XOR DI(597) XOR DI(413) XOR DI(213) XOR DI(4) XOR DI(248) XOR DI(21) XOR DI(72) XOR DI(779) XOR DI(909) XOR DI(400) XOR DI(748) XOR DI(563) XOR DI(106) XOR DI(997) XOR DI(420) XOR DI(442) XOR DI(156) XOR DI(734) XOR DI(468) XOR DI(797) XOR DI(591) XOR DI(309) XOR DI(894) XOR DI(383) XOR DI(109) XOR DI(257) XOR DI(589) XOR DI(333) XOR DI(799) XOR DI(635) XOR DI(53) XOR DI(377) XOR DI(639) XOR DI(491) XOR DI(452) XOR DI(543) XOR DI(940) XOR DI(134) XOR DI(355) XOR DI(188) XOR DI(371) XOR DI(446) XOR DI(654) XOR DI(450) XOR DI(608) XOR DI(928) XOR DI(126) XOR DI(1001) XOR DI(1013) XOR DI(577) XOR DI(858) XOR DI(578) XOR DI(436) XOR DI(292) XOR DI(787) XOR DI(845) XOR DI(786) XOR DI(916) XOR DI(755) XOR DI(96) XOR DI(552) XOR DI(429) XOR DI(694) XOR DI(113) XOR DI(439) XOR DI(153) XOR DI(595) XOR DI(485) XOR DI(56) XOR DI(623) XOR DI(177) XOR DI(97) XOR DI(358) XOR DI(472) XOR DI(903) XOR DI(521) XOR DI(967) XOR DI(887) XOR DI(290) XOR DI(878) XOR DI(737) XOR DI(273) XOR DI(605) XOR DI(475) XOR DI(717) XOR DI(877) XOR DI(240) XOR DI(598) XOR DI(495) XOR DI(456) XOR DI(61) XOR DI(312) XOR DI(813) XOR DI(99) XOR DI(702) XOR DI(918) XOR DI(657) XOR DI(607) XOR DI(390) XOR DI(932) XOR DI(347) XOR DI(187) XOR DI(844) XOR DI(1005) XOR DI(30) XOR DI(73) XOR DI(29) XOR DI(75) XOR DI(339) XOR DI(780) XOR DI(822) XOR DI(285) XOR DI(342) XOR DI(564) XOR DI(897) XOR DI(482) XOR DI(245) XOR DI(961) XOR DI(340) XOR DI(913) XOR DI(771) XOR DI(798) XOR DI(711) XOR DI(404) XOR DI(55) XOR DI(807) XOR DI(983) XOR DI(454) XOR DI(880) XOR DI(651) XOR DI(272) XOR DI(319) XOR DI(927) XOR DI(31) XOR DI(522) XOR DI(334) XOR DI(800) XOR DI(195) XOR DI(428) XOR DI(226) XOR DI(865) XOR DI(636) XOR DI(304) XOR DI(8) XOR DI(54) XOR DI(402) XOR DI(104) XOR DI(544) XOR DI(898) XOR DI(941) XOR DI(356) XOR DI(198) XOR DI(328) XOR DI(519) XOR DI(196) XOR DI(513) XOR DI(441) XOR DI(929) XOR DI(474) XOR DI(675) XOR DI(514) XOR DI(1014) XOR DI(994) XOR DI(742) XOR DI(581) XOR DI(900) XOR DI(80) XOR DI(40) XOR DI(274) XOR DI(862) XOR DI(582) XOR DI(440) XOR DI(83) XOR DI(828) XOR DI(989) XOR DI(39) XOR DI(791) XOR DI(566) XOR DI(47) XOR DI(84) XOR DI(934) XOR DI(85) XOR DI(919) XOR DI(349) XOR DI(683) XOR DI(867) XOR DI(569) XOR DI(790) XOR DI(832) XOR DI(63) XOR DI(327) XOR DI(411) XOR DI(970) XOR DI(728) XOR DI(606) XOR DI(43) XOR DI(100) XOR DI(186) XOR DI(295) XOR DI(835) XOR DI(462) XOR DI(825) XOR DI(546) XOR DI(950) XOR DI(433) XOR DI(632) XOR DI(574) XOR DI(698) XOR DI(731) XOR DI(489) XOR DI(60) XOR DI(181) XOR DI(974) XOR DI(836) XOR DI(101) XOR DI(680) XOR DI(907) XOR DI(992) XOR DI(525) XOR DI(921) XOR DI(255) XOR DI(220) XOR DI(2) XOR DI(971) XOR DI(935) XOR DI(669) XOR DI(754) XOR DI(891) XOR DI(365) XOR DI(781) XOR DI(750) XOR DI(719) XOR DI(167) XOR DI(816) XOR DI(225) XOR DI(51) XOR DI(516) XOR DI(369) XOR DI(699) XOR DI(251) XOR DI(118) XOR DI(882) XOR DI(444) XOR DI(732) XOR DI(233) XOR DI(874) XOR DI(479) XOR DI(883) XOR DI(721) XOR DI(398) XOR DI(10) XOR DI(602) XOR DI(414) XOR DI(488) XOR DI(316) XOR DI(150) XOR DI(70) XOR DI(418) XOR DI(132) XOR DI(681) XOR DI(103) XOR DI(730) XOR DI(407) XOR DI(637) XOR DI(890) XOR DI(169) XOR DI(661) XOR DI(282) XOR DI(26) XOR DI(585) XOR DI(611) XOR DI(329) XOR DI(806) XOR DI(278) XOR DI(539) XOR DI(936) XOR DI(120) XOR DI(610) XOR DI(848) XOR DI(924) XOR DI(469) XOR DI(676) XOR DI(988) XOR DI(74) XOR DI(34) XOR DI(268) XOR DI(77) XOR DI(325) XOR DI(33) XOR DI(560) XOR DI(79) XOR DI(343) XOR DI(677) XOR DI(914) XOR DI(722) XOR DI(289) XOR DI(170) XOR DI(819) XOR DI(427) XOR DI(141) XOR DI(626) XOR DI(111) XOR DI(483) XOR DI(986) XOR DI(372) XOR DI(915) XOR DI(788) XOR DI(214) XOR DI(532) XOR DI(344) XOR DI(121) XOR DI(775) XOR DI(744) XOR DI(713) XOR DI(161) XOR DI(363) XOR DI(205) XOR DI(438) XOR DI(726) XOR DI(473) XOR DI(802) XOR DI(715) XOR DI(392) XOR DI(622) XOR DI(875) XOR DI(238) XOR DI(408) XOR DI(493) XOR DI(59) XOR DI(64) XOR DI(899) XOR DI(811) XOR DI(535) XOR DI(212) XOR DI(458) XOR DI(631) XOR DI(3) XOR DI(884) XOR DI(655) XOR DI(20) XOR DI(388) XOR DI(293) XOR DI(604) XOR DI(931) XOR DI(502) XOR DI(122) XOR DI(463) XOR DI(670) XOR DI(68) XOR DI(28) XOR DI(671) XOR DI(908) XOR DI(716) XOR DI(594) XOR DI(145) XOR DI(203) XOR DI(208) XOR DI(115) XOR DI(419) XOR DI(155) XOR DI(204) XOR DI(720) XOR DI(640) XOR DI(308) XOR DI(58) XOR DI(529) XOR DI(406) XOR DI(981) XOR DI(718) XOR DI(625) XOR DI(649) XOR DI(14) XOR DI(382) XOR DI(172) XOR DI(496) XOR DI(116) XOR DI(256) XOR DI(665) XOR DI(902) XOR DI(952) XOR DI(614) XOR DI(360) XOR DI(202) XOR DI(149) XOR DI(809) XOR DI(461) XOR DI(863) XOR DI(6) XOR DI(523) XOR DI(389) XOR DI(200) XOR DI(311) XOR DI(451) XOR DI(455) XOR DI(697) XOR DI(0) XOR DI(517) XOR DI(613) XOR DI(484) XOR DI(536) XOR DI(137) XOR DI(691) XOR DI(851) XOR DI(511) XOR DI(478) XOR DI(131) XOR DI(524) XOR DI(125) XOR DI(512) XOR DI(500) XOR DI(1006) XOR DI(1018);
   DO(11) <= DI(769) XOR DI(834) XOR DI(87) XOR DI(835) XOR DI(467) XOR DI(149) XOR DI(1000) XOR DI(773) XOR DI(236) XOR DI(838) XOR DI(560) XOR DI(588) XOR DI(302) XOR DI(380) XOR DI(796) XOR DI(50) XOR DI(973) XOR DI(689) XOR DI(774) XOR DI(218) XOR DI(874) XOR DI(840) XOR DI(630) XOR DI(26) XOR DI(683) XOR DI(587) XOR DI(944) XOR DI(425) XOR DI(280) XOR DI(690) XOR DI(510) XOR DI(1011) XOR DI(862) XOR DI(58) XOR DI(830) XOR DI(471) XOR DI(93) XOR DI(664) XOR DI(220) XOR DI(46) XOR DI(613) XOR DI(907) XOR DI(604) XOR DI(186) XOR DI(28) XOR DI(106) XOR DI(963) XOR DI(244) XOR DI(997) XOR DI(770) XOR DI(797) XOR DI(819) XOR DI(225) XOR DI(635) XOR DI(303) XOR DI(53) XOR DI(355) XOR DI(759) XOR DI(270) XOR DI(79) XOR DI(327) XOR DI(562) XOR DI(43) XOR DI(679) XOR DI(786) XOR DI(323) XOR DI(472) XOR DI(580) XOR DI(94) XOR DI(282) XOR DI(163) XOR DI(47) XOR DI(365) XOR DI(418) XOR DI(737) XOR DI(394) XOR DI(648) XOR DI(598) XOR DI(414) XOR DI(214) XOR DI(5) XOR DI(249) XOR DI(22) XOR DI(73) XOR DI(780) XOR DI(910) XOR DI(401) XOR DI(749) XOR DI(564) XOR DI(107) XOR DI(998) XOR DI(421) XOR DI(443) XOR DI(157) XOR DI(735) XOR DI(469) XOR DI(798) XOR DI(592) XOR DI(310) XOR DI(895) XOR DI(384) XOR DI(110) XOR DI(258) XOR DI(590) XOR DI(334) XOR DI(800) XOR DI(636) XOR DI(54) XOR DI(378) XOR DI(640) XOR DI(492) XOR DI(453) XOR DI(544) XOR DI(941) XOR DI(135) XOR DI(356) XOR DI(189) XOR DI(372) XOR DI(447) XOR DI(655) XOR DI(451) XOR DI(609) XOR DI(929) XOR DI(127) XOR DI(1002) XOR DI(1014) XOR DI(578) XOR DI(859) XOR DI(579) XOR DI(437) XOR DI(293) XOR DI(788) XOR DI(846) XOR DI(787) XOR DI(917) XOR DI(756) XOR DI(97) XOR DI(553) XOR DI(430) XOR DI(695) XOR DI(114) XOR DI(440) XOR DI(154) XOR DI(596) XOR DI(486) XOR DI(57) XOR DI(624) XOR DI(178) XOR DI(98) XOR DI(359) XOR DI(473) XOR DI(904) XOR DI(522) XOR DI(968) XOR DI(888) XOR DI(291) XOR DI(879) XOR DI(738) XOR DI(274) XOR DI(606) XOR DI(476) XOR DI(718) XOR DI(878) XOR DI(241) XOR DI(599) XOR DI(496) XOR DI(457) XOR DI(62) XOR DI(313) XOR DI(814) XOR DI(100) XOR DI(703) XOR DI(919) XOR DI(658) XOR DI(608) XOR DI(391) XOR DI(933) XOR DI(348) XOR DI(188) XOR DI(845) XOR DI(1006) XOR DI(31) XOR DI(74) XOR DI(30) XOR DI(76) XOR DI(340) XOR DI(781) XOR DI(823) XOR DI(286) XOR DI(343) XOR DI(565) XOR DI(898) XOR DI(483) XOR DI(246) XOR DI(962) XOR DI(341) XOR DI(914) XOR DI(772) XOR DI(799) XOR DI(712) XOR DI(405) XOR DI(56) XOR DI(808) XOR DI(984) XOR DI(455) XOR DI(881) XOR DI(652) XOR DI(273) XOR DI(320) XOR DI(928) XOR DI(32) XOR DI(523) XOR DI(335) XOR DI(801) XOR DI(196) XOR DI(429) XOR DI(227) XOR DI(866) XOR DI(637) XOR DI(305) XOR DI(9) XOR DI(55) XOR DI(403) XOR DI(105) XOR DI(545) XOR DI(899) XOR DI(942) XOR DI(357) XOR DI(199) XOR DI(329) XOR DI(520) XOR DI(197) XOR DI(514) XOR DI(442) XOR DI(930) XOR DI(475) XOR DI(676) XOR DI(515) XOR DI(1015) XOR DI(995) XOR DI(743) XOR DI(582) XOR DI(901) XOR DI(81) XOR DI(41) XOR DI(275) XOR DI(863) XOR DI(583) XOR DI(441) XOR DI(84) XOR DI(829) XOR DI(990) XOR DI(40) XOR DI(792) XOR DI(567) XOR DI(48) XOR DI(85) XOR DI(935) XOR DI(86) XOR DI(920) XOR DI(350) XOR DI(684) XOR DI(868) XOR DI(570) XOR DI(791) XOR DI(833) XOR DI(64) XOR DI(328) XOR DI(412) XOR DI(971) XOR DI(729) XOR DI(607) XOR DI(44) XOR DI(101) XOR DI(187) XOR DI(296) XOR DI(836) XOR DI(463) XOR DI(826) XOR DI(547) XOR DI(951) XOR DI(434) XOR DI(633) XOR DI(575) XOR DI(699) XOR DI(732) XOR DI(490) XOR DI(61) XOR DI(182) XOR DI(975) XOR DI(837) XOR DI(102) XOR DI(681) XOR DI(908) XOR DI(993) XOR DI(526) XOR DI(922) XOR DI(256) XOR DI(221) XOR DI(3) XOR DI(972) XOR DI(936) XOR DI(670) XOR DI(755) XOR DI(892) XOR DI(366) XOR DI(782) XOR DI(751) XOR DI(720) XOR DI(168) XOR DI(817) XOR DI(226) XOR DI(52) XOR DI(517) XOR DI(370) XOR DI(700) XOR DI(252) XOR DI(119) XOR DI(883) XOR DI(445) XOR DI(733) XOR DI(234) XOR DI(875) XOR DI(480) XOR DI(884) XOR DI(722) XOR DI(399) XOR DI(11) XOR DI(603) XOR DI(415) XOR DI(489) XOR DI(317) XOR DI(151) XOR DI(71) XOR DI(419) XOR DI(133) XOR DI(682) XOR DI(104) XOR DI(731) XOR DI(408) XOR DI(638) XOR DI(891) XOR DI(170) XOR DI(662) XOR DI(283) XOR DI(27) XOR DI(586) XOR DI(612) XOR DI(330) XOR DI(807) XOR DI(279) XOR DI(540) XOR DI(937) XOR DI(121) XOR DI(611) XOR DI(849) XOR DI(925) XOR DI(470) XOR DI(677) XOR DI(989) XOR DI(75) XOR DI(35) XOR DI(269) XOR DI(78) XOR DI(326) XOR DI(34) XOR DI(561) XOR DI(80) XOR DI(344) XOR DI(678) XOR DI(915) XOR DI(723) XOR DI(290) XOR DI(171) XOR DI(820) XOR DI(428) XOR DI(142) XOR DI(627) XOR DI(112) XOR DI(484) XOR DI(987) XOR DI(373) XOR DI(916) XOR DI(789) XOR DI(215) XOR DI(533) XOR DI(345) XOR DI(122) XOR DI(776) XOR DI(745) XOR DI(714) XOR DI(162) XOR DI(364) XOR DI(206) XOR DI(439) XOR DI(727) XOR DI(474) XOR DI(803) XOR DI(716) XOR DI(393) XOR DI(623) XOR DI(876) XOR DI(239) XOR DI(409) XOR DI(494) XOR DI(60) XOR DI(65) XOR DI(900) XOR DI(812) XOR DI(536) XOR DI(213) XOR DI(459) XOR DI(632) XOR DI(4) XOR DI(885) XOR DI(656) XOR DI(21) XOR DI(389) XOR DI(294) XOR DI(605) XOR DI(932) XOR DI(503) XOR DI(123) XOR DI(464) XOR DI(671) XOR DI(69) XOR DI(29) XOR DI(672) XOR DI(909) XOR DI(717) XOR DI(595) XOR DI(146) XOR DI(204) XOR DI(209) XOR DI(116) XOR DI(420) XOR DI(156) XOR DI(205) XOR DI(721) XOR DI(641) XOR DI(309) XOR DI(59) XOR DI(530) XOR DI(407) XOR DI(982) XOR DI(719) XOR DI(626) XOR DI(650) XOR DI(15) XOR DI(383) XOR DI(173) XOR DI(497) XOR DI(117) XOR DI(257) XOR DI(666) XOR DI(903) XOR DI(953) XOR DI(615) XOR DI(361) XOR DI(203) XOR DI(150) XOR DI(810) XOR DI(462) XOR DI(864) XOR DI(7) XOR DI(524) XOR DI(390) XOR DI(201) XOR DI(312) XOR DI(452) XOR DI(456) XOR DI(698) XOR DI(1) XOR DI(518) XOR DI(614) XOR DI(485) XOR DI(537) XOR DI(138) XOR DI(692) XOR DI(852) XOR DI(512) XOR DI(479) XOR DI(132) XOR DI(525) XOR DI(126) XOR DI(513) XOR DI(501) XOR DI(1007) XOR DI(1019);
   DO(12) <= DI(770) XOR DI(835) XOR DI(88) XOR DI(836) XOR DI(468) XOR DI(150) XOR DI(1001) XOR DI(774) XOR DI(237) XOR DI(839) XOR DI(561) XOR DI(589) XOR DI(303) XOR DI(381) XOR DI(797) XOR DI(51) XOR DI(974) XOR DI(690) XOR DI(775) XOR DI(219) XOR DI(875) XOR DI(841) XOR DI(631) XOR DI(27) XOR DI(684) XOR DI(588) XOR DI(945) XOR DI(426) XOR DI(281) XOR DI(691) XOR DI(511) XOR DI(1012) XOR DI(863) XOR DI(59) XOR DI(831) XOR DI(472) XOR DI(94) XOR DI(665) XOR DI(221) XOR DI(47) XOR DI(614) XOR DI(908) XOR DI(605) XOR DI(187) XOR DI(29) XOR DI(107) XOR DI(964) XOR DI(245) XOR DI(998) XOR DI(771) XOR DI(798) XOR DI(820) XOR DI(226) XOR DI(636) XOR DI(304) XOR DI(54) XOR DI(356) XOR DI(760) XOR DI(271) XOR DI(80) XOR DI(328) XOR DI(563) XOR DI(44) XOR DI(680) XOR DI(787) XOR DI(324) XOR DI(473) XOR DI(581) XOR DI(95) XOR DI(283) XOR DI(164) XOR DI(48) XOR DI(366) XOR DI(419) XOR DI(738) XOR DI(395) XOR DI(649) XOR DI(599) XOR DI(415) XOR DI(215) XOR DI(6) XOR DI(250) XOR DI(23) XOR DI(74) XOR DI(781) XOR DI(911) XOR DI(402) XOR DI(750) XOR DI(565) XOR DI(108) XOR DI(999) XOR DI(422) XOR DI(444) XOR DI(158) XOR DI(736) XOR DI(470) XOR DI(799) XOR DI(593) XOR DI(311) XOR DI(896) XOR DI(385) XOR DI(111) XOR DI(259) XOR DI(591) XOR DI(335) XOR DI(801) XOR DI(637) XOR DI(55) XOR DI(379) XOR DI(641) XOR DI(493) XOR DI(454) XOR DI(545) XOR DI(942) XOR DI(136) XOR DI(357) XOR DI(190) XOR DI(373) XOR DI(448) XOR DI(656) XOR DI(452) XOR DI(610) XOR DI(930) XOR DI(128) XOR DI(1003) XOR DI(1015) XOR DI(579) XOR DI(860) XOR DI(580) XOR DI(438) XOR DI(294) XOR DI(789) XOR DI(847) XOR DI(788) XOR DI(918) XOR DI(757) XOR DI(98) XOR DI(554) XOR DI(431) XOR DI(696) XOR DI(115) XOR DI(441) XOR DI(155) XOR DI(597) XOR DI(487) XOR DI(58) XOR DI(625) XOR DI(179) XOR DI(99) XOR DI(360) XOR DI(474) XOR DI(905) XOR DI(523) XOR DI(0) XOR DI(969) XOR DI(889) XOR DI(292) XOR DI(880) XOR DI(739) XOR DI(275) XOR DI(607) XOR DI(477) XOR DI(719) XOR DI(879) XOR DI(242) XOR DI(600) XOR DI(497) XOR DI(458) XOR DI(63) XOR DI(314) XOR DI(815) XOR DI(101) XOR DI(704) XOR DI(920) XOR DI(659) XOR DI(609) XOR DI(392) XOR DI(934) XOR DI(349) XOR DI(189) XOR DI(846) XOR DI(1007) XOR DI(32) XOR DI(75) XOR DI(31) XOR DI(77) XOR DI(341) XOR DI(782) XOR DI(824) XOR DI(287) XOR DI(344) XOR DI(566) XOR DI(899) XOR DI(484) XOR DI(247) XOR DI(963) XOR DI(342) XOR DI(915) XOR DI(773) XOR DI(800) XOR DI(713) XOR DI(406) XOR DI(57) XOR DI(809) XOR DI(985) XOR DI(456) XOR DI(882) XOR DI(653) XOR DI(274) XOR DI(321) XOR DI(929) XOR DI(33) XOR DI(524) XOR DI(336) XOR DI(802) XOR DI(197) XOR DI(430) XOR DI(228) XOR DI(867) XOR DI(638) XOR DI(306) XOR DI(10) XOR DI(56) XOR DI(404) XOR DI(106) XOR DI(546) XOR DI(900) XOR DI(943) XOR DI(358) XOR DI(200) XOR DI(330) XOR DI(521) XOR DI(198) XOR DI(515) XOR DI(443) XOR DI(931) XOR DI(476) XOR DI(677) XOR DI(516) XOR DI(1016) XOR DI(996) XOR DI(744) XOR DI(583) XOR DI(902) XOR DI(82) XOR DI(42) XOR DI(276) XOR DI(864) XOR DI(584) XOR DI(442) XOR DI(85) XOR DI(830) XOR DI(991) XOR DI(41) XOR DI(793) XOR DI(568) XOR DI(49) XOR DI(86) XOR DI(936) XOR DI(87) XOR DI(921) XOR DI(351) XOR DI(685) XOR DI(869) XOR DI(571) XOR DI(792) XOR DI(834) XOR DI(65) XOR DI(329) XOR DI(413) XOR DI(972) XOR DI(730) XOR DI(608) XOR DI(45) XOR DI(102) XOR DI(188) XOR DI(297) XOR DI(837) XOR DI(464) XOR DI(827) XOR DI(548) XOR DI(952) XOR DI(435) XOR DI(634) XOR DI(576) XOR DI(700) XOR DI(733) XOR DI(491) XOR DI(62) XOR DI(183) XOR DI(976) XOR DI(838) XOR DI(103) XOR DI(682) XOR DI(909) XOR DI(994) XOR DI(527) XOR DI(923) XOR DI(257) XOR DI(222) XOR DI(4) XOR DI(973) XOR DI(937) XOR DI(671) XOR DI(756) XOR DI(893) XOR DI(367) XOR DI(783) XOR DI(752) XOR DI(721) XOR DI(169) XOR DI(818) XOR DI(227) XOR DI(53) XOR DI(518) XOR DI(371) XOR DI(701) XOR DI(253) XOR DI(120) XOR DI(884) XOR DI(446) XOR DI(734) XOR DI(235) XOR DI(876) XOR DI(481) XOR DI(885) XOR DI(723) XOR DI(400) XOR DI(12) XOR DI(604) XOR DI(416) XOR DI(490) XOR DI(318) XOR DI(152) XOR DI(72) XOR DI(420) XOR DI(134) XOR DI(683) XOR DI(105) XOR DI(732) XOR DI(409) XOR DI(639) XOR DI(892) XOR DI(171) XOR DI(663) XOR DI(284) XOR DI(28) XOR DI(587) XOR DI(613) XOR DI(331) XOR DI(808) XOR DI(280) XOR DI(541) XOR DI(938) XOR DI(122) XOR DI(612) XOR DI(850) XOR DI(926) XOR DI(471) XOR DI(678) XOR DI(990) XOR DI(76) XOR DI(36) XOR DI(270) XOR DI(79) XOR DI(327) XOR DI(35) XOR DI(562) XOR DI(81) XOR DI(345) XOR DI(679) XOR DI(916) XOR DI(724) XOR DI(291) XOR DI(172) XOR DI(821) XOR DI(429) XOR DI(143) XOR DI(628) XOR DI(113) XOR DI(485) XOR DI(988) XOR DI(374) XOR DI(917) XOR DI(790) XOR DI(216) XOR DI(534) XOR DI(346) XOR DI(123) XOR DI(777) XOR DI(746) XOR DI(715) XOR DI(163) XOR DI(365) XOR DI(207) XOR DI(440) XOR DI(728) XOR DI(475) XOR DI(804) XOR DI(717) XOR DI(394) XOR DI(624) XOR DI(877) XOR DI(240) XOR DI(410) XOR DI(495) XOR DI(61) XOR DI(66) XOR DI(901) XOR DI(813) XOR DI(537) XOR DI(214) XOR DI(460) XOR DI(633) XOR DI(5) XOR DI(886) XOR DI(657) XOR DI(22) XOR DI(390) XOR DI(295) XOR DI(606) XOR DI(933) XOR DI(504) XOR DI(124) XOR DI(465) XOR DI(672) XOR DI(70) XOR DI(30) XOR DI(673) XOR DI(910) XOR DI(718) XOR DI(596) XOR DI(147) XOR DI(205) XOR DI(210) XOR DI(117) XOR DI(421) XOR DI(157) XOR DI(206) XOR DI(722) XOR DI(642) XOR DI(310) XOR DI(60) XOR DI(531) XOR DI(408) XOR DI(983) XOR DI(720) XOR DI(627) XOR DI(651) XOR DI(16) XOR DI(384) XOR DI(174) XOR DI(498) XOR DI(118) XOR DI(258) XOR DI(667) XOR DI(904) XOR DI(954) XOR DI(616) XOR DI(362) XOR DI(204) XOR DI(151) XOR DI(811) XOR DI(463) XOR DI(865) XOR DI(8) XOR DI(525) XOR DI(391) XOR DI(202) XOR DI(313) XOR DI(453) XOR DI(457) XOR DI(699) XOR DI(2) XOR DI(519) XOR DI(615) XOR DI(486) XOR DI(538) XOR DI(139) XOR DI(693) XOR DI(853) XOR DI(513) XOR DI(480) XOR DI(133) XOR DI(526) XOR DI(127) XOR DI(514) XOR DI(502) XOR DI(1008) XOR DI(1020);
   DO(13) <= DI(771) XOR DI(836) XOR DI(89) XOR DI(837) XOR DI(469) XOR DI(151) XOR DI(1002) XOR DI(775) XOR DI(238) XOR DI(840) XOR DI(562) XOR DI(590) XOR DI(304) XOR DI(382) XOR DI(798) XOR DI(52) XOR DI(975) XOR DI(691) XOR DI(776) XOR DI(220) XOR DI(876) XOR DI(842) XOR DI(632) XOR DI(28) XOR DI(685) XOR DI(589) XOR DI(946) XOR DI(427) XOR DI(282) XOR DI(692) XOR DI(512) XOR DI(1013) XOR DI(864) XOR DI(60) XOR DI(832) XOR DI(473) XOR DI(95) XOR DI(666) XOR DI(222) XOR DI(48) XOR DI(615) XOR DI(909) XOR DI(606) XOR DI(188) XOR DI(30) XOR DI(108) XOR DI(965) XOR DI(246) XOR DI(999) XOR DI(772) XOR DI(799) XOR DI(821) XOR DI(227) XOR DI(637) XOR DI(305) XOR DI(55) XOR DI(357) XOR DI(761) XOR DI(272) XOR DI(81) XOR DI(329) XOR DI(564) XOR DI(45) XOR DI(681) XOR DI(788) XOR DI(325) XOR DI(474) XOR DI(582) XOR DI(96) XOR DI(284) XOR DI(165) XOR DI(49) XOR DI(367) XOR DI(420) XOR DI(739) XOR DI(396) XOR DI(650) XOR DI(600) XOR DI(416) XOR DI(216) XOR DI(7) XOR DI(251) XOR DI(24) XOR DI(75) XOR DI(782) XOR DI(912) XOR DI(403) XOR DI(751) XOR DI(566) XOR DI(109) XOR DI(1000) XOR DI(423) XOR DI(445) XOR DI(159) XOR DI(737) XOR DI(471) XOR DI(800) XOR DI(594) XOR DI(312) XOR DI(897) XOR DI(386) XOR DI(112) XOR DI(260) XOR DI(592) XOR DI(336) XOR DI(802) XOR DI(638) XOR DI(56) XOR DI(380) XOR DI(642) XOR DI(494) XOR DI(455) XOR DI(546) XOR DI(943) XOR DI(137) XOR DI(358) XOR DI(191) XOR DI(374) XOR DI(449) XOR DI(657) XOR DI(453) XOR DI(611) XOR DI(931) XOR DI(129) XOR DI(1004) XOR DI(1016) XOR DI(580) XOR DI(861) XOR DI(581) XOR DI(439) XOR DI(295) XOR DI(790) XOR DI(848) XOR DI(789) XOR DI(919) XOR DI(758) XOR DI(99) XOR DI(555) XOR DI(432) XOR DI(697) XOR DI(116) XOR DI(442) XOR DI(156) XOR DI(598) XOR DI(488) XOR DI(59) XOR DI(626) XOR DI(180) XOR DI(100) XOR DI(361) XOR DI(475) XOR DI(906) XOR DI(524) XOR DI(1) XOR DI(970) XOR DI(890) XOR DI(293) XOR DI(881) XOR DI(740) XOR DI(276) XOR DI(608) XOR DI(478) XOR DI(720) XOR DI(880) XOR DI(243) XOR DI(601) XOR DI(498) XOR DI(459) XOR DI(64) XOR DI(315) XOR DI(816) XOR DI(102) XOR DI(705) XOR DI(921) XOR DI(660) XOR DI(610) XOR DI(393) XOR DI(935) XOR DI(350) XOR DI(190) XOR DI(847) XOR DI(1008) XOR DI(33) XOR DI(76) XOR DI(32) XOR DI(78) XOR DI(342) XOR DI(783) XOR DI(825) XOR DI(288) XOR DI(345) XOR DI(567) XOR DI(900) XOR DI(485) XOR DI(248) XOR DI(964) XOR DI(343) XOR DI(916) XOR DI(774) XOR DI(801) XOR DI(714) XOR DI(407) XOR DI(58) XOR DI(810) XOR DI(986) XOR DI(457) XOR DI(883) XOR DI(654) XOR DI(275) XOR DI(322) XOR DI(930) XOR DI(34) XOR DI(525) XOR DI(337) XOR DI(803) XOR DI(198) XOR DI(431) XOR DI(229) XOR DI(868) XOR DI(639) XOR DI(307) XOR DI(11) XOR DI(57) XOR DI(405) XOR DI(107) XOR DI(547) XOR DI(901) XOR DI(944) XOR DI(359) XOR DI(201) XOR DI(331) XOR DI(522) XOR DI(199) XOR DI(516) XOR DI(444) XOR DI(932) XOR DI(477) XOR DI(678) XOR DI(517) XOR DI(1017) XOR DI(997) XOR DI(745) XOR DI(584) XOR DI(903) XOR DI(83) XOR DI(43) XOR DI(277) XOR DI(865) XOR DI(585) XOR DI(443) XOR DI(86) XOR DI(831) XOR DI(992) XOR DI(42) XOR DI(794) XOR DI(569) XOR DI(50) XOR DI(87) XOR DI(937) XOR DI(88) XOR DI(922) XOR DI(352) XOR DI(686) XOR DI(870) XOR DI(572) XOR DI(793) XOR DI(835) XOR DI(66) XOR DI(330) XOR DI(414) XOR DI(973) XOR DI(731) XOR DI(609) XOR DI(46) XOR DI(103) XOR DI(189) XOR DI(298) XOR DI(838) XOR DI(465) XOR DI(828) XOR DI(549) XOR DI(953) XOR DI(436) XOR DI(635) XOR DI(577) XOR DI(701) XOR DI(734) XOR DI(492) XOR DI(63) XOR DI(184) XOR DI(977) XOR DI(839) XOR DI(104) XOR DI(683) XOR DI(910) XOR DI(995) XOR DI(528) XOR DI(924) XOR DI(258) XOR DI(223) XOR DI(5) XOR DI(974) XOR DI(938) XOR DI(672) XOR DI(757) XOR DI(894) XOR DI(368) XOR DI(784) XOR DI(753) XOR DI(722) XOR DI(170) XOR DI(819) XOR DI(228) XOR DI(54) XOR DI(519) XOR DI(372) XOR DI(702) XOR DI(254) XOR DI(121) XOR DI(885) XOR DI(447) XOR DI(735) XOR DI(236) XOR DI(877) XOR DI(482) XOR DI(886) XOR DI(724) XOR DI(401) XOR DI(13) XOR DI(605) XOR DI(417) XOR DI(491) XOR DI(319) XOR DI(153) XOR DI(73) XOR DI(421) XOR DI(135) XOR DI(684) XOR DI(106) XOR DI(733) XOR DI(410) XOR DI(640) XOR DI(893) XOR DI(172) XOR DI(664) XOR DI(285) XOR DI(29) XOR DI(588) XOR DI(614) XOR DI(332) XOR DI(809) XOR DI(281) XOR DI(542) XOR DI(939) XOR DI(123) XOR DI(613) XOR DI(851) XOR DI(927) XOR DI(472) XOR DI(679) XOR DI(991) XOR DI(77) XOR DI(37) XOR DI(271) XOR DI(80) XOR DI(328) XOR DI(36) XOR DI(563) XOR DI(82) XOR DI(346) XOR DI(680) XOR DI(917) XOR DI(725) XOR DI(292) XOR DI(173) XOR DI(822) XOR DI(430) XOR DI(144) XOR DI(629) XOR DI(114) XOR DI(486) XOR DI(989) XOR DI(375) XOR DI(918) XOR DI(791) XOR DI(217) XOR DI(535) XOR DI(347) XOR DI(124) XOR DI(778) XOR DI(747) XOR DI(716) XOR DI(164) XOR DI(366) XOR DI(208) XOR DI(441) XOR DI(729) XOR DI(476) XOR DI(805) XOR DI(718) XOR DI(395) XOR DI(625) XOR DI(878) XOR DI(241) XOR DI(411) XOR DI(496) XOR DI(62) XOR DI(67) XOR DI(902) XOR DI(814) XOR DI(538) XOR DI(215) XOR DI(461) XOR DI(634) XOR DI(6) XOR DI(887) XOR DI(658) XOR DI(23) XOR DI(391) XOR DI(296) XOR DI(607) XOR DI(934) XOR DI(505) XOR DI(125) XOR DI(466) XOR DI(673) XOR DI(71) XOR DI(31) XOR DI(674) XOR DI(911) XOR DI(719) XOR DI(597) XOR DI(148) XOR DI(206) XOR DI(211) XOR DI(118) XOR DI(422) XOR DI(158) XOR DI(207) XOR DI(723) XOR DI(643) XOR DI(311) XOR DI(61) XOR DI(532) XOR DI(409) XOR DI(984) XOR DI(721) XOR DI(628) XOR DI(0) XOR DI(652) XOR DI(17) XOR DI(385) XOR DI(175) XOR DI(499) XOR DI(119) XOR DI(259) XOR DI(668) XOR DI(905) XOR DI(955) XOR DI(617) XOR DI(363) XOR DI(205) XOR DI(152) XOR DI(812) XOR DI(464) XOR DI(866) XOR DI(9) XOR DI(526) XOR DI(392) XOR DI(203) XOR DI(314) XOR DI(454) XOR DI(458) XOR DI(700) XOR DI(3) XOR DI(520) XOR DI(616) XOR DI(487) XOR DI(539) XOR DI(140) XOR DI(694) XOR DI(854) XOR DI(514) XOR DI(481) XOR DI(134) XOR DI(527) XOR DI(128) XOR DI(515) XOR DI(503) XOR DI(1009) XOR DI(1021);
   DO(14) <= DI(772) XOR DI(837) XOR DI(90) XOR DI(838) XOR DI(470) XOR DI(152) XOR DI(1003) XOR DI(776) XOR DI(239) XOR DI(841) XOR DI(563) XOR DI(591) XOR DI(305) XOR DI(383) XOR DI(799) XOR DI(53) XOR DI(976) XOR DI(692) XOR DI(777) XOR DI(221) XOR DI(877) XOR DI(843) XOR DI(633) XOR DI(29) XOR DI(686) XOR DI(590) XOR DI(947) XOR DI(428) XOR DI(283) XOR DI(693) XOR DI(513) XOR DI(1014) XOR DI(865) XOR DI(61) XOR DI(833) XOR DI(474) XOR DI(96) XOR DI(667) XOR DI(223) XOR DI(49) XOR DI(616) XOR DI(910) XOR DI(607) XOR DI(189) XOR DI(31) XOR DI(109) XOR DI(966) XOR DI(247) XOR DI(1000) XOR DI(773) XOR DI(800) XOR DI(822) XOR DI(228) XOR DI(638) XOR DI(306) XOR DI(56) XOR DI(358) XOR DI(762) XOR DI(273) XOR DI(82) XOR DI(330) XOR DI(565) XOR DI(46) XOR DI(682) XOR DI(789) XOR DI(326) XOR DI(475) XOR DI(583) XOR DI(97) XOR DI(285) XOR DI(166) XOR DI(50) XOR DI(368) XOR DI(421) XOR DI(740) XOR DI(397) XOR DI(651) XOR DI(601) XOR DI(417) XOR DI(217) XOR DI(8) XOR DI(252) XOR DI(25) XOR DI(76) XOR DI(783) XOR DI(913) XOR DI(404) XOR DI(752) XOR DI(567) XOR DI(110) XOR DI(1001) XOR DI(424) XOR DI(446) XOR DI(160) XOR DI(738) XOR DI(472) XOR DI(801) XOR DI(595) XOR DI(313) XOR DI(898) XOR DI(387) XOR DI(113) XOR DI(261) XOR DI(593) XOR DI(337) XOR DI(803) XOR DI(639) XOR DI(57) XOR DI(381) XOR DI(643) XOR DI(495) XOR DI(456) XOR DI(547) XOR DI(944) XOR DI(138) XOR DI(359) XOR DI(192) XOR DI(375) XOR DI(450) XOR DI(658) XOR DI(454) XOR DI(612) XOR DI(932) XOR DI(130) XOR DI(1005) XOR DI(1017) XOR DI(581) XOR DI(862) XOR DI(582) XOR DI(440) XOR DI(296) XOR DI(791) XOR DI(849) XOR DI(790) XOR DI(920) XOR DI(759) XOR DI(100) XOR DI(556) XOR DI(433) XOR DI(698) XOR DI(117) XOR DI(443) XOR DI(157) XOR DI(599) XOR DI(489) XOR DI(60) XOR DI(627) XOR DI(181) XOR DI(101) XOR DI(362) XOR DI(476) XOR DI(907) XOR DI(525) XOR DI(2) XOR DI(971) XOR DI(891) XOR DI(294) XOR DI(882) XOR DI(741) XOR DI(277) XOR DI(609) XOR DI(479) XOR DI(721) XOR DI(881) XOR DI(244) XOR DI(602) XOR DI(499) XOR DI(460) XOR DI(65) XOR DI(316) XOR DI(817) XOR DI(103) XOR DI(706) XOR DI(922) XOR DI(661) XOR DI(611) XOR DI(394) XOR DI(936) XOR DI(351) XOR DI(191) XOR DI(848) XOR DI(1009) XOR DI(34) XOR DI(77) XOR DI(33) XOR DI(79) XOR DI(343) XOR DI(784) XOR DI(826) XOR DI(289) XOR DI(346) XOR DI(568) XOR DI(901) XOR DI(486) XOR DI(249) XOR DI(965) XOR DI(344) XOR DI(917) XOR DI(775) XOR DI(802) XOR DI(715) XOR DI(408) XOR DI(59) XOR DI(811) XOR DI(987) XOR DI(458) XOR DI(884) XOR DI(655) XOR DI(276) XOR DI(323) XOR DI(931) XOR DI(35) XOR DI(526) XOR DI(338) XOR DI(804) XOR DI(199) XOR DI(432) XOR DI(230) XOR DI(869) XOR DI(640) XOR DI(308) XOR DI(12) XOR DI(58) XOR DI(406) XOR DI(108) XOR DI(548) XOR DI(902) XOR DI(945) XOR DI(360) XOR DI(202) XOR DI(332) XOR DI(523) XOR DI(200) XOR DI(0) XOR DI(517) XOR DI(445) XOR DI(933) XOR DI(478) XOR DI(679) XOR DI(518) XOR DI(1018) XOR DI(998) XOR DI(746) XOR DI(585) XOR DI(904) XOR DI(84) XOR DI(44) XOR DI(278) XOR DI(866) XOR DI(586) XOR DI(444) XOR DI(87) XOR DI(832) XOR DI(993) XOR DI(43) XOR DI(795) XOR DI(570) XOR DI(51) XOR DI(88) XOR DI(938) XOR DI(89) XOR DI(923) XOR DI(353) XOR DI(687) XOR DI(871) XOR DI(573) XOR DI(794) XOR DI(836) XOR DI(67) XOR DI(331) XOR DI(415) XOR DI(974) XOR DI(732) XOR DI(610) XOR DI(47) XOR DI(104) XOR DI(190) XOR DI(299) XOR DI(839) XOR DI(466) XOR DI(829) XOR DI(550) XOR DI(954) XOR DI(437) XOR DI(636) XOR DI(578) XOR DI(702) XOR DI(735) XOR DI(493) XOR DI(64) XOR DI(185) XOR DI(978) XOR DI(840) XOR DI(105) XOR DI(684) XOR DI(911) XOR DI(996) XOR DI(529) XOR DI(925) XOR DI(259) XOR DI(224) XOR DI(6) XOR DI(975) XOR DI(939) XOR DI(673) XOR DI(758) XOR DI(895) XOR DI(369) XOR DI(785) XOR DI(754) XOR DI(723) XOR DI(171) XOR DI(820) XOR DI(229) XOR DI(55) XOR DI(520) XOR DI(373) XOR DI(703) XOR DI(255) XOR DI(122) XOR DI(886) XOR DI(448) XOR DI(736) XOR DI(237) XOR DI(878) XOR DI(483) XOR DI(887) XOR DI(725) XOR DI(402) XOR DI(14) XOR DI(606) XOR DI(418) XOR DI(492) XOR DI(320) XOR DI(154) XOR DI(74) XOR DI(422) XOR DI(136) XOR DI(685) XOR DI(107) XOR DI(734) XOR DI(411) XOR DI(641) XOR DI(894) XOR DI(173) XOR DI(665) XOR DI(286) XOR DI(30) XOR DI(589) XOR DI(615) XOR DI(333) XOR DI(810) XOR DI(282) XOR DI(543) XOR DI(940) XOR DI(124) XOR DI(614) XOR DI(852) XOR DI(928) XOR DI(473) XOR DI(680) XOR DI(992) XOR DI(78) XOR DI(38) XOR DI(272) XOR DI(81) XOR DI(329) XOR DI(37) XOR DI(564) XOR DI(83) XOR DI(347) XOR DI(681) XOR DI(918) XOR DI(726) XOR DI(293) XOR DI(174) XOR DI(823) XOR DI(431) XOR DI(145) XOR DI(630) XOR DI(115) XOR DI(487) XOR DI(990) XOR DI(376) XOR DI(919) XOR DI(792) XOR DI(218) XOR DI(536) XOR DI(348) XOR DI(125) XOR DI(779) XOR DI(748) XOR DI(717) XOR DI(165) XOR DI(367) XOR DI(209) XOR DI(442) XOR DI(730) XOR DI(477) XOR DI(806) XOR DI(719) XOR DI(396) XOR DI(626) XOR DI(879) XOR DI(242) XOR DI(412) XOR DI(497) XOR DI(63) XOR DI(68) XOR DI(903) XOR DI(815) XOR DI(539) XOR DI(216) XOR DI(462) XOR DI(635) XOR DI(7) XOR DI(888) XOR DI(659) XOR DI(24) XOR DI(392) XOR DI(297) XOR DI(608) XOR DI(935) XOR DI(506) XOR DI(126) XOR DI(467) XOR DI(674) XOR DI(72) XOR DI(32) XOR DI(675) XOR DI(912) XOR DI(720) XOR DI(598) XOR DI(149) XOR DI(207) XOR DI(212) XOR DI(119) XOR DI(423) XOR DI(159) XOR DI(208) XOR DI(724) XOR DI(644) XOR DI(312) XOR DI(62) XOR DI(533) XOR DI(410) XOR DI(985) XOR DI(722) XOR DI(629) XOR DI(1) XOR DI(653) XOR DI(18) XOR DI(386) XOR DI(176) XOR DI(500) XOR DI(120) XOR DI(260) XOR DI(669) XOR DI(906) XOR DI(956) XOR DI(618) XOR DI(364) XOR DI(206) XOR DI(153) XOR DI(813) XOR DI(465) XOR DI(867) XOR DI(10) XOR DI(527) XOR DI(393) XOR DI(204) XOR DI(315) XOR DI(455) XOR DI(459) XOR DI(701) XOR DI(4) XOR DI(521) XOR DI(617) XOR DI(488) XOR DI(540) XOR DI(141) XOR DI(695) XOR DI(855) XOR DI(515) XOR DI(482) XOR DI(135) XOR DI(528) XOR DI(129) XOR DI(516) XOR DI(504) XOR DI(1010) XOR DI(1022);
   DO(15) <= DI(773) XOR DI(838) XOR DI(91) XOR DI(839) XOR DI(471) XOR DI(153) XOR DI(1004) XOR DI(777) XOR DI(240) XOR DI(842) XOR DI(564) XOR DI(592) XOR DI(306) XOR DI(384) XOR DI(800) XOR DI(54) XOR DI(977) XOR DI(693) XOR DI(778) XOR DI(222) XOR DI(878) XOR DI(844) XOR DI(634) XOR DI(30) XOR DI(687) XOR DI(591) XOR DI(948) XOR DI(429) XOR DI(284) XOR DI(694) XOR DI(514) XOR DI(1015) XOR DI(866) XOR DI(62) XOR DI(834) XOR DI(475) XOR DI(97) XOR DI(668) XOR DI(224) XOR DI(50) XOR DI(617) XOR DI(911) XOR DI(608) XOR DI(190) XOR DI(32) XOR DI(110) XOR DI(967) XOR DI(248) XOR DI(1001) XOR DI(774) XOR DI(801) XOR DI(823) XOR DI(229) XOR DI(639) XOR DI(307) XOR DI(57) XOR DI(359) XOR DI(763) XOR DI(274) XOR DI(83) XOR DI(331) XOR DI(566) XOR DI(47) XOR DI(683) XOR DI(790) XOR DI(327) XOR DI(476) XOR DI(584) XOR DI(98) XOR DI(286) XOR DI(167) XOR DI(51) XOR DI(369) XOR DI(422) XOR DI(741) XOR DI(398) XOR DI(652) XOR DI(602) XOR DI(418) XOR DI(218) XOR DI(9) XOR DI(253) XOR DI(26) XOR DI(77) XOR DI(784) XOR DI(914) XOR DI(405) XOR DI(753) XOR DI(568) XOR DI(111) XOR DI(1002) XOR DI(425) XOR DI(447) XOR DI(161) XOR DI(739) XOR DI(473) XOR DI(802) XOR DI(596) XOR DI(314) XOR DI(899) XOR DI(388) XOR DI(114) XOR DI(262) XOR DI(594) XOR DI(338) XOR DI(804) XOR DI(640) XOR DI(58) XOR DI(382) XOR DI(644) XOR DI(496) XOR DI(457) XOR DI(548) XOR DI(945) XOR DI(139) XOR DI(360) XOR DI(193) XOR DI(376) XOR DI(451) XOR DI(659) XOR DI(455) XOR DI(613) XOR DI(933) XOR DI(131) XOR DI(1006) XOR DI(1018) XOR DI(582) XOR DI(863) XOR DI(583) XOR DI(441) XOR DI(297) XOR DI(792) XOR DI(850) XOR DI(791) XOR DI(921) XOR DI(760) XOR DI(101) XOR DI(557) XOR DI(434) XOR DI(699) XOR DI(118) XOR DI(444) XOR DI(158) XOR DI(600) XOR DI(490) XOR DI(61) XOR DI(628) XOR DI(0) XOR DI(182) XOR DI(102) XOR DI(363) XOR DI(477) XOR DI(908) XOR DI(526) XOR DI(3) XOR DI(972) XOR DI(892) XOR DI(295) XOR DI(883) XOR DI(742) XOR DI(278) XOR DI(610) XOR DI(480) XOR DI(722) XOR DI(882) XOR DI(245) XOR DI(603) XOR DI(500) XOR DI(461) XOR DI(66) XOR DI(317) XOR DI(818) XOR DI(104) XOR DI(707) XOR DI(923) XOR DI(662) XOR DI(612) XOR DI(395) XOR DI(937) XOR DI(352) XOR DI(192) XOR DI(849) XOR DI(1010) XOR DI(35) XOR DI(78) XOR DI(34) XOR DI(80) XOR DI(344) XOR DI(785) XOR DI(827) XOR DI(290) XOR DI(347) XOR DI(569) XOR DI(902) XOR DI(487) XOR DI(250) XOR DI(966) XOR DI(345) XOR DI(918) XOR DI(776) XOR DI(803) XOR DI(716) XOR DI(409) XOR DI(60) XOR DI(812) XOR DI(988) XOR DI(459) XOR DI(885) XOR DI(656) XOR DI(277) XOR DI(324) XOR DI(932) XOR DI(36) XOR DI(527) XOR DI(339) XOR DI(805) XOR DI(200) XOR DI(433) XOR DI(231) XOR DI(870) XOR DI(641) XOR DI(309) XOR DI(13) XOR DI(59) XOR DI(407) XOR DI(109) XOR DI(549) XOR DI(903) XOR DI(946) XOR DI(361) XOR DI(203) XOR DI(333) XOR DI(524) XOR DI(201) XOR DI(1) XOR DI(518) XOR DI(446) XOR DI(934) XOR DI(479) XOR DI(680) XOR DI(519) XOR DI(1019) XOR DI(999) XOR DI(747) XOR DI(586) XOR DI(905) XOR DI(85) XOR DI(45) XOR DI(279) XOR DI(867) XOR DI(587) XOR DI(445) XOR DI(88) XOR DI(833) XOR DI(994) XOR DI(44) XOR DI(796) XOR DI(571) XOR DI(52) XOR DI(89) XOR DI(939) XOR DI(90) XOR DI(924) XOR DI(354) XOR DI(688) XOR DI(872) XOR DI(574) XOR DI(795) XOR DI(837) XOR DI(68) XOR DI(332) XOR DI(416) XOR DI(975) XOR DI(733) XOR DI(611) XOR DI(48) XOR DI(105) XOR DI(191) XOR DI(300) XOR DI(840) XOR DI(467) XOR DI(830) XOR DI(551) XOR DI(955) XOR DI(438) XOR DI(637) XOR DI(579) XOR DI(703) XOR DI(736) XOR DI(494) XOR DI(65) XOR DI(186) XOR DI(979) XOR DI(841) XOR DI(106) XOR DI(685) XOR DI(912) XOR DI(997) XOR DI(530) XOR DI(926) XOR DI(260) XOR DI(225) XOR DI(7) XOR DI(976) XOR DI(940) XOR DI(674) XOR DI(759) XOR DI(896) XOR DI(370) XOR DI(786) XOR DI(755) XOR DI(724) XOR DI(172) XOR DI(821) XOR DI(230) XOR DI(56) XOR DI(521) XOR DI(374) XOR DI(704) XOR DI(256) XOR DI(123) XOR DI(887) XOR DI(449) XOR DI(737) XOR DI(238) XOR DI(879) XOR DI(484) XOR DI(888) XOR DI(726) XOR DI(403) XOR DI(15) XOR DI(607) XOR DI(419) XOR DI(493) XOR DI(321) XOR DI(155) XOR DI(75) XOR DI(423) XOR DI(137) XOR DI(686) XOR DI(108) XOR DI(735) XOR DI(412) XOR DI(642) XOR DI(895) XOR DI(174) XOR DI(666) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(616) XOR DI(334) XOR DI(811) XOR DI(283) XOR DI(544) XOR DI(941) XOR DI(125) XOR DI(615) XOR DI(853) XOR DI(929) XOR DI(474) XOR DI(681) XOR DI(993) XOR DI(79) XOR DI(39) XOR DI(273) XOR DI(82) XOR DI(330) XOR DI(38) XOR DI(565) XOR DI(84) XOR DI(348) XOR DI(682) XOR DI(919) XOR DI(727) XOR DI(294) XOR DI(175) XOR DI(824) XOR DI(432) XOR DI(146) XOR DI(631) XOR DI(116) XOR DI(488) XOR DI(991) XOR DI(377) XOR DI(920) XOR DI(793) XOR DI(219) XOR DI(537) XOR DI(349) XOR DI(126) XOR DI(780) XOR DI(749) XOR DI(718) XOR DI(166) XOR DI(368) XOR DI(210) XOR DI(443) XOR DI(731) XOR DI(478) XOR DI(807) XOR DI(720) XOR DI(397) XOR DI(627) XOR DI(880) XOR DI(243) XOR DI(413) XOR DI(498) XOR DI(64) XOR DI(69) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(217) XOR DI(463) XOR DI(636) XOR DI(8) XOR DI(889) XOR DI(660) XOR DI(25) XOR DI(393) XOR DI(298) XOR DI(609) XOR DI(936) XOR DI(507) XOR DI(127) XOR DI(468) XOR DI(675) XOR DI(73) XOR DI(33) XOR DI(676) XOR DI(913) XOR DI(721) XOR DI(599) XOR DI(150) XOR DI(208) XOR DI(213) XOR DI(120) XOR DI(424) XOR DI(160) XOR DI(209) XOR DI(725) XOR DI(645) XOR DI(313) XOR DI(63) XOR DI(534) XOR DI(411) XOR DI(986) XOR DI(723) XOR DI(630) XOR DI(2) XOR DI(654) XOR DI(19) XOR DI(387) XOR DI(177) XOR DI(501) XOR DI(121) XOR DI(261) XOR DI(670) XOR DI(907) XOR DI(957) XOR DI(619) XOR DI(365) XOR DI(207) XOR DI(154) XOR DI(814) XOR DI(466) XOR DI(868) XOR DI(11) XOR DI(528) XOR DI(394) XOR DI(205) XOR DI(316) XOR DI(456) XOR DI(460) XOR DI(702) XOR DI(5) XOR DI(522) XOR DI(618) XOR DI(489) XOR DI(541) XOR DI(142) XOR DI(696) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(136) XOR DI(529) XOR DI(130) XOR DI(517) XOR DI(505) XOR DI(1011) XOR DI(1023);
   DO(16) <= DI(774) XOR DI(839) XOR DI(50) XOR DI(636) XOR DI(356) XOR DI(92) XOR DI(337) XOR DI(840) XOR DI(769) XOR DI(590) XOR DI(798) XOR DI(302) XOR DI(472) XOR DI(93) XOR DI(563) XOR DI(154) XOR DI(359) XOR DI(1005) XOR DI(778) XOR DI(248) XOR DI(241) XOR DI(911) XOR DI(843) XOR DI(565) XOR DI(999) XOR DI(224) XOR DI(712) XOR DI(593) XOR DI(307) XOR DI(385) XOR DI(928) XOR DI(259) XOR DI(801) XOR DI(866) XOR DI(55) XOR DI(978) XOR DI(357) XOR DI(190) XOR DI(1015) XOR DI(898) XOR DI(694) XOR DI(779) XOR DI(814) XOR DI(223) XOR DI(879) XOR DI(845) XOR DI(635) XOR DI(189) XOR DI(31) XOR DI(688) XOR DI(800) XOR DI(929) XOR DI(592) XOR DI(949) XOR DI(197) XOR DI(430) XOR DI(979) XOR DI(285) XOR DI(943) XOR DI(358) XOR DI(695) XOR DI(855) XOR DI(515) XOR DI(482) XOR DI(1016) XOR DI(303) XOR DI(47) XOR DI(867) XOR DI(63) XOR DI(835) XOR DI(963) XOR DI(574) XOR DI(696) XOR DI(476) XOR DI(98) XOR DI(669) XOR DI(431) XOR DI(225) XOR DI(51) XOR DI(618) XOR DI(516) XOR DI(912) XOR DI(422) XOR DI(609) XOR DI(242) XOR DI(706) XOR DI(282) XOR DI(191) XOR DI(268) XOR DI(33) XOR DI(560) XOR DI(111) XOR DI(690) XOR DI(968) XOR DI(249) XOR DI(1002) XOR DI(775) XOR DI(438) XOR DI(473) XOR DI(802) XOR DI(392) XOR DI(18) XOR DI(899) XOR DI(323) XOR DI(164) XOR DI(135) XOR DI(824) XOR DI(338) XOR DI(199) XOR DI(230) XOR DI(640) XOR DI(308) XOR DI(58) XOR DI(625) XOR DI(382) XOR DI(496) XOR DI(665) XOR DI(945) XOR DI(360) XOR DI(451) XOR DI(125) XOR DI(1018) XOR DI(764) XOR DI(275) XOR DI(863) XOR DI(441) XOR DI(84) XOR DI(332) XOR DI(304) XOR DI(567) XOR DI(974) XOR DI(554) XOR DI(48) XOR DI(684) XOR DI(791) XOR DI(833) XOR DI(328) XOR DI(971) XOR DI(729) XOR DI(44) XOR DI(836) XOR DI(964) XOR DI(961) XOR DI(547) XOR DI(951) XOR DI(148) XOR DI(0) XOR DI(182) XOR DI(477) XOR DI(993) XOR DI(493) XOR DI(585) XOR DI(221) XOR DI(709) XOR DI(99) XOR DI(184) XOR DI(432) XOR DI(287) XOR DI(168) XOR DI(52) XOR DI(370) XOR DI(423) XOR DI(742) XOR DI(875) XOR DI(399) XOR DI(653) XOR DI(603) XOR DI(415) XOR DI(25) XOR DI(71) XOR DI(419) XOR DI(767) XOR DI(104) XOR DI(219) XOR DI(707) XOR DI(10) XOR DI(254) XOR DI(283) XOR DI(27) XOR DI(330) XOR DI(470) XOR DI(269) XOR DI(78) XOR DI(344) XOR DI(785) XOR DI(915) XOR DI(406) XOR DI(754) XOR DI(569) XOR DI(112) XOR DI(691) XOR DI(969) XOR DI(250) XOR DI(215) XOR DI(533) XOR DI(918) XOR DI(1003) XOR DI(426) XOR DI(776) XOR DI(745) XOR DI(714) XOR DI(448) XOR DI(162) XOR DI(740) XOR DI(474) XOR DI(803) XOR DI(597) XOR DI(315) XOR DI(19) XOR DI(900) XOR DI(536) XOR DI(887) XOR DI(656) XOR DI(277) XOR DI(389) XOR DI(324) XOR DI(115) XOR DI(605) XOR DI(503) XOR DI(263) XOR DI(292) XOR DI(595) XOR DI(165) XOR DI(339) XOR DI(805) XOR DI(816) XOR DI(505) XOR DI(200) XOR DI(266) XOR DI(641) XOR DI(233) XOR DI(309) XOR DI(13) XOR DI(59) XOR DI(626) XOR DI(650) XOR DI(271) XOR DI(383) XOR DI(645) XOR DI(497) XOR DI(458) XOR DI(549) XOR DI(666) XOR DI(946) XOR DI(140) XOR DI(361) XOR DI(150) XOR DI(194) XOR DI(524) XOR DI(377) XOR DI(452) XOR DI(660) XOR DI(456) XOR DI(614) XOR DI(934) XOR DI(852) XOR DI(132) XOR DI(680) XOR DI(1007) XOR DI(1019) XOR DI(996) XOR DI(583) XOR DI(765) XOR DI(772) XOR DI(42) XOR DI(276) XOR DI(864) XOR DI(584) XOR DI(442) XOR DI(298) XOR DI(376) XOR DI(830) XOR DI(326) XOR DI(41) XOR DI(793) XOR DI(305) XOR DI(851) XOR DI(351) XOR DI(685) XOR DI(792) XOR DI(922) XOR DI(329) XOR DI(761) XOR DI(730) XOR DI(102) XOR DI(297) XOR DI(558) XOR DI(751) XOR DI(827) XOR DI(548) XOR DI(952) XOR DI(435) XOR DI(149) XOR DI(634) XOR DI(354) XOR DI(576) XOR DI(700) XOR DI(119) XOR DI(445) XOR DI(159) XOR DI(217) XOR DI(601) XOR DI(236) XOR DI(491) XOR DI(62) XOR DI(629) XOR DI(1) XOR DI(183) XOR DI(103) XOR DI(364) XOR DI(478) XOR DI(909) XOR DI(527) XOR DI(380) XOR DI(170) XOR DI(923) XOR DI(222) XOR DI(300) XOR DI(4) XOR DI(973) XOR DI(352) XOR DI(185) XOR DI(763) XOR DI(893) XOR DI(296) XOR DI(559) XOR DI(213) XOR DI(120) XOR DI(662) XOR DI(747) XOR DI(884) XOR DI(743) XOR DI(279) XOR DI(611) XOR DI(437) XOR DI(481) XOR DI(810) XOR DI(723) XOR DI(400) XOR DI(883) XOR DI(246) XOR DI(604) XOR DI(501) XOR DI(462) XOR DI(67) XOR DI(318) XOR DI(907) XOR DI(819) XOR DI(957) XOR DI(543) XOR DI(134) XOR DI(105) XOR DI(409) XOR DI(466) XOR DI(708) XOR DI(892) XOR DI(171) XOR DI(924) XOR DI(663) XOR DI(255) XOR DI(28) XOR DI(613) XOR DI(396) XOR DI(862) XOR DI(658) XOR DI(938) XOR DI(353) XOR DI(193) XOR DI(939) XOR DI(850) XOR DI(510) XOR DI(926) XOR DI(1011) XOR DI(990) XOR DI(759) XOR DI(36) XOR DI(858) XOR DI(79) XOR DI(320) XOR DI(35) XOR DI(562) XOR DI(43) XOR DI(81) XOR DI(345) XOR DI(679) XOR DI(786) XOR DI(828) XOR DI(407) XOR DI(966) XOR DI(755) XOR DI(602) XOR DI(291) XOR DI(959) XOR DI(821) XOR DI(429) XOR DI(348) XOR DI(570) XOR DI(153) XOR DI(970) XOR DI(832) XOR DI(903) XOR DI(411) XOR DI(488) XOR DI(790) XOR DI(251) XOR DI(216) XOR DI(967) XOR DI(534) XOR DI(346) XOR DI(919) XOR DI(123) XOR DI(777) XOR DI(715) XOR DI(449) XOR DI(163) XOR DI(823) XOR DI(512) XOR DI(114) XOR DI(741) XOR DI(418) XOR DI(212) XOR DI(238) XOR DI(804) XOR DI(717) XOR DI(624) XOR DI(648) XOR DI(240) XOR DI(316) XOR DI(410) XOR DI(61) XOR DI(146) XOR DI(901) XOR DI(813) XOR DI(989) XOR DI(460) XOR DI(702) XOR DI(633) XOR DI(5) XOR DI(886) XOR DI(657) XOR DI(15) XOR DI(278) XOR DI(325) XOR DI(652) XOR DI(606) XOR DI(933) XOR DI(30) XOR DI(293) XOR DI(556) XOR DI(37) XOR DI(910) XOR DI(401) XOR DI(205) XOR DI(826) XOR DI(405) XOR DI(368) XOR DI(528) XOR DI(340) XOR DI(421) XOR DI(157) XOR DI(806) XOR DI(201) XOR DI(434) XOR DI(232) XOR DI(871) XOR DI(642) XOR DI(310) XOR DI(14) XOR DI(60) XOR DI(408) XOR DI(384) XOR DI(110) XOR DI(174) XOR DI(498) XOR DI(118) XOR DI(459) XOR DI(24) XOR DI(550) XOR DI(904) XOR DI(947) XOR DI(141) XOR DI(362) XOR DI(204) XOR DI(334) XOR DI(428) XOR DI(463) XOR DI(525) XOR DI(202) XOR DI(492) XOR DI(453) XOR DI(544) XOR DI(145) XOR DI(2) XOR DI(519) XOR DI(615) XOR DI(372) XOR DI(447) XOR DI(935) XOR DI(853) XOR DI(513) XOR DI(480) XOR DI(532) XOR DI(133) XOR DI(681) XOR DI(520) XOR DI(514) XOR DI(1008) XOR DI(1014) XOR DI(1020);
   DO(17) <= DI(775) XOR DI(840) XOR DI(51) XOR DI(637) XOR DI(357) XOR DI(93) XOR DI(338) XOR DI(841) XOR DI(770) XOR DI(591) XOR DI(799) XOR DI(303) XOR DI(473) XOR DI(94) XOR DI(564) XOR DI(155) XOR DI(360) XOR DI(1006) XOR DI(779) XOR DI(249) XOR DI(242) XOR DI(912) XOR DI(844) XOR DI(566) XOR DI(1000) XOR DI(225) XOR DI(713) XOR DI(594) XOR DI(308) XOR DI(386) XOR DI(929) XOR DI(260) XOR DI(802) XOR DI(867) XOR DI(56) XOR DI(979) XOR DI(358) XOR DI(191) XOR DI(1016) XOR DI(899) XOR DI(695) XOR DI(780) XOR DI(815) XOR DI(224) XOR DI(880) XOR DI(846) XOR DI(636) XOR DI(190) XOR DI(32) XOR DI(689) XOR DI(801) XOR DI(930) XOR DI(593) XOR DI(950) XOR DI(198) XOR DI(431) XOR DI(980) XOR DI(286) XOR DI(944) XOR DI(359) XOR DI(696) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(1017) XOR DI(304) XOR DI(48) XOR DI(868) XOR DI(64) XOR DI(836) XOR DI(964) XOR DI(575) XOR DI(697) XOR DI(477) XOR DI(99) XOR DI(670) XOR DI(432) XOR DI(226) XOR DI(52) XOR DI(619) XOR DI(517) XOR DI(913) XOR DI(423) XOR DI(610) XOR DI(243) XOR DI(707) XOR DI(283) XOR DI(192) XOR DI(269) XOR DI(34) XOR DI(561) XOR DI(112) XOR DI(691) XOR DI(969) XOR DI(250) XOR DI(1003) XOR DI(776) XOR DI(439) XOR DI(474) XOR DI(803) XOR DI(393) XOR DI(19) XOR DI(900) XOR DI(324) XOR DI(165) XOR DI(136) XOR DI(825) XOR DI(339) XOR DI(200) XOR DI(231) XOR DI(641) XOR DI(309) XOR DI(59) XOR DI(626) XOR DI(383) XOR DI(497) XOR DI(666) XOR DI(946) XOR DI(361) XOR DI(452) XOR DI(126) XOR DI(1019) XOR DI(765) XOR DI(276) XOR DI(864) XOR DI(442) XOR DI(85) XOR DI(333) XOR DI(305) XOR DI(568) XOR DI(975) XOR DI(555) XOR DI(49) XOR DI(685) XOR DI(792) XOR DI(834) XOR DI(329) XOR DI(972) XOR DI(730) XOR DI(45) XOR DI(837) XOR DI(965) XOR DI(962) XOR DI(548) XOR DI(952) XOR DI(149) XOR DI(1) XOR DI(183) XOR DI(478) XOR DI(994) XOR DI(494) XOR DI(586) XOR DI(222) XOR DI(710) XOR DI(100) XOR DI(185) XOR DI(433) XOR DI(288) XOR DI(169) XOR DI(53) XOR DI(371) XOR DI(424) XOR DI(743) XOR DI(876) XOR DI(400) XOR DI(654) XOR DI(604) XOR DI(416) XOR DI(26) XOR DI(72) XOR DI(420) XOR DI(768) XOR DI(105) XOR DI(220) XOR DI(708) XOR DI(11) XOR DI(255) XOR DI(284) XOR DI(28) XOR DI(331) XOR DI(471) XOR DI(270) XOR DI(79) XOR DI(345) XOR DI(786) XOR DI(916) XOR DI(407) XOR DI(755) XOR DI(570) XOR DI(113) XOR DI(692) XOR DI(970) XOR DI(251) XOR DI(216) XOR DI(534) XOR DI(919) XOR DI(1004) XOR DI(427) XOR DI(777) XOR DI(746) XOR DI(715) XOR DI(449) XOR DI(163) XOR DI(741) XOR DI(475) XOR DI(804) XOR DI(598) XOR DI(316) XOR DI(20) XOR DI(901) XOR DI(537) XOR DI(888) XOR DI(657) XOR DI(278) XOR DI(390) XOR DI(325) XOR DI(116) XOR DI(606) XOR DI(504) XOR DI(264) XOR DI(293) XOR DI(596) XOR DI(166) XOR DI(340) XOR DI(806) XOR DI(817) XOR DI(506) XOR DI(201) XOR DI(267) XOR DI(642) XOR DI(234) XOR DI(310) XOR DI(14) XOR DI(60) XOR DI(627) XOR DI(651) XOR DI(272) XOR DI(384) XOR DI(646) XOR DI(498) XOR DI(459) XOR DI(550) XOR DI(667) XOR DI(947) XOR DI(141) XOR DI(362) XOR DI(151) XOR DI(195) XOR DI(525) XOR DI(378) XOR DI(453) XOR DI(661) XOR DI(457) XOR DI(615) XOR DI(935) XOR DI(853) XOR DI(133) XOR DI(681) XOR DI(1008) XOR DI(1020) XOR DI(997) XOR DI(584) XOR DI(766) XOR DI(773) XOR DI(43) XOR DI(277) XOR DI(865) XOR DI(585) XOR DI(443) XOR DI(299) XOR DI(377) XOR DI(831) XOR DI(327) XOR DI(42) XOR DI(794) XOR DI(306) XOR DI(852) XOR DI(352) XOR DI(686) XOR DI(793) XOR DI(923) XOR DI(330) XOR DI(762) XOR DI(731) XOR DI(103) XOR DI(298) XOR DI(559) XOR DI(752) XOR DI(828) XOR DI(549) XOR DI(953) XOR DI(436) XOR DI(150) XOR DI(635) XOR DI(355) XOR DI(577) XOR DI(701) XOR DI(120) XOR DI(446) XOR DI(160) XOR DI(218) XOR DI(602) XOR DI(237) XOR DI(492) XOR DI(63) XOR DI(630) XOR DI(2) XOR DI(184) XOR DI(104) XOR DI(365) XOR DI(479) XOR DI(910) XOR DI(528) XOR DI(381) XOR DI(171) XOR DI(924) XOR DI(223) XOR DI(301) XOR DI(5) XOR DI(974) XOR DI(353) XOR DI(186) XOR DI(764) XOR DI(894) XOR DI(297) XOR DI(560) XOR DI(214) XOR DI(121) XOR DI(663) XOR DI(748) XOR DI(885) XOR DI(744) XOR DI(280) XOR DI(612) XOR DI(438) XOR DI(482) XOR DI(811) XOR DI(724) XOR DI(401) XOR DI(884) XOR DI(247) XOR DI(605) XOR DI(502) XOR DI(463) XOR DI(68) XOR DI(319) XOR DI(908) XOR DI(820) XOR DI(958) XOR DI(544) XOR DI(135) XOR DI(106) XOR DI(410) XOR DI(467) XOR DI(709) XOR DI(893) XOR DI(172) XOR DI(925) XOR DI(664) XOR DI(256) XOR DI(29) XOR DI(614) XOR DI(397) XOR DI(863) XOR DI(659) XOR DI(939) XOR DI(354) XOR DI(194) XOR DI(940) XOR DI(851) XOR DI(511) XOR DI(927) XOR DI(1012) XOR DI(991) XOR DI(760) XOR DI(37) XOR DI(859) XOR DI(80) XOR DI(321) XOR DI(36) XOR DI(563) XOR DI(44) XOR DI(82) XOR DI(346) XOR DI(680) XOR DI(787) XOR DI(829) XOR DI(408) XOR DI(967) XOR DI(756) XOR DI(603) XOR DI(292) XOR DI(960) XOR DI(822) XOR DI(430) XOR DI(349) XOR DI(571) XOR DI(154) XOR DI(971) XOR DI(833) XOR DI(904) XOR DI(412) XOR DI(489) XOR DI(791) XOR DI(252) XOR DI(217) XOR DI(968) XOR DI(535) XOR DI(347) XOR DI(920) XOR DI(124) XOR DI(778) XOR DI(716) XOR DI(450) XOR DI(164) XOR DI(824) XOR DI(513) XOR DI(115) XOR DI(742) XOR DI(419) XOR DI(213) XOR DI(239) XOR DI(805) XOR DI(718) XOR DI(625) XOR DI(649) XOR DI(241) XOR DI(317) XOR DI(411) XOR DI(62) XOR DI(147) XOR DI(902) XOR DI(814) XOR DI(990) XOR DI(461) XOR DI(703) XOR DI(634) XOR DI(6) XOR DI(887) XOR DI(658) XOR DI(16) XOR DI(279) XOR DI(326) XOR DI(653) XOR DI(607) XOR DI(934) XOR DI(31) XOR DI(294) XOR DI(557) XOR DI(38) XOR DI(911) XOR DI(402) XOR DI(206) XOR DI(827) XOR DI(406) XOR DI(369) XOR DI(529) XOR DI(341) XOR DI(422) XOR DI(158) XOR DI(807) XOR DI(202) XOR DI(435) XOR DI(233) XOR DI(872) XOR DI(643) XOR DI(311) XOR DI(15) XOR DI(61) XOR DI(409) XOR DI(0) XOR DI(385) XOR DI(111) XOR DI(175) XOR DI(499) XOR DI(119) XOR DI(460) XOR DI(25) XOR DI(551) XOR DI(905) XOR DI(948) XOR DI(142) XOR DI(363) XOR DI(205) XOR DI(335) XOR DI(429) XOR DI(464) XOR DI(526) XOR DI(203) XOR DI(493) XOR DI(454) XOR DI(545) XOR DI(146) XOR DI(3) XOR DI(520) XOR DI(616) XOR DI(373) XOR DI(448) XOR DI(936) XOR DI(854) XOR DI(514) XOR DI(481) XOR DI(533) XOR DI(134) XOR DI(682) XOR DI(521) XOR DI(515) XOR DI(1009) XOR DI(1015) XOR DI(1021);
   DO(18) <= DI(776) XOR DI(841) XOR DI(52) XOR DI(638) XOR DI(358) XOR DI(94) XOR DI(339) XOR DI(842) XOR DI(771) XOR DI(592) XOR DI(800) XOR DI(304) XOR DI(474) XOR DI(95) XOR DI(565) XOR DI(156) XOR DI(361) XOR DI(1007) XOR DI(780) XOR DI(250) XOR DI(243) XOR DI(913) XOR DI(845) XOR DI(567) XOR DI(1001) XOR DI(226) XOR DI(714) XOR DI(595) XOR DI(309) XOR DI(387) XOR DI(930) XOR DI(261) XOR DI(803) XOR DI(868) XOR DI(57) XOR DI(980) XOR DI(359) XOR DI(192) XOR DI(1017) XOR DI(900) XOR DI(696) XOR DI(781) XOR DI(816) XOR DI(225) XOR DI(881) XOR DI(847) XOR DI(637) XOR DI(191) XOR DI(33) XOR DI(690) XOR DI(802) XOR DI(931) XOR DI(594) XOR DI(951) XOR DI(199) XOR DI(432) XOR DI(981) XOR DI(287) XOR DI(945) XOR DI(360) XOR DI(697) XOR DI(857) XOR DI(517) XOR DI(484) XOR DI(1018) XOR DI(305) XOR DI(49) XOR DI(869) XOR DI(65) XOR DI(837) XOR DI(965) XOR DI(576) XOR DI(698) XOR DI(478) XOR DI(100) XOR DI(671) XOR DI(433) XOR DI(227) XOR DI(53) XOR DI(620) XOR DI(518) XOR DI(914) XOR DI(424) XOR DI(611) XOR DI(244) XOR DI(708) XOR DI(284) XOR DI(193) XOR DI(270) XOR DI(35) XOR DI(562) XOR DI(113) XOR DI(692) XOR DI(970) XOR DI(251) XOR DI(1004) XOR DI(777) XOR DI(440) XOR DI(475) XOR DI(804) XOR DI(394) XOR DI(20) XOR DI(901) XOR DI(325) XOR DI(166) XOR DI(137) XOR DI(826) XOR DI(340) XOR DI(201) XOR DI(232) XOR DI(642) XOR DI(310) XOR DI(60) XOR DI(627) XOR DI(384) XOR DI(498) XOR DI(667) XOR DI(947) XOR DI(362) XOR DI(453) XOR DI(127) XOR DI(1020) XOR DI(766) XOR DI(277) XOR DI(865) XOR DI(443) XOR DI(86) XOR DI(334) XOR DI(306) XOR DI(569) XOR DI(976) XOR DI(556) XOR DI(50) XOR DI(686) XOR DI(793) XOR DI(835) XOR DI(330) XOR DI(973) XOR DI(731) XOR DI(46) XOR DI(838) XOR DI(966) XOR DI(963) XOR DI(549) XOR DI(953) XOR DI(150) XOR DI(2) XOR DI(184) XOR DI(479) XOR DI(995) XOR DI(495) XOR DI(587) XOR DI(223) XOR DI(711) XOR DI(101) XOR DI(186) XOR DI(434) XOR DI(289) XOR DI(170) XOR DI(54) XOR DI(372) XOR DI(425) XOR DI(744) XOR DI(877) XOR DI(401) XOR DI(655) XOR DI(605) XOR DI(417) XOR DI(27) XOR DI(73) XOR DI(421) XOR DI(769) XOR DI(106) XOR DI(221) XOR DI(709) XOR DI(12) XOR DI(256) XOR DI(285) XOR DI(29) XOR DI(332) XOR DI(472) XOR DI(271) XOR DI(80) XOR DI(346) XOR DI(787) XOR DI(917) XOR DI(408) XOR DI(756) XOR DI(571) XOR DI(114) XOR DI(693) XOR DI(971) XOR DI(252) XOR DI(217) XOR DI(535) XOR DI(920) XOR DI(1005) XOR DI(428) XOR DI(778) XOR DI(747) XOR DI(716) XOR DI(450) XOR DI(164) XOR DI(742) XOR DI(476) XOR DI(805) XOR DI(599) XOR DI(317) XOR DI(21) XOR DI(902) XOR DI(538) XOR DI(889) XOR DI(658) XOR DI(279) XOR DI(391) XOR DI(326) XOR DI(117) XOR DI(607) XOR DI(505) XOR DI(265) XOR DI(294) XOR DI(597) XOR DI(167) XOR DI(341) XOR DI(807) XOR DI(818) XOR DI(507) XOR DI(202) XOR DI(268) XOR DI(643) XOR DI(235) XOR DI(311) XOR DI(15) XOR DI(61) XOR DI(628) XOR DI(0) XOR DI(652) XOR DI(273) XOR DI(385) XOR DI(647) XOR DI(499) XOR DI(460) XOR DI(551) XOR DI(668) XOR DI(948) XOR DI(142) XOR DI(363) XOR DI(152) XOR DI(196) XOR DI(526) XOR DI(379) XOR DI(454) XOR DI(662) XOR DI(458) XOR DI(616) XOR DI(936) XOR DI(854) XOR DI(134) XOR DI(682) XOR DI(1009) XOR DI(1021) XOR DI(998) XOR DI(585) XOR DI(767) XOR DI(774) XOR DI(44) XOR DI(278) XOR DI(866) XOR DI(586) XOR DI(444) XOR DI(300) XOR DI(378) XOR DI(832) XOR DI(328) XOR DI(43) XOR DI(795) XOR DI(307) XOR DI(853) XOR DI(353) XOR DI(687) XOR DI(794) XOR DI(924) XOR DI(331) XOR DI(763) XOR DI(732) XOR DI(104) XOR DI(299) XOR DI(560) XOR DI(753) XOR DI(829) XOR DI(550) XOR DI(954) XOR DI(437) XOR DI(151) XOR DI(636) XOR DI(356) XOR DI(578) XOR DI(702) XOR DI(121) XOR DI(447) XOR DI(161) XOR DI(219) XOR DI(603) XOR DI(238) XOR DI(493) XOR DI(64) XOR DI(631) XOR DI(3) XOR DI(185) XOR DI(105) XOR DI(366) XOR DI(480) XOR DI(911) XOR DI(529) XOR DI(382) XOR DI(172) XOR DI(925) XOR DI(224) XOR DI(302) XOR DI(6) XOR DI(975) XOR DI(354) XOR DI(187) XOR DI(765) XOR DI(895) XOR DI(298) XOR DI(561) XOR DI(215) XOR DI(122) XOR DI(664) XOR DI(749) XOR DI(886) XOR DI(745) XOR DI(281) XOR DI(613) XOR DI(439) XOR DI(483) XOR DI(812) XOR DI(725) XOR DI(402) XOR DI(885) XOR DI(248) XOR DI(606) XOR DI(503) XOR DI(464) XOR DI(69) XOR DI(320) XOR DI(909) XOR DI(821) XOR DI(959) XOR DI(545) XOR DI(136) XOR DI(107) XOR DI(411) XOR DI(468) XOR DI(710) XOR DI(894) XOR DI(173) XOR DI(926) XOR DI(665) XOR DI(257) XOR DI(30) XOR DI(615) XOR DI(398) XOR DI(864) XOR DI(660) XOR DI(940) XOR DI(355) XOR DI(195) XOR DI(941) XOR DI(852) XOR DI(512) XOR DI(928) XOR DI(1013) XOR DI(992) XOR DI(761) XOR DI(38) XOR DI(860) XOR DI(81) XOR DI(322) XOR DI(37) XOR DI(564) XOR DI(45) XOR DI(83) XOR DI(347) XOR DI(681) XOR DI(788) XOR DI(830) XOR DI(409) XOR DI(968) XOR DI(757) XOR DI(604) XOR DI(293) XOR DI(961) XOR DI(823) XOR DI(431) XOR DI(350) XOR DI(572) XOR DI(155) XOR DI(972) XOR DI(834) XOR DI(905) XOR DI(413) XOR DI(490) XOR DI(792) XOR DI(253) XOR DI(218) XOR DI(969) XOR DI(536) XOR DI(348) XOR DI(921) XOR DI(125) XOR DI(779) XOR DI(717) XOR DI(451) XOR DI(165) XOR DI(825) XOR DI(514) XOR DI(116) XOR DI(743) XOR DI(420) XOR DI(214) XOR DI(240) XOR DI(806) XOR DI(719) XOR DI(626) XOR DI(650) XOR DI(242) XOR DI(318) XOR DI(412) XOR DI(63) XOR DI(148) XOR DI(903) XOR DI(815) XOR DI(991) XOR DI(462) XOR DI(704) XOR DI(635) XOR DI(7) XOR DI(888) XOR DI(659) XOR DI(17) XOR DI(280) XOR DI(327) XOR DI(654) XOR DI(608) XOR DI(935) XOR DI(32) XOR DI(295) XOR DI(558) XOR DI(39) XOR DI(912) XOR DI(403) XOR DI(207) XOR DI(828) XOR DI(407) XOR DI(370) XOR DI(530) XOR DI(342) XOR DI(423) XOR DI(159) XOR DI(808) XOR DI(203) XOR DI(436) XOR DI(234) XOR DI(873) XOR DI(644) XOR DI(312) XOR DI(16) XOR DI(62) XOR DI(410) XOR DI(1) XOR DI(386) XOR DI(112) XOR DI(176) XOR DI(500) XOR DI(120) XOR DI(461) XOR DI(26) XOR DI(552) XOR DI(906) XOR DI(949) XOR DI(143) XOR DI(364) XOR DI(206) XOR DI(336) XOR DI(430) XOR DI(465) XOR DI(527) XOR DI(204) XOR DI(494) XOR DI(455) XOR DI(546) XOR DI(147) XOR DI(4) XOR DI(521) XOR DI(617) XOR DI(374) XOR DI(449) XOR DI(937) XOR DI(855) XOR DI(515) XOR DI(482) XOR DI(534) XOR DI(135) XOR DI(683) XOR DI(522) XOR DI(516) XOR DI(1010) XOR DI(1016) XOR DI(1022);
   DO(19) <= DI(777) XOR DI(842) XOR DI(53) XOR DI(639) XOR DI(359) XOR DI(95) XOR DI(340) XOR DI(843) XOR DI(772) XOR DI(593) XOR DI(801) XOR DI(305) XOR DI(475) XOR DI(96) XOR DI(566) XOR DI(157) XOR DI(362) XOR DI(1008) XOR DI(781) XOR DI(251) XOR DI(244) XOR DI(914) XOR DI(846) XOR DI(568) XOR DI(1002) XOR DI(227) XOR DI(715) XOR DI(596) XOR DI(310) XOR DI(388) XOR DI(931) XOR DI(262) XOR DI(804) XOR DI(869) XOR DI(58) XOR DI(981) XOR DI(360) XOR DI(193) XOR DI(1018) XOR DI(901) XOR DI(697) XOR DI(782) XOR DI(817) XOR DI(226) XOR DI(882) XOR DI(848) XOR DI(638) XOR DI(192) XOR DI(34) XOR DI(691) XOR DI(803) XOR DI(932) XOR DI(595) XOR DI(952) XOR DI(200) XOR DI(433) XOR DI(982) XOR DI(288) XOR DI(946) XOR DI(361) XOR DI(698) XOR DI(858) XOR DI(518) XOR DI(485) XOR DI(1019) XOR DI(306) XOR DI(50) XOR DI(870) XOR DI(66) XOR DI(838) XOR DI(966) XOR DI(577) XOR DI(699) XOR DI(479) XOR DI(101) XOR DI(672) XOR DI(434) XOR DI(228) XOR DI(54) XOR DI(621) XOR DI(519) XOR DI(915) XOR DI(425) XOR DI(612) XOR DI(245) XOR DI(709) XOR DI(285) XOR DI(194) XOR DI(271) XOR DI(36) XOR DI(563) XOR DI(114) XOR DI(693) XOR DI(971) XOR DI(252) XOR DI(1005) XOR DI(778) XOR DI(441) XOR DI(476) XOR DI(805) XOR DI(395) XOR DI(21) XOR DI(902) XOR DI(326) XOR DI(167) XOR DI(138) XOR DI(827) XOR DI(341) XOR DI(202) XOR DI(233) XOR DI(643) XOR DI(311) XOR DI(61) XOR DI(628) XOR DI(0) XOR DI(385) XOR DI(499) XOR DI(668) XOR DI(948) XOR DI(363) XOR DI(454) XOR DI(128) XOR DI(1021) XOR DI(767) XOR DI(278) XOR DI(866) XOR DI(444) XOR DI(87) XOR DI(335) XOR DI(307) XOR DI(570) XOR DI(977) XOR DI(557) XOR DI(51) XOR DI(687) XOR DI(794) XOR DI(836) XOR DI(331) XOR DI(974) XOR DI(732) XOR DI(47) XOR DI(839) XOR DI(967) XOR DI(964) XOR DI(550) XOR DI(954) XOR DI(151) XOR DI(3) XOR DI(185) XOR DI(480) XOR DI(996) XOR DI(496) XOR DI(588) XOR DI(224) XOR DI(712) XOR DI(102) XOR DI(187) XOR DI(435) XOR DI(290) XOR DI(171) XOR DI(55) XOR DI(373) XOR DI(426) XOR DI(745) XOR DI(878) XOR DI(402) XOR DI(656) XOR DI(606) XOR DI(418) XOR DI(28) XOR DI(74) XOR DI(422) XOR DI(770) XOR DI(107) XOR DI(222) XOR DI(710) XOR DI(13) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(333) XOR DI(473) XOR DI(272) XOR DI(81) XOR DI(347) XOR DI(788) XOR DI(918) XOR DI(409) XOR DI(757) XOR DI(572) XOR DI(115) XOR DI(694) XOR DI(972) XOR DI(253) XOR DI(218) XOR DI(536) XOR DI(921) XOR DI(1006) XOR DI(429) XOR DI(779) XOR DI(748) XOR DI(717) XOR DI(451) XOR DI(165) XOR DI(743) XOR DI(477) XOR DI(806) XOR DI(600) XOR DI(318) XOR DI(22) XOR DI(903) XOR DI(539) XOR DI(890) XOR DI(659) XOR DI(280) XOR DI(392) XOR DI(327) XOR DI(118) XOR DI(608) XOR DI(506) XOR DI(266) XOR DI(295) XOR DI(598) XOR DI(168) XOR DI(342) XOR DI(808) XOR DI(819) XOR DI(508) XOR DI(203) XOR DI(269) XOR DI(644) XOR DI(236) XOR DI(312) XOR DI(16) XOR DI(62) XOR DI(629) XOR DI(1) XOR DI(653) XOR DI(274) XOR DI(386) XOR DI(648) XOR DI(500) XOR DI(461) XOR DI(552) XOR DI(669) XOR DI(949) XOR DI(143) XOR DI(364) XOR DI(153) XOR DI(197) XOR DI(527) XOR DI(380) XOR DI(455) XOR DI(663) XOR DI(459) XOR DI(617) XOR DI(937) XOR DI(855) XOR DI(135) XOR DI(683) XOR DI(1010) XOR DI(1022) XOR DI(999) XOR DI(586) XOR DI(768) XOR DI(775) XOR DI(45) XOR DI(279) XOR DI(867) XOR DI(587) XOR DI(445) XOR DI(301) XOR DI(379) XOR DI(833) XOR DI(329) XOR DI(44) XOR DI(796) XOR DI(308) XOR DI(854) XOR DI(354) XOR DI(688) XOR DI(795) XOR DI(925) XOR DI(332) XOR DI(764) XOR DI(733) XOR DI(105) XOR DI(300) XOR DI(561) XOR DI(754) XOR DI(830) XOR DI(551) XOR DI(955) XOR DI(438) XOR DI(152) XOR DI(637) XOR DI(357) XOR DI(579) XOR DI(703) XOR DI(122) XOR DI(448) XOR DI(162) XOR DI(220) XOR DI(604) XOR DI(239) XOR DI(494) XOR DI(65) XOR DI(632) XOR DI(4) XOR DI(186) XOR DI(106) XOR DI(367) XOR DI(481) XOR DI(912) XOR DI(530) XOR DI(383) XOR DI(173) XOR DI(926) XOR DI(225) XOR DI(303) XOR DI(7) XOR DI(976) XOR DI(355) XOR DI(188) XOR DI(766) XOR DI(896) XOR DI(299) XOR DI(562) XOR DI(216) XOR DI(123) XOR DI(665) XOR DI(750) XOR DI(887) XOR DI(746) XOR DI(282) XOR DI(614) XOR DI(440) XOR DI(484) XOR DI(813) XOR DI(726) XOR DI(403) XOR DI(886) XOR DI(249) XOR DI(607) XOR DI(504) XOR DI(465) XOR DI(70) XOR DI(321) XOR DI(910) XOR DI(822) XOR DI(960) XOR DI(546) XOR DI(137) XOR DI(108) XOR DI(412) XOR DI(469) XOR DI(711) XOR DI(895) XOR DI(174) XOR DI(927) XOR DI(666) XOR DI(258) XOR DI(31) XOR DI(616) XOR DI(399) XOR DI(865) XOR DI(661) XOR DI(941) XOR DI(356) XOR DI(196) XOR DI(942) XOR DI(853) XOR DI(513) XOR DI(929) XOR DI(1014) XOR DI(993) XOR DI(762) XOR DI(39) XOR DI(861) XOR DI(82) XOR DI(323) XOR DI(38) XOR DI(565) XOR DI(46) XOR DI(84) XOR DI(348) XOR DI(682) XOR DI(789) XOR DI(831) XOR DI(410) XOR DI(969) XOR DI(758) XOR DI(605) XOR DI(294) XOR DI(962) XOR DI(824) XOR DI(432) XOR DI(351) XOR DI(573) XOR DI(156) XOR DI(973) XOR DI(835) XOR DI(906) XOR DI(414) XOR DI(491) XOR DI(793) XOR DI(254) XOR DI(219) XOR DI(970) XOR DI(537) XOR DI(349) XOR DI(922) XOR DI(126) XOR DI(780) XOR DI(718) XOR DI(452) XOR DI(166) XOR DI(826) XOR DI(515) XOR DI(117) XOR DI(744) XOR DI(421) XOR DI(215) XOR DI(241) XOR DI(807) XOR DI(720) XOR DI(627) XOR DI(651) XOR DI(243) XOR DI(319) XOR DI(413) XOR DI(64) XOR DI(149) XOR DI(904) XOR DI(816) XOR DI(992) XOR DI(463) XOR DI(705) XOR DI(636) XOR DI(8) XOR DI(889) XOR DI(660) XOR DI(18) XOR DI(281) XOR DI(328) XOR DI(655) XOR DI(609) XOR DI(936) XOR DI(33) XOR DI(296) XOR DI(559) XOR DI(40) XOR DI(913) XOR DI(404) XOR DI(208) XOR DI(829) XOR DI(408) XOR DI(371) XOR DI(531) XOR DI(343) XOR DI(424) XOR DI(160) XOR DI(809) XOR DI(204) XOR DI(437) XOR DI(235) XOR DI(874) XOR DI(645) XOR DI(313) XOR DI(17) XOR DI(63) XOR DI(411) XOR DI(2) XOR DI(387) XOR DI(113) XOR DI(177) XOR DI(501) XOR DI(121) XOR DI(462) XOR DI(27) XOR DI(553) XOR DI(907) XOR DI(950) XOR DI(144) XOR DI(365) XOR DI(207) XOR DI(337) XOR DI(431) XOR DI(466) XOR DI(528) XOR DI(205) XOR DI(495) XOR DI(456) XOR DI(547) XOR DI(148) XOR DI(5) XOR DI(522) XOR DI(618) XOR DI(375) XOR DI(450) XOR DI(938) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(535) XOR DI(136) XOR DI(684) XOR DI(523) XOR DI(517) XOR DI(1011) XOR DI(1017) XOR DI(1023);
   DO(20) <= DI(778) XOR DI(93) XOR DI(591) XOR DI(843) XOR DI(842) XOR DI(54) XOR DI(640) XOR DI(360) XOR DI(96) XOR DI(341) XOR DI(844) XOR DI(773) XOR DI(800) XOR DI(594) XOR DI(802) XOR DI(306) XOR DI(476) XOR DI(97) XOR DI(50) XOR DI(881) XOR DI(787) XOR DI(738) XOR DI(57) XOR DI(980) XOR DI(359) XOR DI(945) XOR DI(863) XOR DI(567) XOR DI(760) XOR DI(158) XOR DI(643) XOR DI(697) XOR DI(0) XOR DI(363) XOR DI(709) XOR DI(128) XOR DI(1009) XOR DI(782) XOR DI(252) XOR DI(245) XOR DI(317) XOR DI(395) XOR DI(192) XOR DI(80) XOR DI(915) XOR DI(847) XOR DI(569) XOR DI(691) XOR DI(987) XOR DI(1003) XOR DI(228) XOR DI(716) XOR DI(597) XOR DI(311) XOR DI(277) XOR DI(389) XOR DI(932) XOR DI(263) XOR DI(805) XOR DI(200) XOR DI(870) XOR DI(233) XOR DI(59) XOR DI(982) XOR DI(271) XOR DI(361) XOR DI(194) XOR DI(479) XOR DI(1019) XOR DI(772) XOR DI(902) XOR DI(326) XOR DI(305) XOR DI(86) XOR DI(869) XOR DI(952) XOR DI(576) XOR DI(698) XOR DI(838) XOR DI(262) XOR DI(671) XOR DI(756) XOR DI(783) XOR DI(288) XOR DI(818) XOR DI(227) XOR DI(53) XOR DI(620) XOR DI(883) XOR DI(849) XOR DI(639) XOR DI(892) XOR DI(284) XOR DI(658) XOR DI(193) XOR DI(612) XOR DI(499) XOR DI(76) XOR DI(858) XOR DI(35) XOR DI(966) XOR DI(602) XOR DI(692) XOR DI(715) XOR DI(741) XOR DI(475) XOR DI(804) XOR DI(20) XOR DI(901) XOR DI(933) XOR DI(556) XOR DI(401) XOR DI(596) XOR DI(953) XOR DI(201) XOR DI(434) XOR DI(983) XOR DI(289) XOR DI(947) XOR DI(362) XOR DI(699) XOR DI(859) XOR DI(519) XOR DI(486) XOR DI(1008) XOR DI(1020) XOR DI(444) XOR DI(378) XOR DI(335) XOR DI(307) XOR DI(51) XOR DI(687) XOR DI(871) XOR DI(91) XOR DI(67) XOR DI(331) XOR DI(732) XOR DI(104) XOR DI(190) XOR DI(839) XOR DI(967) XOR DI(964) XOR DI(151) XOR DI(578) XOR DI(700) XOR DI(185) XOR DI(480) XOR DI(996) XOR DI(382) XOR DI(798) XOR DI(224) XOR DI(634) XOR DI(102) XOR DI(131) XOR DI(673) XOR DI(435) XOR DI(369) XOR DI(171) XOR DI(229) XOR DI(55) XOR DI(622) XOR DI(520) XOR DI(916) XOR DI(426) XOR DI(613) XOR DI(246) XOR DI(812) XOR DI(248) XOR DI(418) XOR DI(503) XOR DI(74) XOR DI(959) XOR DI(545) XOR DI(222) XOR DI(710) XOR DI(13) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(398) XOR DI(195) XOR DI(473) XOR DI(680) XOR DI(272) XOR DI(37) XOR DI(564) XOR DI(918) XOR DI(293) XOR DI(572) XOR DI(115) XOR DI(694) XOR DI(972) XOR DI(990) XOR DI(490) XOR DI(253) XOR DI(218) XOR DI(921) XOR DI(1006) XOR DI(429) XOR DI(779) XOR DI(748) XOR DI(165) XOR DI(442) XOR DI(730) XOR DI(231) XOR DI(477) XOR DI(806) XOR DI(396) XOR DI(626) XOR DI(650) XOR DI(600) XOR DI(22) XOR DI(903) XOR DI(392) XOR DI(327) XOR DI(182) XOR DI(506) XOR DI(266) XOR DI(168) XOR DI(139) XOR DI(828) XOR DI(899) XOR DI(407) XOR DI(342) XOR DI(508) XOR DI(203) XOR DI(269) XOR DI(234) XOR DI(873) XOR DI(644) XOR DI(312) XOR DI(16) XOR DI(62) XOR DI(722) XOR DI(629) XOR DI(1) XOR DI(274) XOR DI(386) XOR DI(648) XOR DI(176) XOR DI(500) XOR DI(461) XOR DI(26) XOR DI(669) XOR DI(949) XOR DI(143) XOR DI(364) XOR DI(707) XOR DI(455) XOR DI(459) XOR DI(141) XOR DI(135) XOR DI(129) XOR DI(677) XOR DI(510) XOR DI(1022) XOR DI(575) XOR DI(268) XOR DI(999) XOR DI(768) XOR DI(279) XOR DI(867) XOR DI(445) XOR DI(88) XOR DI(336) XOR DI(833) XOR DI(44) XOR DI(308) XOR DI(184) XOR DI(571) XOR DI(978) XOR DI(558) XOR DI(52) XOR DI(89) XOR DI(49) XOR DI(170) XOR DI(90) XOR DI(354) XOR DI(688) XOR DI(795) XOR DI(925) XOR DI(837) XOR DI(332) XOR DI(975) XOR DI(733) XOR DI(48) XOR DI(840) XOR DI(995) XOR DI(968) XOR DI(965) XOR DI(551) XOR DI(958) XOR DI(955) XOR DI(152) XOR DI(703) XOR DI(736) XOR DI(239) XOR DI(494) XOR DI(632) XOR DI(4) XOR DI(186) XOR DI(979) XOR DI(841) XOR DI(481) XOR DI(997) XOR DI(420) XOR DI(530) XOR DI(173) XOR DI(497) XOR DI(589) XOR DI(225) XOR DI(303) XOR DI(976) XOR DI(713) XOR DI(103) XOR DI(543) XOR DI(940) XOR DI(188) XOR DI(436) XOR DI(299) XOR DI(724) XOR DI(291) XOR DI(172) XOR DI(821) XOR DI(542) XOR DI(56) XOR DI(374) XOR DI(665) XOR DI(750) XOR DI(427) XOR DI(746) XOR DI(533) XOR DI(512) XOR DI(737) XOR DI(212) XOR DI(238) XOR DI(728) XOR DI(879) XOR DI(726) XOR DI(403) XOR DI(657) XOR DI(15) XOR DI(607) XOR DI(419) XOR DI(493) XOR DI(70) XOR DI(852) XOR DI(29) XOR DI(155) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(423) XOR DI(147) XOR DI(686) XOR DI(998) XOR DI(771) XOR DI(108) XOR DI(223) XOR DI(469) XOR DI(711) XOR DI(14) XOR DI(24) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(616) XOR DI(334) XOR DI(428) XOR DI(544) XOR DI(941) XOR DI(125) XOR DI(853) XOR DI(513) XOR DI(929) XOR DI(133) XOR DI(474) XOR DI(1014) XOR DI(273) XOR DI(82) XOR DI(323) XOR DI(43) XOR DI(164) XOR DI(348) XOR DI(682) XOR DI(789) XOR DI(919) XOR DI(410) XOR DI(969) XOR DI(758) XOR DI(42) XOR DI(146) XOR DI(631) XOR DI(351) XOR DI(573) XOR DI(116) XOR DI(156) XOR DI(214) XOR DI(695) XOR DI(973) XOR DI(679) XOR DI(906) XOR DI(920) XOR DI(254) XOR DI(219) XOR DI(537) XOR DI(922) XOR DI(126) XOR DI(1007) XOR DI(430) XOR DI(780) XOR DI(749) XOR DI(718) XOR DI(452) XOR DI(166) XOR DI(815) XOR DI(826) XOR DI(210) XOR DI(117) XOR DI(744) XOR DI(421) XOR DI(276) XOR DI(215) XOR DI(478) XOR DI(807) XOR DI(880) XOR DI(601) XOR DI(319) XOR DI(498) XOR DI(23) XOR DI(69) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(417) XOR DI(891) XOR DI(992) XOR DI(729) XOR DI(705) XOR DI(636) XOR DI(889) XOR DI(660) XOR DI(281) XOR DI(25) XOR DI(393) XOR DI(328) XOR DI(655) XOR DI(119) XOR DI(609) XOR DI(507) XOR DI(468) XOR DI(675) XOR DI(267) XOR DI(296) XOR DI(559) XOR DI(676) XOR DI(599) XOR DI(169) XOR DI(625) XOR DI(371) XOR DI(213) XOR DI(343) XOR DI(120) XOR DI(424) XOR DI(809) XOR DI(820) XOR DI(509) XOR DI(204) XOR DI(270) XOR DI(437) XOR DI(725) XOR DI(714) XOR DI(645) XOR DI(237) XOR DI(313) XOR DI(17) XOR DI(63) XOR DI(898) XOR DI(534) XOR DI(211) XOR DI(630) XOR DI(2) XOR DI(654) XOR DI(12) XOR DI(275) XOR DI(387) XOR DI(292) XOR DI(649) XOR DI(501) XOR DI(121) XOR DI(462) XOR DI(261) XOR DI(553) XOR DI(670) XOR DI(957) XOR DI(950) XOR DI(134) XOR DI(144) XOR DI(365) XOR DI(337) XOR DI(154) XOR DI(198) XOR DI(431) XOR DI(528) XOR DI(394) XOR DI(624) XOR DI(381) XOR DI(316) XOR DI(456) XOR DI(664) XOR DI(148) XOR DI(460) XOR DI(702) XOR DI(522) XOR DI(199) XOR DI(618) XOR DI(375) XOR DI(489) XOR DI(450) XOR DI(541) XOR DI(938) XOR DI(696) XOR DI(856) XOR DI(535) XOR DI(136) XOR DI(690) XOR DI(684) XOR DI(1011) XOR DI(1023);
   DO(21) <= DI(93) XOR DI(776) XOR DI(779) XOR DI(638) XOR DI(94) XOR DI(798) XOR DI(592) XOR DI(800) XOR DI(767) XOR DI(844) XOR DI(843) XOR DI(55) XOR DI(943) XOR DI(580) XOR DI(439) XOR DI(641) XOR DI(361) XOR DI(707) XOR DI(97) XOR DI(250) XOR DI(873) XOR DI(190) XOR DI(342) XOR DI(845) XOR DI(248) XOR DI(774) XOR DI(801) XOR DI(595) XOR DI(803) XOR DI(231) XOR DI(307) XOR DI(107) XOR DI(359) XOR DI(192) XOR DI(477) XOR DI(566) XOR DI(176) XOR DI(836) XOR DI(98) XOR DI(51) XOR DI(882) XOR DI(444) XOR DI(242) XOR DI(74) XOR DI(34) XOR DI(964) XOR DI(788) XOR DI(739) XOR DI(473) XOR DI(875) XOR DI(58) XOR DI(981) XOR DI(945) XOR DI(360) XOR DI(946) XOR DI(524) XOR DI(1018) XOR DI(765) XOR DI(864) XOR DI(305) XOR DI(568) XOR DI(869) XOR DI(761) XOR DI(178) XOR DI(548) XOR DI(952) XOR DI(159) XOR DI(644) XOR DI(698) XOR DI(1) XOR DI(364) XOR DI(380) XOR DI(257) XOR DI(222) XOR DI(710) XOR DI(129) XOR DI(1010) XOR DI(763) XOR DI(433) XOR DI(783) XOR DI(620) XOR DI(518) XOR DI(914) XOR DI(253) XOR DI(244) XOR DI(246) XOR DI(318) XOR DI(732) XOR DI(284) XOR DI(28) XOR DI(396) XOR DI(331) XOR DI(193) XOR DI(858) XOR DI(81) XOR DI(916) XOR DI(407) XOR DI(848) XOR DI(570) XOR DI(485) XOR DI(692) XOR DI(988) XOR DI(1004) XOR DI(741) XOR DI(229) XOR DI(717) XOR DI(648) XOR DI(598) XOR DI(312) XOR DI(20) XOR DI(901) XOR DI(278) XOR DI(390) XOR DI(295) XOR DI(606) XOR DI(933) XOR DI(264) XOR DI(405) XOR DI(806) XOR DI(506) XOR DI(201) XOR DI(871) XOR DI(234) XOR DI(60) XOR DI(983) XOR DI(272) XOR DI(384) XOR DI(459) XOR DI(667) XOR DI(141) XOR DI(362) XOR DI(151) XOR DI(195) XOR DI(378) XOR DI(480) XOR DI(1020) XOR DI(266) XOR DI(773) XOR DI(903) XOR DI(86) XOR DI(327) XOR DI(794) XOR DI(306) XOR DI(182) XOR DI(556) XOR DI(87) XOR DI(937) XOR DI(47) XOR DI(870) XOR DI(66) XOR DI(855) XOR DI(953) XOR DI(577) XOR DI(218) XOR DI(699) XOR DI(839) XOR DI(263) XOR DI(672) XOR DI(757) XOR DI(784) XOR DI(722) XOR DI(289) XOR DI(819) XOR DI(228) XOR DI(54) XOR DI(621) XOR DI(748) XOR DI(612) XOR DI(236) XOR DI(401) XOR DI(884) XOR DI(850) XOR DI(908) XOR DI(709) XOR DI(640) XOR DI(893) XOR DI(285) XOR DI(588) XOR DI(863) XOR DI(659) XOR DI(143) XOR DI(194) XOR DI(613) XOR DI(131) XOR DI(500) XOR DI(760) XOR DI(77) XOR DI(859) XOR DI(80) XOR DI(36) XOR DI(563) XOR DI(787) XOR DI(967) XOR DI(756) XOR DI(603) XOR DI(987) XOR DI(114) XOR DI(693) XOR DI(971) XOR DI(918) XOR DI(716) XOR DI(742) XOR DI(441) XOR DI(476) XOR DI(805) XOR DI(496) XOR DI(21) XOR DI(902) XOR DI(415) XOR DI(990) XOR DI(634) XOR DI(6) XOR DI(326) XOR DI(934) XOR DI(557) XOR DI(402) XOR DI(961) XOR DI(597) XOR DI(954) XOR DI(138) XOR DI(206) XOR DI(369) XOR DI(202) XOR DI(435) XOR DI(233) XOR DI(643) XOR DI(409) XOR DI(984) XOR DI(398) XOR DI(628) XOR DI(0) XOR DI(652) XOR DI(290) XOR DI(948) XOR DI(161) XOR DI(363) XOR DI(812) XOR DI(464) XOR DI(866) XOR DI(9) XOR DI(392) XOR DI(662) XOR DI(700) XOR DI(860) XOR DI(520) XOR DI(197) XOR DI(487) XOR DI(128) XOR DI(503) XOR DI(1009) XOR DI(1021) XOR DI(575) XOR DI(41) XOR DI(85) XOR DI(587) XOR DI(445) XOR DI(301) XOR DI(379) XOR DI(336) XOR DI(833) XOR DI(994) XOR DI(308) XOR DI(184) XOR DI(52) XOR DI(354) XOR DI(688) XOR DI(872) XOR DI(92) XOR DI(925) XOR DI(68) XOR DI(332) XOR DI(733) XOR DI(105) XOR DI(191) XOR DI(840) XOR DI(467) XOR DI(995) XOR DI(968) XOR DI(965) XOR DI(830) XOR DI(152) XOR DI(357) XOR DI(579) XOR DI(736) XOR DI(65) XOR DI(701) XOR DI(186) XOR DI(106) XOR DI(481) XOR DI(997) XOR DI(797) XOR DI(530) XOR DI(383) XOR DI(799) XOR DI(225) XOR DI(635) XOR DI(303) XOR DI(103) XOR DI(940) XOR DI(928) XOR DI(132) XOR DI(674) XOR DI(896) XOR DI(436) XOR DI(370) XOR DI(299) XOR DI(562) XOR DI(755) XOR DI(724) XOR DI(172) XOR DI(230) XOR DI(56) XOR DI(623) XOR DI(832) XOR DI(358) XOR DI(521) XOR DI(917) XOR DI(123) XOR DI(887) XOR DI(427) XOR DI(449) XOR DI(533) XOR DI(221) XOR DI(614) XOR DI(512) XOR DI(247) XOR DI(728) XOR DI(484) XOR DI(813) XOR DI(888) XOR DI(249) XOR DI(419) XOR DI(504) XOR DI(493) XOR DI(852) XOR DI(75) XOR DI(910) XOR DI(960) XOR DI(546) XOR DI(686) XOR DI(897) XOR DI(412) XOR DI(223) XOR DI(711) XOR DI(14) XOR DI(927) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(616) XOR DI(399) XOR DI(283) XOR DI(125) XOR DI(356) XOR DI(196) XOR DI(615) XOR DI(532) XOR DI(929) XOR DI(133) XOR DI(474) XOR DI(681) XOR DI(1014) XOR DI(39) XOR DI(273) XOR DI(330) XOR DI(323) XOR DI(38) XOR DI(302) XOR DI(565) XOR DI(46) XOR DI(164) XOR DI(682) XOR DI(919) XOR DI(831) XOR DI(605) XOR DI(42) XOR DI(294) XOR DI(175) XOR DI(146) XOR DI(351) XOR DI(573) XOR DI(116) XOR DI(695) XOR DI(973) XOR DI(679) XOR DI(906) XOR DI(991) XOR DI(414) XOR DI(491) XOR DI(254) XOR DI(219) XOR DI(922) XOR DI(1007) XOR DI(430) XOR DI(780) XOR DI(749) XOR DI(166) XOR DI(815) XOR DI(826) XOR DI(368) XOR DI(210) XOR DI(443) XOR DI(731) XOR DI(232) XOR DI(478) XOR DI(807) XOR DI(397) XOR DI(627) XOR DI(651) XOR DI(601) XOR DI(413) XOR DI(23) XOR DI(69) XOR DI(904) XOR DI(417) XOR DI(992) XOR DI(217) XOR DI(705) XOR DI(636) XOR DI(8) XOR DI(889) XOR DI(393) XOR DI(328) XOR DI(350) XOR DI(183) XOR DI(507) XOR DI(468) XOR DI(675) XOR DI(267) XOR DI(40) XOR DI(913) XOR DI(825) XOR DI(963) XOR DI(721) XOR DI(169) XOR DI(140) XOR DI(150) XOR DI(208) XOR DI(829) XOR DI(900) XOR DI(408) XOR DI(371) XOR DI(343) XOR DI(509) XOR DI(204) XOR DI(270) XOR DI(209) XOR DI(235) XOR DI(874) XOR DI(645) XOR DI(313) XOR DI(492) XOR DI(17) XOR DI(63) XOR DI(898) XOR DI(723) XOR DI(400) XOR DI(630) XOR DI(2) XOR DI(12) XOR DI(275) XOR DI(19) XOR DI(387) XOR DI(322) XOR DI(649) XOR DI(177) XOR DI(501) XOR DI(462) XOR DI(27) XOR DI(261) XOR DI(670) XOR DI(957) XOR DI(950) XOR DI(163) XOR DI(144) XOR DI(365) XOR DI(814) XOR DI(466) XOR DI(708) XOR DI(624) XOR DI(316) XOR DI(456) XOR DI(547) XOR DI(460) XOR DI(702) XOR DI(862) XOR DI(522) XOR DI(489) XOR DI(450) XOR DI(142) XOR DI(516) XOR DI(136) XOR DI(690) XOR DI(130) XOR DI(124) XOR DI(678) XOR DI(517) XOR DI(511) XOR DI(505) XOR DI(1023);
   DO(22) <= DI(562) XOR DI(94) XOR DI(777) XOR DI(780) XOR DI(980) XOR DI(842) XOR DI(590) XOR DI(1014) XOR DI(639) XOR DI(95) XOR DI(999) XOR DI(772) XOR DI(799) XOR DI(593) XOR DI(591) XOR DI(801) XOR DI(305) XOR DI(768) XOR DI(667) XOR DI(49) XOR DI(880) XOR DI(845) XOR DI(844) XOR DI(1000) XOR DI(56) XOR DI(979) XOR DI(944) XOR DI(581) XOR DI(862) XOR DI(440) XOR DI(790) XOR DI(970) XOR DI(759) XOR DI(157) XOR DI(642) XOR DI(362) XOR DI(708) XOR DI(98) XOR DI(127) XOR DI(453) XOR DI(251) XOR DI(741) XOR DI(874) XOR DI(881) XOR DI(244) XOR DI(316) XOR DI(191) XOR DI(343) XOR DI(846) XOR DI(690) XOR DI(249) XOR DI(775) XOR DI(802) XOR DI(715) XOR DI(596) XOR DI(338) XOR DI(804) XOR DI(199) XOR DI(869) XOR DI(232) XOR DI(308) XOR DI(108) XOR DI(945) XOR DI(360) XOR DI(193) XOR DI(478) XOR DI(1018) XOR DI(567) XOR DI(85) XOR DI(868) XOR DI(177) XOR DI(575) XOR DI(697) XOR DI(837) XOR DI(261) XOR DI(99) XOR DI(755) XOR DI(892) XOR DI(432) XOR DI(751) XOR DI(817) XOR DI(52) XOR DI(619) XOR DI(913) XOR DI(661) XOR DI(883) XOR DI(445) XOR DI(243) XOR DI(638) XOR DI(283) XOR DI(424) XOR DI(498) XOR DI(75) XOR DI(35) XOR DI(857) XOR DI(34) XOR DI(965) XOR DI(484) XOR DI(789) XOR DI(776) XOR DI(714) XOR DI(740) XOR DI(474) XOR DI(876) XOR DI(19) XOR DI(65) XOR DI(952) XOR DI(156) XOR DI(200) XOR DI(433) XOR DI(59) XOR DI(982) XOR DI(8) XOR DI(109) XOR DI(666) XOR DI(946) XOR DI(361) XOR DI(524) XOR DI(620) XOR DI(947) XOR DI(858) XOR DI(525) XOR DI(1019) XOR DI(766) XOR DI(277) XOR DI(865) XOR DI(306) XOR DI(569) XOR DI(976) XOR DI(556) XOR DI(50) XOR DI(686) XOR DI(870) XOR DI(90) XOR DI(330) XOR DI(762) XOR DI(46) XOR DI(189) XOR DI(838) XOR DI(559) XOR DI(963) XOR DI(179) XOR DI(549) XOR DI(953) XOR DI(150) XOR DI(160) XOR DI(645) XOR DI(699) XOR DI(2) XOR DI(365) XOR DI(910) XOR DI(381) XOR DI(495) XOR DI(587) XOR DI(797) XOR DI(258) XOR DI(223) XOR DI(633) XOR DI(5) XOR DI(711) XOR DI(130) XOR DI(1011) XOR DI(764) XOR DI(434) XOR DI(368) XOR DI(784) XOR DI(621) XOR DI(519) XOR DI(915) XOR DI(254) XOR DI(425) XOR DI(612) XOR DI(245) XOR DI(438) XOR DI(655) XOR DI(247) XOR DI(605) XOR DI(417) XOR DI(319) XOR DI(544) XOR DI(421) XOR DI(769) XOR DI(733) XOR DI(221) XOR DI(12) XOR DI(285) XOR DI(29) XOR DI(397) XOR DI(332) XOR DI(194) XOR DI(760) XOR DI(859) XOR DI(80) XOR DI(82) XOR DI(787) XOR DI(917) XOR DI(408) XOR DI(292) XOR DI(987) XOR DI(849) XOR DI(822) XOR DI(571) XOR DI(114) XOR DI(486) XOR DI(693) XOR DI(971) XOR DI(989) XOR DI(375) XOR DI(489) XOR DI(217) XOR DI(535) XOR DI(1005) XOR DI(747) XOR DI(742) XOR DI(738) XOR DI(441) XOR DI(239) XOR DI(230) XOR DI(718) XOR DI(395) XOR DI(649) XOR DI(599) XOR DI(313) XOR DI(21) XOR DI(902) XOR DI(538) XOR DI(404) XOR DI(658) XOR DI(279) XOR DI(391) XOR DI(326) XOR DI(296) XOR DI(607) XOR DI(934) XOR DI(71) XOR DI(265) XOR DI(138) XOR DI(406) XOR DI(807) XOR DI(507) XOR DI(202) XOR DI(470) XOR DI(872) XOR DI(643) XOR DI(235) XOR DI(61) XOR DI(984) XOR DI(721) XOR DI(0) XOR DI(273) XOR DI(385) XOR DI(175) XOR DI(499) XOR DI(460) XOR DI(25) XOR DI(668) XOR DI(142) XOR DI(363) XOR DI(152) XOR DI(196) XOR DI(379) XOR DI(662) XOR DI(942) XOR DI(854) XOR DI(481) XOR DI(128) XOR DI(1021) XOR DI(267) XOR DI(767) XOR DI(774) XOR DI(904) XOR DI(44) XOR DI(866) XOR DI(705) XOR DI(87) XOR DI(378) XOR DI(335) XOR DI(328) XOR DI(795) XOR DI(307) XOR DI(183) XOR DI(977) XOR DI(557) XOR DI(88) XOR DI(938) XOR DI(48) XOR DI(89) XOR DI(871) XOR DI(91) XOR DI(794) XOR DI(836) XOR DI(67) XOR DI(763) XOR DI(610) XOR DI(190) XOR DI(299) XOR DI(466) XOR DI(994) XOR DI(856) XOR DI(560) XOR DI(957) XOR DI(954) XOR DI(356) XOR DI(578) XOR DI(121) XOR DI(161) XOR DI(219) XOR DI(238) XOR DI(700) XOR DI(908) XOR DI(840) XOR DI(796) XOR DI(529) XOR DI(382) XOR DI(925) XOR DI(496) XOR DI(634) XOR DI(6) XOR DI(264) XOR DI(542) XOR DI(939) XOR DI(354) XOR DI(927) XOR DI(673) XOR DI(1012) XOR DI(758) XOR DI(765) XOR DI(785) XOR DI(723) XOR DI(290) XOR DI(171) XOR DI(820) XOR DI(541) XOR DI(229) XOR DI(55) XOR DI(622) XOR DI(215) XOR DI(122) XOR DI(749) XOR DI(745) XOR DI(532) XOR DI(613) XOR DI(736) XOR DI(439) XOR DI(237) XOR DI(727) XOR DI(812) XOR DI(887) XOR DI(402) XOR DI(632) XOR DI(885) XOR DI(656) XOR DI(503) XOR DI(464) XOR DI(851) XOR DI(320) XOR DI(74) XOR DI(909) XOR DI(821) XOR DI(959) XOR DI(545) XOR DI(422) XOR DI(146) XOR DI(685) XOR DI(896) XOR DI(411) XOR DI(710) XOR DI(641) XOR DI(894) XOR DI(665) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(589) XOR DI(810) XOR DI(864) XOR DI(282) XOR DI(543) XOR DI(660) XOR DI(940) XOR DI(144) XOR DI(195) XOR DI(614) XOR DI(852) XOR DI(132) XOR DI(473) XOR DI(501) XOR DI(761) XOR DI(78) XOR DI(860) XOR DI(81) XOR DI(322) XOR DI(37) XOR DI(301) XOR DI(564) XOR DI(45) XOR DI(163) XOR DI(83) XOR DI(788) XOR DI(968) XOR DI(757) XOR DI(726) XOR DI(604) XOR DI(293) XOR DI(988) XOR DI(554) XOR DI(174) XOR DI(823) XOR DI(350) XOR DI(572) XOR DI(115) XOR DI(155) XOR DI(213) XOR DI(694) XOR DI(972) XOR DI(990) XOR DI(376) XOR DI(919) XOR DI(536) XOR DI(921) XOR DI(429) XOR DI(748) XOR DI(717) XOR DI(825) XOR DI(514) XOR DI(743) XOR DI(442) XOR DI(214) XOR DI(240) XOR DI(730) XOR DI(477) XOR DI(806) XOR DI(719) XOR DI(626) XOR DI(242) XOR DI(600) XOR DI(412) XOR DI(497) XOR DI(22) XOR DI(148) XOR DI(903) XOR DI(416) XOR DI(991) XOR DI(728) XOR DI(405) XOR DI(216) XOR DI(704) XOR DI(635) XOR DI(7) XOR DI(280) XOR DI(392) XOR DI(327) XOR DI(297) XOR DI(118) XOR DI(349) XOR DI(182) XOR DI(608) XOR DI(935) XOR DI(266) XOR DI(558) XOR DI(403) XOR DI(962) XOR DI(598) XOR DI(955) XOR DI(139) XOR DI(149) XOR DI(207) XOR DI(407) XOR DI(370) XOR DI(212) XOR DI(530) XOR DI(203) XOR DI(269) XOR DI(436) XOR DI(208) XOR DI(234) XOR DI(644) XOR DI(16) XOR DI(410) XOR DI(985) XOR DI(399) XOR DI(629) XOR DI(1) XOR DI(653) XOR DI(291) XOR DI(648) XOR DI(120) XOR DI(26) XOR DI(552) XOR DI(906) XOR DI(956) XOR DI(949) XOR DI(162) XOR DI(364) XOR DI(206) XOR DI(813) XOR DI(465) XOR DI(707) XOR DI(867) XOR DI(10) XOR DI(393) XOR DI(663) XOR DI(943) XOR DI(459) XOR DI(701) XOR DI(861) XOR DI(521) XOR DI(198) XOR DI(488) XOR DI(449) XOR DI(937) XOR DI(855) XOR DI(135) XOR DI(129) XOR DI(123) XOR DI(677) XOR DI(516) XOR DI(504) XOR DI(1010) XOR DI(1022);
   DO(23) <= DI(563) XOR DI(95) XOR DI(778) XOR DI(781) XOR DI(981) XOR DI(843) XOR DI(591) XOR DI(1015) XOR DI(640) XOR DI(96) XOR DI(1000) XOR DI(773) XOR DI(800) XOR DI(594) XOR DI(592) XOR DI(802) XOR DI(306) XOR DI(769) XOR DI(668) XOR DI(50) XOR DI(881) XOR DI(846) XOR DI(845) XOR DI(1001) XOR DI(57) XOR DI(980) XOR DI(945) XOR DI(582) XOR DI(863) XOR DI(441) XOR DI(791) XOR DI(971) XOR DI(760) XOR DI(158) XOR DI(643) XOR DI(0) XOR DI(363) XOR DI(709) XOR DI(99) XOR DI(128) XOR DI(454) XOR DI(252) XOR DI(742) XOR DI(875) XOR DI(882) XOR DI(245) XOR DI(317) XOR DI(192) XOR DI(344) XOR DI(847) XOR DI(691) XOR DI(250) XOR DI(776) XOR DI(803) XOR DI(716) XOR DI(597) XOR DI(339) XOR DI(805) XOR DI(200) XOR DI(870) XOR DI(233) XOR DI(309) XOR DI(109) XOR DI(946) XOR DI(361) XOR DI(194) XOR DI(479) XOR DI(1019) XOR DI(568) XOR DI(86) XOR DI(869) XOR DI(178) XOR DI(576) XOR DI(698) XOR DI(838) XOR DI(262) XOR DI(100) XOR DI(756) XOR DI(893) XOR DI(433) XOR DI(752) XOR DI(818) XOR DI(53) XOR DI(620) XOR DI(914) XOR DI(662) XOR DI(884) XOR DI(446) XOR DI(244) XOR DI(639) XOR DI(284) XOR DI(425) XOR DI(499) XOR DI(76) XOR DI(36) XOR DI(858) XOR DI(35) XOR DI(966) XOR DI(485) XOR DI(790) XOR DI(777) XOR DI(715) XOR DI(741) XOR DI(475) XOR DI(877) XOR DI(20) XOR DI(66) XOR DI(953) XOR DI(157) XOR DI(201) XOR DI(434) XOR DI(60) XOR DI(983) XOR DI(9) XOR DI(110) XOR DI(667) XOR DI(947) XOR DI(362) XOR DI(525) XOR DI(621) XOR DI(948) XOR DI(859) XOR DI(526) XOR DI(1020) XOR DI(767) XOR DI(278) XOR DI(866) XOR DI(307) XOR DI(570) XOR DI(977) XOR DI(557) XOR DI(51) XOR DI(687) XOR DI(871) XOR DI(91) XOR DI(331) XOR DI(763) XOR DI(47) XOR DI(190) XOR DI(839) XOR DI(560) XOR DI(964) XOR DI(180) XOR DI(550) XOR DI(954) XOR DI(151) XOR DI(161) XOR DI(646) XOR DI(700) XOR DI(3) XOR DI(366) XOR DI(911) XOR DI(382) XOR DI(496) XOR DI(588) XOR DI(798) XOR DI(259) XOR DI(224) XOR DI(634) XOR DI(6) XOR DI(712) XOR DI(131) XOR DI(1012) XOR DI(765) XOR DI(435) XOR DI(369) XOR DI(785) XOR DI(622) XOR DI(520) XOR DI(916) XOR DI(255) XOR DI(426) XOR DI(613) XOR DI(246) XOR DI(439) XOR DI(656) XOR DI(248) XOR DI(606) XOR DI(418) XOR DI(320) XOR DI(545) XOR DI(422) XOR DI(770) XOR DI(734) XOR DI(222) XOR DI(13) XOR DI(286) XOR DI(30) XOR DI(398) XOR DI(333) XOR DI(195) XOR DI(761) XOR DI(860) XOR DI(81) XOR DI(83) XOR DI(788) XOR DI(918) XOR DI(409) XOR DI(293) XOR DI(988) XOR DI(850) XOR DI(823) XOR DI(572) XOR DI(115) XOR DI(487) XOR DI(694) XOR DI(972) XOR DI(990) XOR DI(376) XOR DI(490) XOR DI(218) XOR DI(536) XOR DI(1006) XOR DI(748) XOR DI(743) XOR DI(739) XOR DI(442) XOR DI(240) XOR DI(231) XOR DI(719) XOR DI(396) XOR DI(650) XOR DI(600) XOR DI(314) XOR DI(22) XOR DI(903) XOR DI(539) XOR DI(405) XOR DI(659) XOR DI(280) XOR DI(392) XOR DI(327) XOR DI(297) XOR DI(608) XOR DI(935) XOR DI(72) XOR DI(266) XOR DI(139) XOR DI(407) XOR DI(808) XOR DI(508) XOR DI(203) XOR DI(471) XOR DI(873) XOR DI(644) XOR DI(236) XOR DI(62) XOR DI(985) XOR DI(722) XOR DI(1) XOR DI(274) XOR DI(386) XOR DI(176) XOR DI(500) XOR DI(461) XOR DI(26) XOR DI(669) XOR DI(143) XOR DI(364) XOR DI(153) XOR DI(197) XOR DI(380) XOR DI(663) XOR DI(943) XOR DI(855) XOR DI(482) XOR DI(129) XOR DI(1022) XOR DI(268) XOR DI(768) XOR DI(775) XOR DI(905) XOR DI(45) XOR DI(867) XOR DI(706) XOR DI(88) XOR DI(379) XOR DI(336) XOR DI(329) XOR DI(796) XOR DI(308) XOR DI(184) XOR DI(978) XOR DI(558) XOR DI(89) XOR DI(939) XOR DI(49) XOR DI(90) XOR DI(872) XOR DI(92) XOR DI(795) XOR DI(837) XOR DI(68) XOR DI(764) XOR DI(611) XOR DI(191) XOR DI(300) XOR DI(467) XOR DI(995) XOR DI(857) XOR DI(561) XOR DI(958) XOR DI(955) XOR DI(357) XOR DI(579) XOR DI(122) XOR DI(162) XOR DI(220) XOR DI(239) XOR DI(701) XOR DI(909) XOR DI(841) XOR DI(797) XOR DI(530) XOR DI(383) XOR DI(926) XOR DI(497) XOR DI(635) XOR DI(7) XOR DI(265) XOR DI(543) XOR DI(940) XOR DI(355) XOR DI(928) XOR DI(674) XOR DI(1013) XOR DI(759) XOR DI(766) XOR DI(786) XOR DI(724) XOR DI(291) XOR DI(172) XOR DI(821) XOR DI(542) XOR DI(230) XOR DI(56) XOR DI(623) XOR DI(216) XOR DI(123) XOR DI(750) XOR DI(746) XOR DI(533) XOR DI(614) XOR DI(737) XOR DI(440) XOR DI(238) XOR DI(728) XOR DI(813) XOR DI(888) XOR DI(403) XOR DI(633) XOR DI(886) XOR DI(657) XOR DI(504) XOR DI(465) XOR DI(852) XOR DI(321) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(960) XOR DI(546) XOR DI(423) XOR DI(147) XOR DI(686) XOR DI(897) XOR DI(412) XOR DI(711) XOR DI(642) XOR DI(895) XOR DI(666) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(811) XOR DI(865) XOR DI(283) XOR DI(544) XOR DI(661) XOR DI(941) XOR DI(145) XOR DI(196) XOR DI(615) XOR DI(853) XOR DI(133) XOR DI(474) XOR DI(502) XOR DI(762) XOR DI(79) XOR DI(861) XOR DI(82) XOR DI(323) XOR DI(38) XOR DI(302) XOR DI(565) XOR DI(46) XOR DI(164) XOR DI(84) XOR DI(789) XOR DI(969) XOR DI(758) XOR DI(727) XOR DI(605) XOR DI(294) XOR DI(989) XOR DI(555) XOR DI(175) XOR DI(824) XOR DI(351) XOR DI(573) XOR DI(116) XOR DI(156) XOR DI(214) XOR DI(695) XOR DI(973) XOR DI(991) XOR DI(377) XOR DI(920) XOR DI(537) XOR DI(922) XOR DI(430) XOR DI(749) XOR DI(718) XOR DI(826) XOR DI(515) XOR DI(744) XOR DI(443) XOR DI(215) XOR DI(241) XOR DI(731) XOR DI(478) XOR DI(807) XOR DI(720) XOR DI(627) XOR DI(243) XOR DI(601) XOR DI(413) XOR DI(498) XOR DI(23) XOR DI(149) XOR DI(904) XOR DI(417) XOR DI(992) XOR DI(729) XOR DI(406) XOR DI(217) XOR DI(705) XOR DI(636) XOR DI(8) XOR DI(281) XOR DI(393) XOR DI(328) XOR DI(298) XOR DI(119) XOR DI(350) XOR DI(183) XOR DI(609) XOR DI(936) XOR DI(267) XOR DI(559) XOR DI(404) XOR DI(963) XOR DI(599) XOR DI(956) XOR DI(140) XOR DI(150) XOR DI(208) XOR DI(408) XOR DI(371) XOR DI(213) XOR DI(531) XOR DI(204) XOR DI(270) XOR DI(437) XOR DI(209) XOR DI(235) XOR DI(645) XOR DI(17) XOR DI(411) XOR DI(986) XOR DI(400) XOR DI(630) XOR DI(2) XOR DI(654) XOR DI(292) XOR DI(649) XOR DI(121) XOR DI(27) XOR DI(553) XOR DI(907) XOR DI(957) XOR DI(950) XOR DI(163) XOR DI(365) XOR DI(207) XOR DI(814) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(11) XOR DI(394) XOR DI(664) XOR DI(944) XOR DI(460) XOR DI(702) XOR DI(862) XOR DI(522) XOR DI(199) XOR DI(489) XOR DI(450) XOR DI(938) XOR DI(856) XOR DI(136) XOR DI(130) XOR DI(124) XOR DI(678) XOR DI(517) XOR DI(505) XOR DI(1011) XOR DI(1023);
   DO(24) <= DI(564) XOR DI(96) XOR DI(779) XOR DI(782) XOR DI(982) XOR DI(844) XOR DI(109) XOR DI(1000) XOR DI(800) XOR DI(592) XOR DI(638) XOR DI(943) XOR DI(1016) XOR DI(439) XOR DI(641) XOR DI(97) XOR DI(224) XOR DI(250) XOR DI(190) XOR DI(248) XOR DI(1001) XOR DI(774) XOR DI(226) XOR DI(801) XOR DI(595) XOR DI(930) XOR DI(593) XOR DI(803) XOR DI(307) XOR DI(980) XOR DI(107) XOR DI(359) XOR DI(770) XOR DI(836) XOR DI(669) XOR DI(781) XOR DI(51) XOR DI(882) XOR DI(881) XOR DI(847) XOR DI(890) XOR DI(656) XOR DI(74) XOR DI(34) XOR DI(846) XOR DI(626) XOR DI(344) XOR DI(1002) XOR DI(473) XOR DI(875) XOR DI(899) XOR DI(338) XOR DI(58) XOR DI(981) XOR DI(382) XOR DI(946) XOR DI(697) XOR DI(536) XOR DI(691) XOR DI(524) XOR DI(1018) XOR DI(583) XOR DI(772) XOR DI(864) XOR DI(442) XOR DI(376) XOR DI(333) XOR DI(305) XOR DI(792) XOR DI(834) XOR DI(972) XOR DI(761) XOR DI(608) XOR DI(178) XOR DI(548) XOR DI(952) XOR DI(576) XOR DI(159) XOR DI(644) XOR DI(1) XOR DI(364) XOR DI(257) XOR DI(222) XOR DI(710) XOR DI(262) XOR DI(100) XOR DI(129) XOR DI(671) XOR DI(433) XOR DI(455) XOR DI(53) XOR DI(620) XOR DI(914) XOR DI(253) XOR DI(743) XOR DI(876) XOR DI(810) XOR DI(883) XOR DI(246) XOR DI(318) XOR DI(26) XOR DI(892) XOR DI(255) XOR DI(331) XOR DI(193) XOR DI(345) XOR DI(848) XOR DI(552) XOR DI(485) XOR DI(692) XOR DI(251) XOR DI(777) XOR DI(715) XOR DI(741) XOR DI(804) XOR DI(717) XOR DI(648) XOR DI(598) XOR DI(20) XOR DI(901) XOR DI(30) XOR DI(340) XOR DI(806) XOR DI(817) XOR DI(201) XOR DI(388) XOR DI(871) XOR DI(234) XOR DI(310) XOR DI(110) XOR DI(459) XOR DI(947) XOR DI(362) XOR DI(195) XOR DI(453) XOR DI(457) XOR DI(480) XOR DI(508) XOR DI(1008) XOR DI(1020) XOR DI(277) XOR DI(86) XOR DI(794) XOR DI(182) XOR DI(569) XOR DI(87) XOR DI(870) XOR DI(572) XOR DI(66) XOR DI(855) XOR DI(966) XOR DI(179) XOR DI(577) XOR DI(446) XOR DI(734) XOR DI(699) XOR DI(977) XOR DI(839) XOR DI(104) XOR DI(683) XOR DI(171) XOR DI(263) XOR DI(101) XOR DI(757) XOR DI(894) XOR DI(434) XOR DI(297) XOR DI(753) XOR DI(722) XOR DI(819) XOR DI(54) XOR DI(621) XOR DI(915) XOR DI(663) XOR DI(748) XOR DI(885) XOR DI(425) XOR DI(280) XOR DI(447) XOR DI(510) XOR DI(245) XOR DI(482) XOR DI(13) XOR DI(153) XOR DI(135) XOR DI(640) XOR DI(285) XOR DI(588) XOR DI(426) XOR DI(143) XOR DI(187) XOR DI(500) XOR DI(77) XOR DI(37) XOR DI(859) XOR DI(36) XOR DI(563) XOR DI(680) XOR DI(967) XOR DI(756) XOR DI(114) XOR DI(486) XOR DI(971) XOR DI(677) XOR DI(918) XOR DI(791) XOR DI(778) XOR DI(716) XOR DI(742) XOR DI(274) XOR DI(476) XOR DI(878) XOR DI(317) XOR DI(496) XOR DI(21) XOR DI(67) XOR DI(415) XOR DI(6) XOR DI(16) XOR DI(326) XOR DI(71) XOR DI(954) XOR DI(167) XOR DI(138) XOR DI(206) XOR DI(369) XOR DI(118) XOR DI(422) XOR DI(158) XOR DI(202) XOR DI(435) XOR DI(233) XOR DI(470) XOR DI(61) XOR DI(984) XOR DI(398) XOR DI(0) XOR DI(652) XOR DI(10) XOR DI(320) XOR DI(111) XOR DI(668) XOR DI(948) XOR DI(161) XOR DI(617) XOR DI(363) XOR DI(335) XOR DI(429) XOR DI(464) XOR DI(526) XOR DI(392) XOR DI(622) XOR DI(314) XOR DI(949) XOR DI(860) XOR DI(514) XOR DI(527) XOR DI(128) XOR DI(1015) XOR DI(1021) XOR DI(575) XOR DI(999) XOR DI(41) XOR DI(768) XOR DI(45) XOR DI(279) XOR DI(867) XOR DI(587) XOR DI(833) XOR DI(994) XOR DI(44) XOR DI(308) XOR DI(571) XOR DI(978) XOR DI(558) XOR DI(52) XOR DI(49) XOR DI(170) XOR DI(354) XOR DI(688) XOR DI(872) XOR DI(92) XOR DI(925) XOR DI(332) XOR DI(764) XOR DI(48) XOR DI(191) XOR DI(300) XOR DI(840) XOR DI(995) XOR DI(561) XOR DI(965) XOR DI(181) XOR DI(830) XOR DI(551) XOR DI(955) XOR DI(152) XOR DI(357) XOR DI(162) XOR DI(220) XOR DI(736) XOR DI(647) XOR DI(494) XOR DI(65) XOR DI(701) XOR DI(632) XOR DI(4) XOR DI(841) XOR DI(106) XOR DI(685) XOR DI(367) XOR DI(912) XOR DI(420) XOR DI(530) XOR DI(383) XOR DI(926) XOR DI(497) XOR DI(589) XOR DI(799) XOR DI(260) XOR DI(225) XOR DI(635) XOR DI(7) XOR DI(976) XOR DI(713) XOR DI(355) XOR DI(928) XOR DI(132) XOR DI(1013) XOR DI(766) XOR DI(436) XOR DI(370) XOR DI(786) XOR DI(755) XOR DI(724) XOR DI(821) XOR DI(542) XOR DI(623) XOR DI(832) XOR DI(521) XOR DI(917) XOR DI(704) XOR DI(256) XOR DI(427) XOR DI(449) XOR DI(533) XOR DI(614) XOR DI(512) XOR DI(247) XOR DI(737) XOR DI(440) XOR DI(212) XOR DI(238) XOR DI(484) XOR DI(888) XOR DI(726) XOR DI(633) XOR DI(657) XOR DI(15) XOR DI(249) XOR DI(607) XOR DI(419) XOR DI(493) XOR DI(70) XOR DI(852) XOR DI(321) XOR DI(155) XOR DI(546) XOR DI(423) XOR DI(147) XOR DI(686) XOR DI(897) XOR DI(998) XOR DI(771) XOR DI(735) XOR DI(223) XOR DI(469) XOR DI(14) XOR DI(174) XOR DI(666) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(399) XOR DI(334) XOR DI(428) XOR DI(304) XOR DI(283) XOR DI(661) XOR DI(145) XOR DI(189) XOR DI(196) XOR DI(513) XOR DI(133) XOR DI(502) XOR DI(762) XOR DI(861) XOR DI(82) XOR DI(323) XOR DI(302) XOR DI(43) XOR DI(84) XOR DI(682) XOR DI(789) XOR DI(919) XOR DI(831) XOR DI(410) XOR DI(969) XOR DI(727) XOR DI(605) XOR DI(42) XOR DI(294) XOR DI(989) XOR DI(851) XOR DI(175) XOR DI(824) XOR DI(432) XOR DI(573) XOR DI(116) XOR DI(156) XOR DI(488) XOR DI(695) XOR DI(973) XOR DI(991) XOR DI(377) XOR DI(920) XOR DI(491) XOR DI(219) XOR DI(537) XOR DI(349) XOR DI(126) XOR DI(1007) XOR DI(749) XOR DI(826) XOR DI(368) XOR DI(744) XOR DI(421) XOR DI(740) XOR DI(276) XOR DI(443) XOR DI(241) XOR DI(232) XOR DI(720) XOR DI(397) XOR DI(880) XOR DI(651) XOR DI(601) XOR DI(64) XOR DI(315) XOR DI(23) XOR DI(149) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(417) XOR DI(406) XOR DI(463) XOR DI(705) XOR DI(660) XOR DI(281) XOR DI(25) XOR DI(393) XOR DI(328) XOR DI(298) XOR DI(350) XOR DI(609) XOR DI(936) XOR DI(127) XOR DI(73) XOR DI(267) XOR DI(40) XOR DI(676) XOR DI(913) XOR DI(963) XOR DI(140) XOR DI(625) XOR DI(689) XOR DI(408) XOR DI(371) XOR DI(213) XOR DI(809) XOR DI(509) XOR DI(204) XOR DI(437) XOR DI(472) XOR DI(714) XOR DI(874) XOR DI(645) XOR DI(237) XOR DI(492) XOR DI(63) XOR DI(411) XOR DI(986) XOR DI(723) XOR DI(400) XOR DI(211) XOR DI(2) XOR DI(275) XOR DI(19) XOR DI(387) XOR DI(177) XOR DI(501) XOR DI(121) XOR DI(462) XOR DI(27) XOR DI(261) XOR DI(670) XOR DI(907) XOR DI(619) XOR DI(144) XOR DI(365) XOR DI(154) XOR DI(198) XOR DI(381) XOR DI(316) XOR DI(495) XOR DI(664) XOR DI(944) XOR DI(5) XOR DI(522) XOR DI(199) XOR DI(375) XOR DI(489) XOR DI(450) XOR DI(541) XOR DI(856) XOR DI(483) XOR DI(535) XOR DI(690) XOR DI(529) XOR DI(130) XOR DI(517) XOR DI(1023);
   DO(25) <= DI(580) XOR DI(565) XOR DI(475) XOR DI(97) XOR DI(780) XOR DI(880) XOR DI(76) XOR DI(783) XOR DI(983) XOR DI(845) XOR DI(110) XOR DI(1001) XOR DI(801) XOR DI(930) XOR DI(593) XOR DI(337) XOR DI(639) XOR DI(57) XOR DI(980) XOR DI(944) XOR DI(359) XOR DI(1017) XOR DI(440) XOR DI(566) XOR DI(759) XOR DI(642) XOR DI(98) XOR DI(781) XOR DI(453) XOR DI(225) XOR DI(251) XOR DI(244) XOR DI(70) XOR DI(637) XOR DI(191) XOR DI(469) XOR DI(249) XOR DI(1002) XOR DI(775) XOR DI(227) XOR DI(802) XOR DI(596) XOR DI(931) XOR DI(594) XOR DI(338) XOR DI(804) XOR DI(869) XOR DI(308) XOR DI(981) XOR DI(108) XOR DI(548) XOR DI(360) XOR DI(137) XOR DI(1018) XOR DI(771) XOR DI(901) XOR DI(304) XOR DI(826) XOR DI(951) XOR DI(575) XOR DI(697) XOR DI(837) XOR DI(670) XOR DI(755) XOR DI(892) XOR DI(432) XOR DI(782) XOR DI(751) XOR DI(52) XOR DI(619) XOR DI(517) XOR DI(883) XOR DI(882) XOR DI(848) XOR DI(638) XOR DI(891) XOR DI(283) XOR DI(657) XOR DI(75) XOR DI(35) XOR DI(34) XOR DI(344) XOR DI(847) XOR DI(627) XOR DI(345) XOR DI(1003) XOR DI(776) XOR DI(474) XOR DI(876) XOR DI(19) XOR DI(900) XOR DI(952) XOR DI(339) XOR DI(816) XOR DI(59) XOR DI(982) XOR DI(383) XOR DI(109) XOR DI(666) XOR DI(524) XOR DI(947) XOR DI(698) XOR DI(858) XOR DI(537) XOR DI(692) XOR DI(525) XOR DI(1019) XOR DI(584) XOR DI(773) XOR DI(865) XOR DI(443) XOR DI(86) XOR DI(377) XOR DI(334) XOR DI(306) XOR DI(976) XOR DI(556) XOR DI(90) XOR DI(793) XOR DI(835) XOR DI(330) XOR DI(414) XOR DI(973) XOR DI(762) XOR DI(609) XOR DI(189) XOR DI(838) XOR DI(963) XOR DI(179) XOR DI(549) XOR DI(953) XOR DI(577) XOR DI(446) XOR DI(160) XOR DI(645) XOR DI(2) XOR DI(184) XOR DI(907) XOR DI(365) XOR DI(479) XOR DI(910) XOR DI(587) XOR DI(797) XOR DI(258) XOR DI(223) XOR DI(711) XOR DI(263) XOR DI(101) XOR DI(130) XOR DI(672) XOR DI(434) XOR DI(456) XOR DI(170) XOR DI(54) XOR DI(621) XOR DI(915) XOR DI(254) XOR DI(425) XOR DI(744) XOR DI(612) XOR DI(877) XOR DI(811) XOR DI(884) XOR DI(655) XOR DI(247) XOR DI(605) XOR DI(323) XOR DI(417) XOR DI(319) XOR DI(27) XOR DI(958) XOR DI(544) XOR DI(106) XOR DI(709) XOR DI(12) XOR DI(893) XOR DI(256) XOR DI(332) XOR DI(863) XOR DI(194) XOR DI(679) XOR DI(760) XOR DI(271) XOR DI(80) XOR DI(563) XOR DI(346) XOR DI(292) XOR DI(849) XOR DI(553) XOR DI(114) XOR DI(486) XOR DI(693) XOR DI(971) XOR DI(375) XOR DI(252) XOR DI(217) XOR DI(535) XOR DI(778) XOR DI(747) XOR DI(716) XOR DI(164) XOR DI(742) XOR DI(729) XOR DI(805) XOR DI(718) XOR DI(395) XOR DI(625) XOR DI(649) XOR DI(599) XOR DI(21) XOR DI(902) XOR DI(404) XOR DI(326) XOR DI(505) XOR DI(31) XOR DI(167) XOR DI(138) XOR DI(341) XOR DI(807) XOR DI(818) XOR DI(202) XOR DI(389) XOR DI(872) XOR DI(643) XOR DI(235) XOR DI(311) XOR DI(628) XOR DI(0) XOR DI(111) XOR DI(499) XOR DI(460) XOR DI(25) XOR DI(948) XOR DI(363) XOR DI(196) XOR DI(9) XOR DI(454) XOR DI(942) XOR DI(458) XOR DI(616) XOR DI(854) XOR DI(481) XOR DI(682) XOR DI(676) XOR DI(509) XOR DI(1009) XOR DI(1015) XOR DI(1021) XOR DI(998) XOR DI(40) XOR DI(352) XOR DI(278) XOR DI(866) XOR DI(300) XOR DI(87) XOR DI(993) XOR DI(795) XOR DI(183) XOR DI(570) XOR DI(88) XOR DI(89) XOR DI(923) XOR DI(871) XOR DI(91) XOR DI(573) XOR DI(794) XOR DI(836) XOR DI(67) XOR DI(331) XOR DI(415) XOR DI(732) XOR DI(47) XOR DI(104) XOR DI(466) XOR DI(994) XOR DI(856) XOR DI(560) XOR DI(967) XOR DI(180) XOR DI(957) XOR DI(151) XOR DI(578) XOR DI(121) XOR DI(447) XOR DI(161) XOR DI(735) XOR DI(700) XOR DI(631) XOR DI(185) XOR DI(978) XOR DI(840) XOR DI(105) XOR DI(684) XOR DI(911) XOR DI(796) XOR DI(529) XOR DI(172) XOR DI(925) XOR DI(798) XOR DI(259) XOR DI(302) XOR DI(712) XOR DI(264) XOR DI(102) XOR DI(939) XOR DI(354) XOR DI(187) XOR DI(1012) XOR DI(758) XOR DI(895) XOR DI(435) XOR DI(298) XOR DI(754) XOR DI(723) XOR DI(457) XOR DI(820) XOR DI(55) XOR DI(622) XOR DI(357) XOR DI(916) XOR DI(215) XOR DI(703) XOR DI(255) XOR DI(664) XOR DI(749) XOR DI(886) XOR DI(426) XOR DI(281) XOR DI(448) XOR DI(532) XOR DI(511) XOR DI(246) XOR DI(439) XOR DI(211) XOR DI(483) XOR DI(812) XOR DI(887) XOR DI(632) XOR DI(656) XOR DI(14) XOR DI(69) XOR DI(320) XOR DI(154) XOR DI(821) XOR DI(959) XOR DI(545) XOR DI(136) XOR DI(685) XOR DI(896) XOR DI(734) XOR DI(222) XOR DI(468) XOR DI(641) XOR DI(13) XOR DI(173) XOR DI(286) XOR DI(30) XOR DI(589) XOR DI(427) XOR DI(940) XOR DI(124) XOR DI(144) XOR DI(188) XOR DI(941) XOR DI(512) XOR DI(928) XOR DI(680) XOR DI(501) XOR DI(78) XOR DI(38) XOR DI(860) XOR DI(37) XOR DI(564) XOR DI(681) XOR DI(830) XOR DI(968) XOR DI(757) XOR DI(726) XOR DI(293) XOR DI(554) XOR DI(961) XOR DI(174) XOR DI(823) XOR DI(431) XOR DI(115) XOR DI(487) XOR DI(972) XOR DI(678) XOR DI(413) XOR DI(919) XOR DI(792) XOR DI(218) XOR DI(969) XOR DI(125) XOR DI(779) XOR DI(748) XOR DI(717) XOR DI(165) XOR DI(814) XOR DI(209) XOR DI(743) XOR DI(275) XOR DI(240) XOR DI(730) XOR DI(231) XOR DI(477) XOR DI(719) XOR DI(879) XOR DI(650) XOR DI(600) XOR DI(318) XOR DI(497) XOR DI(314) XOR DI(22) XOR DI(68) XOR DI(815) XOR DI(416) XOR DI(890) XOR DI(405) XOR DI(216) XOR DI(704) XOR DI(7) XOR DI(888) XOR DI(17) XOR DI(392) XOR DI(327) XOR DI(297) XOR DI(118) XOR DI(349) XOR DI(506) XOR DI(126) XOR DI(467) XOR DI(72) XOR DI(266) XOR DI(39) XOR DI(675) XOR DI(955) XOR DI(168) XOR DI(139) XOR DI(149) XOR DI(207) XOR DI(899) XOR DI(370) XOR DI(119) XOR DI(423) XOR DI(159) XOR DI(808) XOR DI(508) XOR DI(203) XOR DI(269) XOR DI(436) XOR DI(208) XOR DI(234) XOR DI(471) XOR DI(236) XOR DI(62) XOR DI(897) XOR DI(533) XOR DI(985) XOR DI(722) XOR DI(399) XOR DI(210) XOR DI(1) XOR DI(653) XOR DI(11) XOR DI(274) XOR DI(18) XOR DI(321) XOR DI(112) XOR DI(120) XOR DI(461) XOR DI(669) XOR DI(906) XOR DI(949) XOR DI(162) XOR DI(618) XOR DI(143) XOR DI(364) XOR DI(206) XOR DI(336) XOR DI(430) XOR DI(465) XOR DI(707) XOR DI(527) XOR DI(393) XOR DI(623) XOR DI(380) XOR DI(315) XOR DI(950) XOR DI(943) XOR DI(147) XOR DI(459) XOR DI(861) XOR DI(617) XOR DI(449) XOR DI(855) XOR DI(515) XOR DI(482) XOR DI(135) XOR DI(528) XOR DI(129) XOR DI(123) XOR DI(516) XOR DI(1016) XOR DI(1022);
   DO(26) <= DI(581) XOR DI(566) XOR DI(476) XOR DI(98) XOR DI(781) XOR DI(881) XOR DI(77) XOR DI(784) XOR DI(984) XOR DI(846) XOR DI(111) XOR DI(1002) XOR DI(802) XOR DI(931) XOR DI(594) XOR DI(338) XOR DI(640) XOR DI(58) XOR DI(981) XOR DI(945) XOR DI(360) XOR DI(1018) XOR DI(441) XOR DI(567) XOR DI(760) XOR DI(643) XOR DI(99) XOR DI(782) XOR DI(454) XOR DI(226) XOR DI(252) XOR DI(245) XOR DI(71) XOR DI(638) XOR DI(192) XOR DI(470) XOR DI(250) XOR DI(1003) XOR DI(776) XOR DI(228) XOR DI(803) XOR DI(597) XOR DI(932) XOR DI(595) XOR DI(339) XOR DI(805) XOR DI(870) XOR DI(309) XOR DI(982) XOR DI(109) XOR DI(549) XOR DI(361) XOR DI(138) XOR DI(1019) XOR DI(772) XOR DI(902) XOR DI(305) XOR DI(827) XOR DI(952) XOR DI(576) XOR DI(698) XOR DI(838) XOR DI(671) XOR DI(756) XOR DI(893) XOR DI(433) XOR DI(783) XOR DI(752) XOR DI(53) XOR DI(620) XOR DI(518) XOR DI(884) XOR DI(883) XOR DI(849) XOR DI(639) XOR DI(892) XOR DI(284) XOR DI(658) XOR DI(76) XOR DI(36) XOR DI(35) XOR DI(345) XOR DI(848) XOR DI(628) XOR DI(346) XOR DI(1004) XOR DI(777) XOR DI(475) XOR DI(877) XOR DI(20) XOR DI(901) XOR DI(953) XOR DI(340) XOR DI(817) XOR DI(60) XOR DI(983) XOR DI(384) XOR DI(110) XOR DI(667) XOR DI(525) XOR DI(948) XOR DI(699) XOR DI(859) XOR DI(538) XOR DI(693) XOR DI(526) XOR DI(1020) XOR DI(585) XOR DI(774) XOR DI(866) XOR DI(444) XOR DI(87) XOR DI(378) XOR DI(335) XOR DI(307) XOR DI(977) XOR DI(557) XOR DI(91) XOR DI(794) XOR DI(836) XOR DI(331) XOR DI(415) XOR DI(974) XOR DI(763) XOR DI(610) XOR DI(190) XOR DI(839) XOR DI(964) XOR DI(180) XOR DI(550) XOR DI(954) XOR DI(578) XOR DI(447) XOR DI(161) XOR DI(646) XOR DI(3) XOR DI(185) XOR DI(908) XOR DI(366) XOR DI(480) XOR DI(911) XOR DI(588) XOR DI(798) XOR DI(259) XOR DI(224) XOR DI(712) XOR DI(264) XOR DI(102) XOR DI(131) XOR DI(673) XOR DI(435) XOR DI(457) XOR DI(171) XOR DI(55) XOR DI(622) XOR DI(916) XOR DI(255) XOR DI(426) XOR DI(745) XOR DI(613) XOR DI(878) XOR DI(812) XOR DI(885) XOR DI(656) XOR DI(248) XOR DI(606) XOR DI(324) XOR DI(418) XOR DI(320) XOR DI(28) XOR DI(959) XOR DI(545) XOR DI(107) XOR DI(710) XOR DI(13) XOR DI(894) XOR DI(257) XOR DI(333) XOR DI(864) XOR DI(195) XOR DI(680) XOR DI(761) XOR DI(272) XOR DI(81) XOR DI(564) XOR DI(347) XOR DI(293) XOR DI(850) XOR DI(554) XOR DI(115) XOR DI(487) XOR DI(694) XOR DI(972) XOR DI(376) XOR DI(253) XOR DI(218) XOR DI(536) XOR DI(779) XOR DI(748) XOR DI(717) XOR DI(165) XOR DI(743) XOR DI(730) XOR DI(806) XOR DI(719) XOR DI(396) XOR DI(626) XOR DI(650) XOR DI(600) XOR DI(22) XOR DI(903) XOR DI(405) XOR DI(327) XOR DI(506) XOR DI(32) XOR DI(168) XOR DI(139) XOR DI(342) XOR DI(808) XOR DI(819) XOR DI(203) XOR DI(390) XOR DI(873) XOR DI(644) XOR DI(236) XOR DI(312) XOR DI(629) XOR DI(1) XOR DI(112) XOR DI(500) XOR DI(461) XOR DI(26) XOR DI(949) XOR DI(364) XOR DI(197) XOR DI(10) XOR DI(455) XOR DI(943) XOR DI(459) XOR DI(617) XOR DI(855) XOR DI(482) XOR DI(683) XOR DI(677) XOR DI(510) XOR DI(1010) XOR DI(1016) XOR DI(1022) XOR DI(999) XOR DI(41) XOR DI(353) XOR DI(279) XOR DI(867) XOR DI(301) XOR DI(88) XOR DI(994) XOR DI(796) XOR DI(184) XOR DI(571) XOR DI(89) XOR DI(90) XOR DI(924) XOR DI(872) XOR DI(92) XOR DI(574) XOR DI(795) XOR DI(837) XOR DI(68) XOR DI(332) XOR DI(416) XOR DI(733) XOR DI(48) XOR DI(105) XOR DI(467) XOR DI(995) XOR DI(857) XOR DI(561) XOR DI(968) XOR DI(181) XOR DI(958) XOR DI(152) XOR DI(579) XOR DI(122) XOR DI(448) XOR DI(162) XOR DI(736) XOR DI(701) XOR DI(632) XOR DI(186) XOR DI(979) XOR DI(841) XOR DI(106) XOR DI(685) XOR DI(912) XOR DI(797) XOR DI(530) XOR DI(173) XOR DI(926) XOR DI(799) XOR DI(260) XOR DI(303) XOR DI(713) XOR DI(265) XOR DI(103) XOR DI(940) XOR DI(355) XOR DI(188) XOR DI(1013) XOR DI(759) XOR DI(896) XOR DI(436) XOR DI(299) XOR DI(755) XOR DI(724) XOR DI(458) XOR DI(821) XOR DI(56) XOR DI(623) XOR DI(358) XOR DI(917) XOR DI(216) XOR DI(704) XOR DI(256) XOR DI(665) XOR DI(750) XOR DI(887) XOR DI(427) XOR DI(282) XOR DI(449) XOR DI(533) XOR DI(512) XOR DI(247) XOR DI(440) XOR DI(212) XOR DI(484) XOR DI(813) XOR DI(888) XOR DI(633) XOR DI(657) XOR DI(15) XOR DI(70) XOR DI(321) XOR DI(155) XOR DI(822) XOR DI(960) XOR DI(546) XOR DI(137) XOR DI(686) XOR DI(897) XOR DI(735) XOR DI(223) XOR DI(469) XOR DI(642) XOR DI(14) XOR DI(174) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(428) XOR DI(941) XOR DI(125) XOR DI(145) XOR DI(189) XOR DI(942) XOR DI(513) XOR DI(929) XOR DI(681) XOR DI(502) XOR DI(79) XOR DI(39) XOR DI(861) XOR DI(38) XOR DI(565) XOR DI(682) XOR DI(831) XOR DI(969) XOR DI(758) XOR DI(727) XOR DI(294) XOR DI(555) XOR DI(962) XOR DI(175) XOR DI(824) XOR DI(432) XOR DI(116) XOR DI(488) XOR DI(973) XOR DI(679) XOR DI(414) XOR DI(920) XOR DI(793) XOR DI(219) XOR DI(970) XOR DI(126) XOR DI(780) XOR DI(749) XOR DI(718) XOR DI(166) XOR DI(815) XOR DI(210) XOR DI(744) XOR DI(276) XOR DI(241) XOR DI(731) XOR DI(232) XOR DI(478) XOR DI(720) XOR DI(880) XOR DI(651) XOR DI(601) XOR DI(319) XOR DI(498) XOR DI(315) XOR DI(23) XOR DI(69) XOR DI(816) XOR DI(417) XOR DI(891) XOR DI(406) XOR DI(217) XOR DI(705) XOR DI(8) XOR DI(889) XOR DI(18) XOR DI(393) XOR DI(328) XOR DI(298) XOR DI(119) XOR DI(350) XOR DI(507) XOR DI(127) XOR DI(468) XOR DI(73) XOR DI(267) XOR DI(40) XOR DI(676) XOR DI(956) XOR DI(169) XOR DI(140) XOR DI(150) XOR DI(208) XOR DI(900) XOR DI(371) XOR DI(120) XOR DI(424) XOR DI(160) XOR DI(809) XOR DI(509) XOR DI(204) XOR DI(270) XOR DI(437) XOR DI(209) XOR DI(235) XOR DI(472) XOR DI(237) XOR DI(63) XOR DI(898) XOR DI(534) XOR DI(986) XOR DI(723) XOR DI(400) XOR DI(211) XOR DI(2) XOR DI(654) XOR DI(12) XOR DI(275) XOR DI(19) XOR DI(322) XOR DI(113) XOR DI(121) XOR DI(462) XOR DI(670) XOR DI(907) XOR DI(950) XOR DI(163) XOR DI(619) XOR DI(144) XOR DI(365) XOR DI(207) XOR DI(337) XOR DI(431) XOR DI(466) XOR DI(708) XOR DI(528) XOR DI(394) XOR DI(624) XOR DI(381) XOR DI(316) XOR DI(951) XOR DI(944) XOR DI(148) XOR DI(460) XOR DI(862) XOR DI(618) XOR DI(450) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(136) XOR DI(529) XOR DI(130) XOR DI(124) XOR DI(517) XOR DI(1017) XOR DI(1023);
   DO(27) <= DI(582) XOR DI(567) XOR DI(554) XOR DI(836) XOR DI(964) XOR DI(444) XOR DI(600) XOR DI(697) XOR DI(477) XOR DI(99) XOR DI(782) XOR DI(226) XOR DI(610) XOR DI(875) XOR DI(882) XOR DI(767) XOR DI(707) XOR DI(638) XOR DI(192) XOR DI(269) XOR DI(78) XOR DI(34) XOR DI(344) XOR DI(785) XOR DI(985) XOR DI(847) XOR DI(112) XOR DI(691) XOR DI(250) XOR DI(1003) XOR DI(776) XOR DI(439) XOR DI(803) XOR DI(536) XOR DI(656) XOR DI(324) XOR DI(932) XOR DI(595) XOR DI(165) XOR DI(339) XOR DI(200) XOR DI(231) XOR DI(641) XOR DI(309) XOR DI(59) XOR DI(982) XOR DI(626) XOR DI(650) XOR DI(109) XOR DI(946) XOR DI(361) XOR DI(524) XOR DI(1019) XOR DI(765) XOR DI(772) XOR DI(442) XOR DI(376) XOR DI(305) XOR DI(568) XOR DI(869) XOR DI(834) XOR DI(761) XOR DI(730) XOR DI(608) XOR DI(178) XOR DI(548) XOR DI(576) XOR DI(644) XOR DI(380) XOR DI(222) XOR DI(262) XOR DI(100) XOR DI(763) XOR DI(783) XOR DI(455) XOR DI(227) XOR DI(53) XOR DI(914) XOR DI(253) XOR DI(244) XOR DI(246) XOR DI(26) XOR DI(72) XOR DI(639) XOR DI(255) XOR DI(284) XOR DI(28) XOR DI(331) XOR DI(808) XOR DI(193) XOR DI(471) XOR DI(76) XOR DI(552) XOR DI(790) XOR DI(251) XOR DI(1004) XOR DI(777) XOR DI(715) XOR DI(741) XOR DI(229) XOR DI(475) XOR DI(804) XOR DI(648) XOR DI(240) XOR DI(598) XOR DI(606) XOR DI(933) XOR DI(30) XOR DI(293) XOR DI(596) XOR DI(405) XOR DI(340) XOR DI(157) XOR DI(806) XOR DI(506) XOR DI(388) XOR DI(871) XOR DI(310) XOR DI(983) XOR DI(384) XOR DI(646) XOR DI(110) XOR DI(550) XOR DI(667) XOR DI(362) XOR DI(378) XOR DI(453) XOR DI(457) XOR DI(139) XOR DI(1008) XOR DI(1020) XOR DI(773) XOR DI(903) XOR DI(83) XOR DI(86) XOR DI(306) XOR DI(50) XOR DI(937) XOR DI(47) XOR DI(352) XOR DI(923) XOR DI(66) XOR DI(855) XOR DI(966) XOR DI(828) XOR DI(953) XOR DI(577) XOR DI(446) XOR DI(699) XOR DI(977) XOR DI(839) XOR DI(171) XOR DI(672) XOR DI(757) XOR DI(894) XOR DI(434) XOR DI(297) XOR DI(560) XOR DI(784) XOR DI(753) XOR DI(722) XOR DI(54) XOR DI(621) XOR DI(519) XOR DI(748) XOR DI(885) XOR DI(612) XOR DI(482) XOR DI(884) XOR DI(850) XOR DI(135) XOR DI(769) XOR DI(640) XOR DI(893) XOR DI(285) XOR DI(588) XOR DI(659) XOR DI(143) XOR DI(1012) XOR DI(77) XOR DI(37) XOR DI(36) XOR DI(563) XOR DI(346) XOR DI(787) XOR DI(849) XOR DI(629) XOR DI(347) XOR DI(1005) XOR DI(778) XOR DI(738) XOR DI(274) XOR DI(476) XOR DI(878) XOR DI(496) XOR DI(21) XOR DI(902) XOR DI(538) XOR DI(990) XOR DI(6) XOR DI(326) XOR DI(911) XOR DI(954) XOR DI(206) XOR DI(827) XOR DI(369) XOR DI(341) XOR DI(118) XOR DI(422) XOR DI(818) XOR DI(712) XOR DI(490) XOR DI(61) XOR DI(409) XOR DI(984) XOR DI(398) XOR DI(628) XOR DI(385) XOR DI(111) XOR DI(259) XOR DI(668) XOR DI(617) XOR DI(335) XOR DI(812) XOR DI(464) XOR DI(866) XOR DI(526) XOR DI(392) XOR DI(314) XOR DI(545) XOR DI(662) XOR DI(949) XOR DI(700) XOR DI(860) XOR DI(197) XOR DI(539) XOR DI(694) XOR DI(527) XOR DI(1015) XOR DI(1021) XOR DI(999) XOR DI(747) XOR DI(586) XOR DI(775) XOR DI(905) XOR DI(85) XOR DI(45) XOR DI(867) XOR DI(587) XOR DI(445) XOR DI(301) XOR DI(88) XOR DI(379) XOR DI(336) XOR DI(833) XOR DI(994) XOR DI(44) XOR DI(308) XOR DI(184) XOR DI(854) XOR DI(978) XOR DI(558) XOR DI(939) XOR DI(92) XOR DI(574) XOR DI(795) XOR DI(837) XOR DI(332) XOR DI(416) XOR DI(975) XOR DI(764) XOR DI(611) XOR DI(191) XOR DI(840) XOR DI(965) XOR DI(181) XOR DI(830) XOR DI(551) XOR DI(958) XOR DI(955) XOR DI(637) XOR DI(357) XOR DI(579) XOR DI(703) XOR DI(448) XOR DI(162) XOR DI(647) XOR DI(239) XOR DI(494) XOR DI(65) XOR DI(632) XOR DI(4) XOR DI(186) XOR DI(909) XOR DI(979) XOR DI(841) XOR DI(685) XOR DI(367) XOR DI(481) XOR DI(912) XOR DI(420) XOR DI(173) XOR DI(926) XOR DI(589) XOR DI(799) XOR DI(260) XOR DI(225) XOR DI(303) XOR DI(976) XOR DI(713) XOR DI(265) XOR DI(103) XOR DI(543) XOR DI(940) XOR DI(355) XOR DI(928) XOR DI(132) XOR DI(674) XOR DI(896) XOR DI(436) XOR DI(755) XOR DI(458) XOR DI(172) XOR DI(821) XOR DI(542) XOR DI(56) XOR DI(623) XOR DI(358) XOR DI(917) XOR DI(216) XOR DI(704) XOR DI(256) XOR DI(665) XOR DI(887) XOR DI(427) XOR DI(746) XOR DI(282) XOR DI(533) XOR DI(221) XOR DI(614) XOR DI(512) XOR DI(879) XOR DI(813) XOR DI(726) XOR DI(886) XOR DI(657) XOR DI(249) XOR DI(607) XOR DI(325) XOR DI(419) XOR DI(493) XOR DI(852) XOR DI(321) XOR DI(29) XOR DI(155) XOR DI(910) XOR DI(960) XOR DI(546) XOR DI(147) XOR DI(998) XOR DI(108) XOR DI(412) XOR DI(711) XOR DI(14) XOR DI(895) XOR DI(258) XOR DI(590) XOR DI(616) XOR DI(334) XOR DI(865) XOR DI(544) XOR DI(661) XOR DI(196) XOR DI(615) XOR DI(853) XOR DI(532) XOR DI(929) XOR DI(133) XOR DI(681) XOR DI(502) XOR DI(993) XOR DI(762) XOR DI(273) XOR DI(82) XOR DI(330) XOR DI(565) XOR DI(46) XOR DI(43) XOR DI(348) XOR DI(831) XOR DI(727) XOR DI(605) XOR DI(294) XOR DI(851) XOR DI(555) XOR DI(631) XOR DI(116) XOR DI(214) XOR DI(488) XOR DI(695) XOR DI(973) XOR DI(679) XOR DI(906) XOR DI(414) XOR DI(377) XOR DI(920) XOR DI(254) XOR DI(219) XOR DI(537) XOR DI(349) XOR DI(780) XOR DI(749) XOR DI(718) XOR DI(166) XOR DI(815) XOR DI(826) XOR DI(368) XOR DI(744) XOR DI(421) XOR DI(215) XOR DI(731) XOR DI(807) XOR DI(720) XOR DI(397) XOR DI(627) XOR DI(880) XOR DI(651) XOR DI(601) XOR DI(413) XOR DI(498) XOR DI(23) XOR DI(904) XOR DI(992) XOR DI(729) XOR DI(406) XOR DI(636) XOR DI(8) XOR DI(18) XOR DI(25) XOR DI(328) XOR DI(350) XOR DI(507) XOR DI(675) XOR DI(33) XOR DI(559) XOR DI(676) XOR DI(404) XOR DI(956) XOR DI(169) XOR DI(140) XOR DI(150) XOR DI(689) XOR DI(371) XOR DI(343) XOR DI(424) XOR DI(809) XOR DI(820) XOR DI(204) XOR DI(391) XOR DI(874) XOR DI(645) XOR DI(237) XOR DI(313) XOR DI(492) XOR DI(411) XOR DI(400) XOR DI(630) XOR DI(2) XOR DI(12) XOR DI(292) XOR DI(113) XOR DI(501) XOR DI(462) XOR DI(27) XOR DI(907) XOR DI(950) XOR DI(134) XOR DI(365) XOR DI(337) XOR DI(198) XOR DI(431) XOR DI(466) XOR DI(11) XOR DI(495) XOR DI(456) XOR DI(944) XOR DI(148) XOR DI(460) XOR DI(5) XOR DI(522) XOR DI(199) XOR DI(618) XOR DI(375) XOR DI(541) XOR DI(696) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(690) XOR DI(684) XOR DI(523) XOR DI(124) XOR DI(678) XOR DI(511) XOR DI(505) XOR DI(1011) XOR DI(1017) XOR DI(1023);
   DO(28) <= DI(583) XOR DI(772) XOR DI(276) XOR DI(85) XOR DI(305) XOR DI(568) XOR DI(555) XOR DI(49) XOR DI(869) XOR DI(65) XOR DI(837) XOR DI(965) XOR DI(751) XOR DI(178) XOR DI(548) XOR DI(952) XOR DI(576) XOR DI(445) XOR DI(601) XOR DI(698) XOR DI(478) XOR DI(262) XOR DI(100) XOR DI(671) XOR DI(433) XOR DI(783) XOR DI(288) XOR DI(227) XOR DI(53) XOR DI(620) XOR DI(518) XOR DI(371) XOR DI(914) XOR DI(424) XOR DI(611) XOR DI(244) XOR DI(876) XOR DI(400) XOR DI(883) XOR DI(768) XOR DI(708) XOR DI(639) XOR DI(892) XOR DI(284) XOR DI(862) XOR DI(193) XOR DI(759) XOR DI(76) XOR DI(270) XOR DI(858) XOR DI(79) XOR DI(35) XOR DI(562) XOR DI(345) XOR DI(786) XOR DI(755) XOR DI(986) XOR DI(848) XOR DI(113) XOR DI(485) XOR DI(692) XOR DI(970) XOR DI(790) XOR DI(251) XOR DI(1004) XOR DI(777) XOR DI(715) XOR DI(741) XOR DI(737) XOR DI(440) XOR DI(475) XOR DI(804) XOR DI(394) XOR DI(316) XOR DI(20) XOR DI(901) XOR DI(537) XOR DI(657) XOR DI(325) XOR DI(933) XOR DI(70) XOR DI(596) XOR DI(166) XOR DI(137) XOR DI(826) XOR DI(340) XOR DI(157) XOR DI(817) XOR DI(201) XOR DI(232) XOR DI(469) XOR DI(388) XOR DI(642) XOR DI(310) XOR DI(60) XOR DI(983) XOR DI(627) XOR DI(651) XOR DI(384) XOR DI(110) XOR DI(498) XOR DI(667) XOR DI(947) XOR DI(362) XOR DI(8) XOR DI(525) XOR DI(453) XOR DI(661) XOR DI(127) XOR DI(1008) XOR DI(1014) XOR DI(1020) XOR DI(766) XOR DI(773) XOR DI(277) XOR DI(443) XOR DI(377) XOR DI(306) XOR DI(569) XOR DI(50) XOR DI(870) XOR DI(90) XOR DI(835) XOR DI(330) XOR DI(762) XOR DI(731) XOR DI(609) XOR DI(189) XOR DI(963) XOR DI(179) XOR DI(549) XOR DI(150) XOR DI(577) XOR DI(645) XOR DI(184) XOR DI(479) XOR DI(381) XOR DI(797) XOR DI(223) XOR DI(263) XOR DI(101) XOR DI(764) XOR DI(784) XOR DI(456) XOR DI(228) XOR DI(54) XOR DI(915) XOR DI(254) XOR DI(245) XOR DI(438) XOR DI(655) XOR DI(247) XOR DI(605) XOR DI(323) XOR DI(27) XOR DI(73) XOR DI(958) XOR DI(769) XOR DI(106) XOR DI(221) XOR DI(709) XOR DI(640) XOR DI(256) XOR DI(285) XOR DI(29) XOR DI(332) XOR DI(809) XOR DI(863) XOR DI(194) XOR DI(472) XOR DI(760) XOR DI(77) XOR DI(271) XOR DI(80) XOR DI(563) XOR DI(787) XOR DI(292) XOR DI(987) XOR DI(553) XOR DI(971) XOR DI(833) XOR DI(375) XOR DI(791) XOR DI(252) XOR DI(535) XOR DI(920) XOR DI(1005) XOR DI(778) XOR DI(716) XOR DI(450) XOR DI(164) XOR DI(742) XOR DI(738) XOR DI(441) XOR DI(239) XOR DI(729) XOR DI(230) XOR DI(476) XOR DI(805) XOR DI(395) XOR DI(625) XOR DI(649) XOR DI(241) XOR DI(599) XOR DI(317) XOR DI(889) XOR DI(404) XOR DI(607) XOR DI(934) XOR DI(505) XOR DI(71) XOR DI(31) XOR DI(294) XOR DI(597) XOR DI(138) XOR DI(898) XOR DI(406) XOR DI(341) XOR DI(158) XOR DI(807) XOR DI(507) XOR DI(268) XOR DI(233) XOR DI(470) XOR DI(389) XOR DI(872) XOR DI(643) XOR DI(311) XOR DI(984) XOR DI(0) XOR DI(385) XOR DI(647) XOR DI(111) XOR DI(175) XOR DI(25) XOR DI(551) XOR DI(668) XOR DI(363) XOR DI(706) XOR DI(379) XOR DI(454) XOR DI(942) XOR DI(458) XOR DI(140) XOR DI(128) XOR DI(1009) XOR DI(1015) XOR DI(1021) XOR DI(574) XOR DI(998) XOR DI(40) XOR DI(352) XOR DI(767) XOR DI(774) XOR DI(904) XOR DI(84) XOR DI(444) XOR DI(300) XOR DI(87) XOR DI(43) XOR DI(307) XOR DI(51) XOR DI(938) XOR DI(48) XOR DI(923) XOR DI(353) XOR DI(687) XOR DI(91) XOR DI(794) XOR DI(924) XOR DI(836) XOR DI(67) XOR DI(610) XOR DI(190) XOR DI(299) XOR DI(466) XOR DI(856) XOR DI(967) XOR DI(964) XOR DI(829) XOR DI(954) XOR DI(636) XOR DI(578) XOR DI(702) XOR DI(121) XOR DI(447) XOR DI(161) XOR DI(64) XOR DI(700) XOR DI(978) XOR DI(840) XOR DI(996) XOR DI(529) XOR DI(382) XOR DI(172) XOR DI(925) XOR DI(798) XOR DI(224) XOR DI(634) XOR DI(939) XOR DI(354) XOR DI(131) XOR DI(673) XOR DI(758) XOR DI(895) XOR DI(435) XOR DI(298) XOR DI(561) XOR DI(785) XOR DI(754) XOR DI(723) XOR DI(171) XOR DI(541) XOR DI(55) XOR DI(622) XOR DI(357) XOR DI(520) XOR DI(703) XOR DI(122) XOR DI(749) XOR DI(886) XOR DI(532) XOR DI(613) XOR DI(736) XOR DI(439) XOR DI(211) XOR DI(483) XOR DI(812) XOR DI(725) XOR DI(885) XOR DI(656) XOR DI(248) XOR DI(324) XOR DI(418) XOR DI(464) XOR DI(492) XOR DI(69) XOR DI(851) XOR DI(320) XOR DI(74) XOR DI(136) XOR DI(146) XOR DI(770) XOR DI(107) XOR DI(734) XOR DI(411) XOR DI(468) XOR DI(641) XOR DI(894) XOR DI(926) XOR DI(665) XOR DI(286) XOR DI(589) XOR DI(303) XOR DI(282) XOR DI(660) XOR DI(124) XOR DI(355) XOR DI(144) XOR DI(531) XOR DI(928) XOR DI(473) XOR DI(1013) XOR DI(992) XOR DI(78) XOR DI(38) XOR DI(37) XOR DI(301) XOR DI(564) XOR DI(42) XOR DI(347) XOR DI(788) XOR DI(830) XOR DI(409) XOR DI(726) XOR DI(41) XOR DI(850) XOR DI(554) XOR DI(823) XOR DI(431) XOR DI(145) XOR DI(630) XOR DI(572) XOR DI(155) XOR DI(213) XOR DI(990) XOR DI(490) XOR DI(218) XOR DI(969) XOR DI(536) XOR DI(348) XOR DI(1006) XOR DI(429) XOR DI(779) XOR DI(451) XOR DI(165) XOR DI(825) XOR DI(514) XOR DI(209) XOR DI(739) XOR DI(275) XOR DI(214) XOR DI(231) XOR DI(477) XOR DI(626) XOR DI(879) XOR DI(650) XOR DI(242) XOR DI(600) XOR DI(497) XOR DI(22) XOR DI(903) XOR DI(815) XOR DI(539) XOR DI(890) XOR DI(991) XOR DI(7) XOR DI(280) XOR DI(327) XOR DI(297) XOR DI(118) XOR DI(126) XOR DI(32) XOR DI(39) XOR DI(912) XOR DI(955) XOR DI(207) XOR DI(828) XOR DI(899) XOR DI(370) XOR DI(212) XOR DI(530) XOR DI(342) XOR DI(119) XOR DI(423) XOR DI(819) XOR DI(269) XOR DI(208) XOR DI(724) XOR DI(713) XOR DI(873) XOR DI(236) XOR DI(491) XOR DI(16) XOR DI(62) XOR DI(410) XOR DI(985) XOR DI(722) XOR DI(399) XOR DI(210) XOR DI(629) XOR DI(18) XOR DI(386) XOR DI(112) XOR DI(176) XOR DI(120) XOR DI(260) XOR DI(669) XOR DI(618) XOR DI(143) XOR DI(206) XOR DI(336) XOR DI(153) XOR DI(813) XOR DI(465) XOR DI(707) XOR DI(867) XOR DI(527) XOR DI(393) XOR DI(315) XOR DI(546) XOR DI(663) XOR DI(950) XOR DI(943) XOR DI(147) XOR DI(701) XOR DI(861) XOR DI(198) XOR DI(540) XOR DI(937) XOR DI(695) XOR DI(689) XOR DI(528) XOR DI(683) XOR DI(522) XOR DI(123) XOR DI(516) XOR DI(510) XOR DI(1016) XOR DI(1022);
   DO(29) <= DI(584) XOR DI(773) XOR DI(277) XOR DI(86) XOR DI(306) XOR DI(569) XOR DI(556) XOR DI(50) XOR DI(870) XOR DI(66) XOR DI(838) XOR DI(966) XOR DI(752) XOR DI(179) XOR DI(549) XOR DI(953) XOR DI(577) XOR DI(446) XOR DI(602) XOR DI(699) XOR DI(479) XOR DI(263) XOR DI(101) XOR DI(672) XOR DI(434) XOR DI(784) XOR DI(289) XOR DI(228) XOR DI(54) XOR DI(621) XOR DI(519) XOR DI(372) XOR DI(915) XOR DI(425) XOR DI(612) XOR DI(245) XOR DI(877) XOR DI(401) XOR DI(884) XOR DI(769) XOR DI(709) XOR DI(640) XOR DI(893) XOR DI(285) XOR DI(863) XOR DI(194) XOR DI(760) XOR DI(77) XOR DI(271) XOR DI(859) XOR DI(80) XOR DI(36) XOR DI(563) XOR DI(346) XOR DI(787) XOR DI(756) XOR DI(987) XOR DI(849) XOR DI(114) XOR DI(486) XOR DI(693) XOR DI(971) XOR DI(791) XOR DI(252) XOR DI(1005) XOR DI(778) XOR DI(716) XOR DI(742) XOR DI(738) XOR DI(441) XOR DI(476) XOR DI(805) XOR DI(395) XOR DI(317) XOR DI(21) XOR DI(902) XOR DI(538) XOR DI(658) XOR DI(326) XOR DI(934) XOR DI(71) XOR DI(597) XOR DI(167) XOR DI(138) XOR DI(827) XOR DI(341) XOR DI(158) XOR DI(818) XOR DI(202) XOR DI(233) XOR DI(470) XOR DI(389) XOR DI(643) XOR DI(311) XOR DI(61) XOR DI(984) XOR DI(628) XOR DI(0) XOR DI(652) XOR DI(385) XOR DI(111) XOR DI(499) XOR DI(668) XOR DI(948) XOR DI(363) XOR DI(9) XOR DI(526) XOR DI(454) XOR DI(662) XOR DI(128) XOR DI(1009) XOR DI(1015) XOR DI(1021) XOR DI(767) XOR DI(774) XOR DI(278) XOR DI(444) XOR DI(378) XOR DI(307) XOR DI(570) XOR DI(51) XOR DI(871) XOR DI(91) XOR DI(836) XOR DI(331) XOR DI(763) XOR DI(732) XOR DI(610) XOR DI(190) XOR DI(964) XOR DI(180) XOR DI(550) XOR DI(151) XOR DI(578) XOR DI(646) XOR DI(185) XOR DI(480) XOR DI(382) XOR DI(798) XOR DI(224) XOR DI(264) XOR DI(102) XOR DI(765) XOR DI(785) XOR DI(457) XOR DI(229) XOR DI(55) XOR DI(916) XOR DI(255) XOR DI(246) XOR DI(439) XOR DI(656) XOR DI(248) XOR DI(606) XOR DI(324) XOR DI(28) XOR DI(74) XOR DI(959) XOR DI(770) XOR DI(107) XOR DI(222) XOR DI(710) XOR DI(641) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(333) XOR DI(810) XOR DI(864) XOR DI(195) XOR DI(473) XOR DI(761) XOR DI(78) XOR DI(272) XOR DI(81) XOR DI(564) XOR DI(788) XOR DI(293) XOR DI(988) XOR DI(554) XOR DI(972) XOR DI(834) XOR DI(376) XOR DI(792) XOR DI(253) XOR DI(536) XOR DI(921) XOR DI(1006) XOR DI(779) XOR DI(717) XOR DI(451) XOR DI(165) XOR DI(743) XOR DI(739) XOR DI(442) XOR DI(240) XOR DI(730) XOR DI(231) XOR DI(477) XOR DI(806) XOR DI(396) XOR DI(626) XOR DI(650) XOR DI(242) XOR DI(600) XOR DI(318) XOR DI(890) XOR DI(405) XOR DI(608) XOR DI(935) XOR DI(506) XOR DI(72) XOR DI(32) XOR DI(295) XOR DI(598) XOR DI(139) XOR DI(899) XOR DI(407) XOR DI(342) XOR DI(159) XOR DI(808) XOR DI(508) XOR DI(269) XOR DI(234) XOR DI(471) XOR DI(390) XOR DI(873) XOR DI(644) XOR DI(312) XOR DI(985) XOR DI(1) XOR DI(386) XOR DI(648) XOR DI(112) XOR DI(176) XOR DI(26) XOR DI(552) XOR DI(669) XOR DI(364) XOR DI(707) XOR DI(380) XOR DI(455) XOR DI(943) XOR DI(459) XOR DI(141) XOR DI(129) XOR DI(1010) XOR DI(1016) XOR DI(1022) XOR DI(575) XOR DI(999) XOR DI(41) XOR DI(353) XOR DI(768) XOR DI(775) XOR DI(905) XOR DI(85) XOR DI(445) XOR DI(301) XOR DI(88) XOR DI(44) XOR DI(308) XOR DI(52) XOR DI(939) XOR DI(49) XOR DI(924) XOR DI(354) XOR DI(688) XOR DI(92) XOR DI(795) XOR DI(925) XOR DI(837) XOR DI(68) XOR DI(611) XOR DI(191) XOR DI(300) XOR DI(467) XOR DI(857) XOR DI(968) XOR DI(965) XOR DI(830) XOR DI(955) XOR DI(637) XOR DI(579) XOR DI(703) XOR DI(122) XOR DI(448) XOR DI(162) XOR DI(65) XOR DI(701) XOR DI(979) XOR DI(841) XOR DI(997) XOR DI(530) XOR DI(383) XOR DI(173) XOR DI(926) XOR DI(799) XOR DI(225) XOR DI(635) XOR DI(940) XOR DI(355) XOR DI(132) XOR DI(674) XOR DI(759) XOR DI(896) XOR DI(436) XOR DI(299) XOR DI(562) XOR DI(786) XOR DI(755) XOR DI(724) XOR DI(172) XOR DI(542) XOR DI(56) XOR DI(623) XOR DI(358) XOR DI(521) XOR DI(704) XOR DI(123) XOR DI(750) XOR DI(887) XOR DI(533) XOR DI(614) XOR DI(737) XOR DI(440) XOR DI(212) XOR DI(484) XOR DI(813) XOR DI(726) XOR DI(886) XOR DI(657) XOR DI(249) XOR DI(325) XOR DI(419) XOR DI(465) XOR DI(493) XOR DI(70) XOR DI(852) XOR DI(321) XOR DI(75) XOR DI(137) XOR DI(147) XOR DI(771) XOR DI(108) XOR DI(735) XOR DI(412) XOR DI(469) XOR DI(642) XOR DI(895) XOR DI(927) XOR DI(666) XOR DI(287) XOR DI(590) XOR DI(304) XOR DI(283) XOR DI(661) XOR DI(125) XOR DI(356) XOR DI(145) XOR DI(532) XOR DI(929) XOR DI(474) XOR DI(1014) XOR DI(993) XOR DI(79) XOR DI(39) XOR DI(38) XOR DI(302) XOR DI(565) XOR DI(43) XOR DI(348) XOR DI(789) XOR DI(831) XOR DI(410) XOR DI(727) XOR DI(42) XOR DI(851) XOR DI(555) XOR DI(824) XOR DI(432) XOR DI(146) XOR DI(631) XOR DI(573) XOR DI(156) XOR DI(214) XOR DI(991) XOR DI(491) XOR DI(219) XOR DI(970) XOR DI(537) XOR DI(349) XOR DI(1007) XOR DI(430) XOR DI(780) XOR DI(452) XOR DI(166) XOR DI(826) XOR DI(515) XOR DI(210) XOR DI(740) XOR DI(276) XOR DI(215) XOR DI(232) XOR DI(478) XOR DI(627) XOR DI(880) XOR DI(651) XOR DI(243) XOR DI(601) XOR DI(498) XOR DI(23) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(891) XOR DI(992) XOR DI(8) XOR DI(281) XOR DI(328) XOR DI(298) XOR DI(119) XOR DI(127) XOR DI(33) XOR DI(40) XOR DI(913) XOR DI(956) XOR DI(208) XOR DI(829) XOR DI(900) XOR DI(371) XOR DI(213) XOR DI(531) XOR DI(343) XOR DI(120) XOR DI(424) XOR DI(820) XOR DI(270) XOR DI(209) XOR DI(725) XOR DI(714) XOR DI(874) XOR DI(237) XOR DI(492) XOR DI(17) XOR DI(63) XOR DI(411) XOR DI(986) XOR DI(723) XOR DI(400) XOR DI(211) XOR DI(630) XOR DI(19) XOR DI(387) XOR DI(113) XOR DI(177) XOR DI(121) XOR DI(261) XOR DI(670) XOR DI(619) XOR DI(144) XOR DI(207) XOR DI(337) XOR DI(154) XOR DI(814) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(528) XOR DI(394) XOR DI(316) XOR DI(547) XOR DI(664) XOR DI(951) XOR DI(944) XOR DI(148) XOR DI(702) XOR DI(862) XOR DI(199) XOR DI(541) XOR DI(938) XOR DI(696) XOR DI(690) XOR DI(529) XOR DI(684) XOR DI(523) XOR DI(124) XOR DI(517) XOR DI(511) XOR DI(1017) XOR DI(1023);
   DO(30) <= DI(352) XOR DI(585) XOR DI(767) XOR DI(774) XOR DI(278) XOR DI(866) XOR DI(444) XOR DI(87) XOR DI(378) XOR DI(335) XOR DI(307) XOR DI(570) XOR DI(977) XOR DI(557) XOR DI(51) XOR DI(923) XOR DI(687) XOR DI(871) XOR DI(91) XOR DI(794) XOR DI(836) XOR DI(67) XOR DI(331) XOR DI(415) XOR DI(974) XOR DI(763) XOR DI(732) XOR DI(610) XOR DI(47) XOR DI(104) XOR DI(190) XOR DI(839) XOR DI(560) XOR DI(967) XOR DI(964) XOR DI(753) XOR DI(180) XOR DI(550) XOR DI(954) XOR DI(151) XOR DI(578) XOR DI(447) XOR DI(161) XOR DI(603) XOR DI(646) XOR DI(700) XOR DI(3) XOR DI(185) XOR DI(908) XOR DI(366) XOR DI(480) XOR DI(911) XOR DI(996) XOR DI(382) XOR DI(496) XOR DI(588) XOR DI(798) XOR DI(259) XOR DI(224) XOR DI(634) XOR DI(6) XOR DI(712) XOR DI(264) XOR DI(102) XOR DI(187) XOR DI(131) XOR DI(673) XOR DI(1012) XOR DI(765) XOR DI(435) XOR DI(369) XOR DI(785) XOR DI(290) XOR DI(457) XOR DI(171) XOR DI(229) XOR DI(55) XOR DI(622) XOR DI(520) XOR DI(373) XOR DI(916) XOR DI(255) XOR DI(426) XOR DI(745) XOR DI(613) XOR DI(246) XOR DI(439) XOR DI(878) XOR DI(812) XOR DI(402) XOR DI(885) XOR DI(656) XOR DI(248) XOR DI(606) XOR DI(324) XOR DI(418) XOR DI(503) XOR DI(464) XOR DI(320) XOR DI(28) XOR DI(74) XOR DI(959) XOR DI(545) XOR DI(422) XOR DI(770) XOR DI(107) XOR DI(734) XOR DI(222) XOR DI(710) XOR DI(641) XOR DI(13) XOR DI(894) XOR DI(257) XOR DI(286) XOR DI(30) XOR DI(398) XOR DI(333) XOR DI(810) XOR DI(864) XOR DI(195) XOR DI(473) XOR DI(680) XOR DI(761) XOR DI(78) XOR DI(272) XOR DI(860) XOR DI(81) XOR DI(37) XOR DI(564) XOR DI(83) XOR DI(347) XOR DI(788) XOR DI(918) XOR DI(409) XOR DI(757) XOR DI(293) XOR DI(988) XOR DI(850) XOR DI(554) XOR DI(961) XOR DI(823) XOR DI(572) XOR DI(115) XOR DI(487) XOR DI(694) XOR DI(972) XOR DI(834) XOR DI(990) XOR DI(376) XOR DI(490) XOR DI(792) XOR DI(253) XOR DI(218) XOR DI(536) XOR DI(921) XOR DI(1006) XOR DI(429) XOR DI(779) XOR DI(748) XOR DI(717) XOR DI(451) XOR DI(165) XOR DI(514) XOR DI(743) XOR DI(739) XOR DI(442) XOR DI(240) XOR DI(730) XOR DI(231) XOR DI(477) XOR DI(806) XOR DI(719) XOR DI(396) XOR DI(626) XOR DI(650) XOR DI(242) XOR DI(600) XOR DI(318) XOR DI(314) XOR DI(22) XOR DI(903) XOR DI(539) XOR DI(890) XOR DI(405) XOR DI(659) XOR DI(280) XOR DI(392) XOR DI(327) XOR DI(297) XOR DI(118) XOR DI(182) XOR DI(608) XOR DI(935) XOR DI(506) XOR DI(72) XOR DI(32) XOR DI(266) XOR DI(295) XOR DI(598) XOR DI(168) XOR DI(139) XOR DI(828) XOR DI(899) XOR DI(407) XOR DI(342) XOR DI(159) XOR DI(808) XOR DI(819) XOR DI(508) XOR DI(203) XOR DI(269) XOR DI(234) XOR DI(471) XOR DI(390) XOR DI(873) XOR DI(644) XOR DI(236) XOR DI(312) XOR DI(16) XOR DI(62) XOR DI(985) XOR DI(722) XOR DI(629) XOR DI(1) XOR DI(653) XOR DI(274) XOR DI(386) XOR DI(648) XOR DI(112) XOR DI(176) XOR DI(500) XOR DI(461) XOR DI(26) XOR DI(552) XOR DI(669) XOR DI(949) XOR DI(143) XOR DI(364) XOR DI(206) XOR DI(153) XOR DI(197) XOR DI(707) XOR DI(10) XOR DI(527) XOR DI(380) XOR DI(455) XOR DI(663) XOR DI(943) XOR DI(459) XOR DI(617) XOR DI(937) XOR DI(141) XOR DI(855) XOR DI(482) XOR DI(135) XOR DI(129) XOR DI(683) XOR DI(677) XOR DI(510) XOR DI(1010) XOR DI(1016) XOR DI(1022) XOR DI(575) XOR DI(268) XOR DI(999) XOR DI(747) XOR DI(768) XOR DI(775) XOR DI(85) XOR DI(279) XOR DI(706) XOR DI(587) XOR DI(445) XOR DI(379) XOR DI(833) XOR DI(308) XOR DI(184) XOR DI(854) XOR DI(571) XOR DI(52) XOR DI(49) XOR DI(170) XOR DI(90) XOR DI(872) XOR DI(92) XOR DI(837) XOR DI(332) XOR DI(764) XOR DI(733) XOR DI(611) XOR DI(191) XOR DI(995) XOR DI(857) XOR DI(965) XOR DI(181) XOR DI(551) XOR DI(958) XOR DI(438) XOR DI(152) XOR DI(637) XOR DI(579) XOR DI(647) XOR DI(239) XOR DI(65) XOR DI(186) XOR DI(979) XOR DI(841) XOR DI(106) XOR DI(481) XOR DI(797) XOR DI(383) XOR DI(799) XOR DI(225) XOR DI(976) XOR DI(265) XOR DI(103) XOR DI(759) XOR DI(766) XOR DI(562) XOR DI(786) XOR DI(755) XOR DI(458) XOR DI(230) XOR DI(56) XOR DI(358) XOR DI(917) XOR DI(256) XOR DI(750) XOR DI(221) XOR DI(247) XOR DI(737) XOR DI(440) XOR DI(484) XOR DI(633) XOR DI(657) XOR DI(15) XOR DI(249) XOR DI(607) XOR DI(325) XOR DI(70) XOR DI(29) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(960) XOR DI(137) XOR DI(686) XOR DI(771) XOR DI(108) XOR DI(223) XOR DI(469) XOR DI(711) XOR DI(642) XOR DI(666) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(616) XOR DI(334) XOR DI(811) XOR DI(428) XOR DI(865) XOR DI(304) XOR DI(283) XOR DI(544) XOR DI(661) XOR DI(189) XOR DI(196) XOR DI(942) XOR DI(513) XOR DI(929) XOR DI(474) XOR DI(502) XOR DI(1014) XOR DI(762) XOR DI(79) XOR DI(273) XOR DI(82) XOR DI(330) XOR DI(323) XOR DI(565) XOR DI(46) XOR DI(164) XOR DI(682) XOR DI(789) XOR DI(605) XOR DI(294) XOR DI(989) XOR DI(555) XOR DI(175) XOR DI(432) XOR DI(351) XOR DI(156) XOR DI(973) XOR DI(835) XOR DI(679) XOR DI(414) XOR DI(377) XOR DI(920) XOR DI(793) XOR DI(254) XOR DI(970) XOR DI(537) XOR DI(922) XOR DI(1007) XOR DI(780) XOR DI(718) XOR DI(452) XOR DI(166) XOR DI(826) XOR DI(368) XOR DI(117) XOR DI(744) XOR DI(421) XOR DI(740) XOR DI(276) XOR DI(443) XOR DI(241) XOR DI(731) XOR DI(232) XOR DI(478) XOR DI(807) XOR DI(397) XOR DI(627) XOR DI(880) XOR DI(651) XOR DI(243) XOR DI(601) XOR DI(319) XOR DI(498) XOR DI(816) XOR DI(417) XOR DI(891) XOR DI(729) XOR DI(406) XOR DI(217) XOR DI(463) XOR DI(8) XOR DI(889) XOR DI(25) XOR DI(655) XOR DI(609) XOR DI(936) XOR DI(507) XOR DI(127) XOR DI(73) XOR DI(33) XOR DI(296) XOR DI(559) XOR DI(676) XOR DI(913) XOR DI(404) XOR DI(963) XOR DI(721) XOR DI(599) XOR DI(140) XOR DI(625) XOR DI(150) XOR DI(900) XOR DI(408) XOR DI(371) XOR DI(343) XOR DI(424) XOR DI(160) XOR DI(809) XOR DI(509) XOR DI(270) XOR DI(235) XOR DI(472) XOR DI(714) XOR DI(391) XOR DI(874) XOR DI(645) XOR DI(313) XOR DI(898) XOR DI(986) XOR DI(400) XOR DI(2) XOR DI(12) XOR DI(19) XOR DI(387) XOR DI(292) XOR DI(649) XOR DI(113) XOR DI(177) XOR DI(27) XOR DI(261) XOR DI(553) XOR DI(670) XOR DI(907) XOR DI(134) XOR DI(619) XOR DI(365) XOR DI(337) XOR DI(708) XOR DI(868) XOR DI(394) XOR DI(205) XOR DI(381) XOR DI(316) XOR DI(495) XOR DI(456) XOR DI(547) XOR DI(951) XOR DI(944) XOR DI(460) XOR DI(862) XOR DI(5) XOR DI(199) XOR DI(375) XOR DI(489) XOR DI(450) XOR DI(142) XOR DI(696) XOR DI(535) XOR DI(690) XOR DI(130) XOR DI(523) XOR DI(517) XOR DI(505) XOR DI(1011) XOR DI(1017) XOR DI(1023);
   DO(31) <= DI(575) XOR DI(268) XOR DI(999) XOR DI(41) XOR DI(747) XOR DI(353) XOR DI(586) XOR DI(768) XOR DI(775) XOR DI(905) XOR DI(85) XOR DI(45) XOR DI(279) XOR DI(867) XOR DI(706) XOR DI(587) XOR DI(445) XOR DI(301) XOR DI(88) XOR DI(379) XOR DI(336) XOR DI(833) XOR DI(994) XOR DI(329) XOR DI(44) XOR DI(796) XOR DI(308) XOR DI(184) XOR DI(854) XOR DI(571) XOR DI(978) XOR DI(558) XOR DI(52) XOR DI(89) XOR DI(939) XOR DI(49) XOR DI(170) XOR DI(90) XOR DI(924) XOR DI(354) XOR DI(688) XOR DI(872) XOR DI(92) XOR DI(574) XOR DI(795) XOR DI(925) XOR DI(837) XOR DI(68) XOR DI(332) XOR DI(416) XOR DI(975) XOR DI(764) XOR DI(733) XOR DI(611) XOR DI(48) XOR DI(105) XOR DI(191) XOR DI(300) XOR DI(840) XOR DI(467) XOR DI(995) XOR DI(857) XOR DI(561) XOR DI(968) XOR DI(965) XOR DI(754) XOR DI(181) XOR DI(830) XOR DI(551) XOR DI(958) XOR DI(955) XOR DI(438) XOR DI(152) XOR DI(637) XOR DI(357) XOR DI(579) XOR DI(703) XOR DI(122) XOR DI(448) XOR DI(162) XOR DI(220) XOR DI(736) XOR DI(604) XOR DI(647) XOR DI(239) XOR DI(494) XOR DI(65) XOR DI(701) XOR DI(632) XOR DI(4) XOR DI(186) XOR DI(909) XOR DI(979) XOR DI(841) XOR DI(106) XOR DI(685) XOR DI(367) XOR DI(481) XOR DI(912) XOR DI(997) XOR DI(420) XOR DI(797) XOR DI(530) XOR DI(383) XOR DI(173) XOR DI(926) XOR DI(497) XOR DI(589) XOR DI(799) XOR DI(260) XOR DI(225) XOR DI(635) XOR DI(303) XOR DI(7) XOR DI(976) XOR DI(713) XOR DI(265) XOR DI(103) XOR DI(543) XOR DI(940) XOR DI(355) XOR DI(188) XOR DI(928) XOR DI(132) XOR DI(674) XOR DI(1013) XOR DI(759) XOR DI(766) XOR DI(896) XOR DI(436) XOR DI(370) XOR DI(299) XOR DI(562) XOR DI(786) XOR DI(755) XOR DI(724) XOR DI(291) XOR DI(458) XOR DI(172) XOR DI(821) XOR DI(542) XOR DI(230) XOR DI(56) XOR DI(623) XOR DI(832) XOR DI(358) XOR DI(521) XOR DI(374) XOR DI(917) XOR DI(216) XOR DI(704) XOR DI(256) XOR DI(123) XOR DI(665) XOR DI(750) XOR DI(887) XOR DI(427) XOR DI(746) XOR DI(282) XOR DI(449) XOR DI(533) XOR DI(221) XOR DI(614) XOR DI(512) XOR DI(247) XOR DI(737) XOR DI(440) XOR DI(212) XOR DI(238) XOR DI(728) XOR DI(879) XOR DI(484) XOR DI(813) XOR DI(888) XOR DI(726) XOR DI(403) XOR DI(633) XOR DI(886) XOR DI(657) XOR DI(15) XOR DI(249) XOR DI(607) XOR DI(325) XOR DI(419) XOR DI(504) XOR DI(465) XOR DI(493) XOR DI(70) XOR DI(852) XOR DI(321) XOR DI(29) XOR DI(155) XOR DI(75) XOR DI(910) XOR DI(822) XOR DI(960) XOR DI(546) XOR DI(423) XOR DI(137) XOR DI(147) XOR DI(686) XOR DI(897) XOR DI(998) XOR DI(771) XOR DI(108) XOR DI(735) XOR DI(412) XOR DI(223) XOR DI(469) XOR DI(711) XOR DI(642) XOR DI(14) XOR DI(895) XOR DI(174) XOR DI(927) XOR DI(666) XOR DI(24) XOR DI(258) XOR DI(287) XOR DI(31) XOR DI(590) XOR DI(616) XOR DI(399) XOR DI(334) XOR DI(811) XOR DI(428) XOR DI(865) XOR DI(304) XOR DI(283) XOR DI(544) XOR DI(661) XOR DI(941) XOR DI(125) XOR DI(356) XOR DI(145) XOR DI(189) XOR DI(196) XOR DI(615) XOR DI(942) XOR DI(853) XOR DI(513) XOR DI(532) XOR DI(929) XOR DI(133) XOR DI(474) XOR DI(681) XOR DI(502) XOR DI(1014) XOR DI(993) XOR DI(762) XOR DI(79) XOR DI(39) XOR DI(273) XOR DI(861) XOR DI(82) XOR DI(330) XOR DI(323) XOR DI(38) XOR DI(302) XOR DI(565) XOR DI(46) XOR DI(43) XOR DI(164) XOR DI(84) XOR DI(348) XOR DI(682) XOR DI(789) XOR DI(919) XOR DI(831) XOR DI(410) XOR DI(969) XOR DI(758) XOR DI(727) XOR DI(605) XOR DI(42) XOR DI(294) XOR DI(989) XOR DI(851) XOR DI(555) XOR DI(962) XOR DI(175) XOR DI(824) XOR DI(432) XOR DI(146) XOR DI(631) XOR DI(351) XOR DI(573) XOR DI(116) XOR DI(156) XOR DI(214) XOR DI(488) XOR DI(695) XOR DI(973) XOR DI(835) XOR DI(679) XOR DI(906) XOR DI(991) XOR DI(414) XOR DI(377) XOR DI(920) XOR DI(491) XOR DI(793) XOR DI(254) XOR DI(219) XOR DI(970) XOR DI(537) XOR DI(349) XOR DI(922) XOR DI(126) XOR DI(1007) XOR DI(430) XOR DI(780) XOR DI(749) XOR DI(718) XOR DI(452) XOR DI(166) XOR DI(815) XOR DI(826) XOR DI(515) XOR DI(368) XOR DI(210) XOR DI(117) XOR DI(744) XOR DI(421) XOR DI(740) XOR DI(276) XOR DI(443) XOR DI(215) XOR DI(241) XOR DI(731) XOR DI(232) XOR DI(478) XOR DI(807) XOR DI(720) XOR DI(397) XOR DI(627) XOR DI(880) XOR DI(651) XOR DI(243) XOR DI(601) XOR DI(319) XOR DI(413) XOR DI(498) XOR DI(64) XOR DI(315) XOR DI(23) XOR DI(149) XOR DI(69) XOR DI(904) XOR DI(816) XOR DI(540) XOR DI(417) XOR DI(891) XOR DI(992) XOR DI(729) XOR DI(406) XOR DI(217) XOR DI(463) XOR DI(705) XOR DI(636) XOR DI(8) XOR DI(889) XOR DI(660) XOR DI(18) XOR DI(281) XOR DI(25) XOR DI(393) XOR DI(328) XOR DI(298) XOR DI(655) XOR DI(119) XOR DI(350) XOR DI(183) XOR DI(609) XOR DI(936) XOR DI(507) XOR DI(127) XOR DI(468) XOR DI(675) XOR DI(73) XOR DI(33) XOR DI(267) XOR DI(296) XOR DI(559) XOR DI(40) XOR DI(676) XOR DI(913) XOR DI(825) XOR DI(404) XOR DI(963) XOR DI(721) XOR DI(599) XOR DI(956) XOR DI(169) XOR DI(140) XOR DI(625) XOR DI(150) XOR DI(208) XOR DI(689) XOR DI(829) XOR DI(900) XOR DI(408) XOR DI(371) XOR DI(213) XOR DI(531) XOR DI(343) XOR DI(120) XOR DI(424) XOR DI(160) XOR DI(809) XOR DI(820) XOR DI(509) XOR DI(204) XOR DI(270) XOR DI(437) XOR DI(209) XOR DI(235) XOR DI(725) XOR DI(472) XOR DI(714) XOR DI(391) XOR DI(874) XOR DI(645) XOR DI(237) XOR DI(313) XOR DI(492) XOR DI(17) XOR DI(63) XOR DI(898) XOR DI(534) XOR DI(411) XOR DI(986) XOR DI(723) XOR DI(400) XOR DI(211) XOR DI(630) XOR DI(2) XOR DI(654) XOR DI(12) XOR DI(275) XOR DI(19) XOR DI(387) XOR DI(322) XOR DI(292) XOR DI(649) XOR DI(113) XOR DI(177) XOR DI(501) XOR DI(121) XOR DI(462) XOR DI(27) XOR DI(261) XOR DI(553) XOR DI(670) XOR DI(907) XOR DI(957) XOR DI(950) XOR DI(163) XOR DI(134) XOR DI(619) XOR DI(144) XOR DI(365) XOR DI(207) XOR DI(337) XOR DI(154) XOR DI(814) XOR DI(198) XOR DI(431) XOR DI(466) XOR DI(708) XOR DI(868) XOR DI(11) XOR DI(528) XOR DI(394) XOR DI(205) XOR DI(624) XOR DI(381) XOR DI(316) XOR DI(495) XOR DI(456) XOR DI(547) XOR DI(664) XOR DI(951) XOR DI(944) XOR DI(148) XOR DI(460) XOR DI(702) XOR DI(862) XOR DI(5) XOR DI(522) XOR DI(199) XOR DI(618) XOR DI(375) XOR DI(489) XOR DI(450) XOR DI(541) XOR DI(938) XOR DI(142) XOR DI(696) XOR DI(856) XOR DI(516) XOR DI(483) XOR DI(535) XOR DI(136) XOR DI(690) XOR DI(529) XOR DI(130) XOR DI(684) XOR DI(523) XOR DI(124) XOR DI(678) XOR DI(517) XOR DI(511) XOR DI(505) XOR DI(1011) XOR DI(1017) XOR DI(1023);
end architecture;