library ieee;
use ieee.std_logic_1164.all;

entity top is
 port(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146: in std_logic;
po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341: std_logic;

begin

w0 <= not pi013 and not pi014;
w1 <= not pi006 and not pi007;
w2 <= w0 and w1;
w3 <= not pi017 and not pi021;
w4 <= not pi008 and w3;
w5 <= not pi012 and w4;
w6 <= w2 and w5;
w7 <= not pi018 and not pi019;
w8 <= not pi004 and not pi016;
w9 <= w7 and w8;
w10 <= not pi005 and not pi022;
w11 <= not pi009 and not pi011;
w12 <= w10 and w11;
w13 <= w9 and w12;
w14 <= w6 and w13;
w15 <= pi054 and not w14;
w16 <= not pi000 and not w15;
w17 <= w10 and not w11;
w18 <= not pi056 and w17;
w19 <= not pi056 and not w10;
w20 <= not pi008 and not pi021;
w21 <= not pi007 and pi013;
w22 <= w20 and w21;
w23 <= not pi007 and w20;
w24 <= pi007 and not w20;
w25 <= not w23 and not w24;
w26 <= pi008 and pi021;
w27 <= not pi013 and not w26;
w28 <= w25 and w27;
w29 <= not w22 and not w28;
w30 <= not pi014 and not w29;
w31 <= not pi013 and pi014;
w32 <= w23 and w31;
w33 <= not w30 and not w32;
w34 <= not pi010 and not w33;
w35 <= pi010 and w0;
w36 <= w23 and w35;
w37 <= not w34 and not w36;
w38 <= w10 and not w37;
w39 <= w9 and w38;
w40 <= not pi017 and w39;
w41 <= not pi006 and not pi012;
w42 <= w40 and w41;
w43 <= not w19 and not w42;
w44 <= w11 and not w43;
w45 <= not w18 and not w44;
w46 <= pi054 and not w45;
w47 <= not w16 and not w46;
w48 <= not pi129 and not w47;
w49 <= not pi003 and w48;
w50 <= not pi011 and not pi012;
w51 <= w20 and w50;
w52 <= w9 and w51;
w53 <= not pi010 and not pi022;
w54 <= not pi007 and not pi013;
w55 <= not pi005 and not pi006;
w56 <= w54 and w55;
w57 <= not pi014 and w56;
w58 <= w53 and w57;
w59 <= w52 and w58;
w60 <= not pi017 and pi054;
w61 <= not w59 and w60;
w62 <= not pi001 and not w61;
w63 <= not pi014 and pi054;
w64 <= not pi008 and not pi011;
w65 <= w3 and w64;
w66 <= not pi005 and w41;
w67 <= pi005 and not w41;
w68 <= not w66 and not w67;
w69 <= pi006 and pi012;
w70 <= not pi007 and not w69;
w71 <= w68 and w70;
w72 <= pi007 and w66;
w73 <= not w71 and not w72;
w74 <= not pi013 and not w73;
w75 <= w21 and w66;
w76 <= not w74 and not w75;
w77 <= not pi009 and not w76;
w78 <= w54 and w66;
w79 <= pi009 and w78;
w80 <= not w77 and not w79;
w81 <= w9 and not w80;
w82 <= w65 and w81;
w83 <= w63 and w82;
w84 <= w53 and w83;
w85 <= not w62 and not w84;
w86 <= not pi129 and not w85;
w87 <= not pi003 and w86;
w88 <= pi122 and pi127;
w89 <= not pi045 and not pi048;
w90 <= not pi043 and not pi047;
w91 <= w89 and w90;
w92 <= not pi015 and not pi020;
w93 <= not pi024 and not pi049;
w94 <= w92 and w93;
w95 <= w91 and w94;
w96 <= not pi041 and not pi046;
w97 <= not pi038 and not pi050;
w98 <= w96 and w97;
w99 <= not pi042 and not pi044;
w100 <= not pi040 and w99;
w101 <= not pi002 and w100;
w102 <= w98 and w101;
w103 <= w95 and w102;
w104 <= pi082 and not w103;
w105 <= not w88 and not w104;
w106 <= not pi065 and w105;
w107 <= not pi024 and not pi045;
w108 <= not pi047 and not pi048;
w109 <= w107 and w108;
w110 <= not pi049 and w92;
w111 <= w109 and w110;
w112 <= not pi038 and not pi040;
w113 <= w99 and w112;
w114 <= not pi046 and not pi050;
w115 <= not pi041 and w114;
w116 <= w113 and w115;
w117 <= not pi043 and w116;
w118 <= w111 and w117;
w119 <= pi082 and not w118;
w120 <= not pi082 and w88;
w121 <= not w119 and not w120;
w122 <= pi002 and not w121;
w123 <= not w106 and not w122;
w124 <= not pi129 and not w123;
w125 <= not pi009 and not pi014;
w126 <= w53 and w125;
w127 <= w56 and w126;
w128 <= not pi008 and not pi017;
w129 <= w50 and w128;
w130 <= not pi021 and w9;
w131 <= w129 and w130;
w132 <= w127 and w131;
w133 <= not pi061 and not pi118;
w134 <= not w132 and w133;
w135 <= pi000 and not pi123;
w136 <= not pi113 and w135;
w137 <= not w134 and not w136;
w138 <= not pi129 and not w137;
w139 <= pi010 and not pi022;
w140 <= w125 and w139;
w141 <= w78 and w140;
w142 <= pi054 and w9;
w143 <= w65 and w142;
w144 <= w141 and w143;
w145 <= pi004 and not pi054;
w146 <= not w144 and not w145;
w147 <= not pi129 and not w146;
w148 <= not pi003 and w147;
w149 <= pi005 and not pi054;
w150 <= not pi007 and w41;
w151 <= not pi025 and not pi029;
w152 <= pi028 and w151;
w153 <= w150 and w152;
w154 <= not pi013 and w126;
w155 <= w153 and w154;
w156 <= not pi059 and w65;
w157 <= not pi016 and pi054;
w158 <= not pi004 and not pi019;
w159 <= not pi018 and w158;
w160 <= not pi005 and w159;
w161 <= w157 and w160;
w162 <= w156 and w161;
w163 <= w155 and w162;
w164 <= not w149 and not w163;
w165 <= not pi129 and not w164;
w166 <= not pi003 and w165;
w167 <= pi006 and not pi054;
w168 <= not pi005 and not pi007;
w169 <= pi025 and not pi029;
w170 <= not pi028 and w169;
w171 <= not pi012 and w170;
w172 <= w168 and w171;
w173 <= w154 and w172;
w174 <= not pi006 and w159;
w175 <= w157 and w174;
w176 <= w156 and w175;
w177 <= w173 and w176;
w178 <= not w167 and not w177;
w179 <= not pi129 and not w178;
w180 <= not pi003 and w179;
w181 <= pi007 and not pi054;
w182 <= not pi018 and not pi021;
w183 <= pi008 and not pi017;
w184 <= w182 and w183;
w185 <= not pi007 and w158;
w186 <= w157 and w185;
w187 <= w184 and w186;
w188 <= not pi006 and w50;
w189 <= not pi005 and w188;
w190 <= w154 and w189;
w191 <= w187 and w190;
w192 <= not w181 and not w191;
w193 <= not pi129 and not w192;
w194 <= not pi003 and w193;
w195 <= pi008 and not pi054;
w196 <= w78 and w126;
w197 <= not pi017 and not pi018;
w198 <= not pi011 and pi021;
w199 <= w197 and w198;
w200 <= not pi008 and w158;
w201 <= w157 and w200;
w202 <= w199 and w201;
w203 <= w196 and w202;
w204 <= not w195 and not w203;
w205 <= not pi129 and not w204;
w206 <= not pi003 and w205;
w207 <= pi009 and not pi054;
w208 <= w0 and w53;
w209 <= pi011 and w168;
w210 <= w41 and w209;
w211 <= w208 and w210;
w212 <= w128 and w182;
w213 <= not pi009 and w158;
w214 <= w157 and w213;
w215 <= w212 and w214;
w216 <= w211 and w215;
w217 <= not w207 and not w216;
w218 <= not pi129 and not w217;
w219 <= not pi003 and w218;
w220 <= pi010 and not pi054;
w221 <= not pi010 and w158;
w222 <= w157 and w221;
w223 <= w212 and w222;
w224 <= w168 and w188;
w225 <= not pi009 and not pi022;
w226 <= w31 and w225;
w227 <= w224 and w226;
w228 <= w223 and w227;
w229 <= not w220 and not w228;
w230 <= not pi129 and not w229;
w231 <= not pi003 and w230;
w232 <= pi011 and not pi054;
w233 <= not pi011 and w158;
w234 <= w157 and w233;
w235 <= w212 and w234;
w236 <= not pi010 and pi022;
w237 <= w125 and w236;
w238 <= w78 and w237;
w239 <= w235 and w238;
w240 <= not w232 and not w239;
w241 <= not pi129 and not w240;
w242 <= not pi003 and w241;
w243 <= pi012 and not pi054;
w244 <= not pi012 and w158;
w245 <= w157 and w244;
w246 <= pi018 and w4;
w247 <= w245 and w246;
w248 <= not pi011 and w127;
w249 <= w247 and w248;
w250 <= not w243 and not w249;
w251 <= not pi129 and not w250;
w252 <= not pi003 and w251;
w253 <= pi013 and not pi054;
w254 <= not pi013 and w159;
w255 <= w157 and w254;
w256 <= w156 and w255;
w257 <= not pi025 and pi029;
w258 <= not pi028 and w257;
w259 <= w66 and w258;
w260 <= not pi007 and w126;
w261 <= w259 and w260;
w262 <= w256 and w261;
w263 <= not w253 and not w262;
w264 <= not pi129 and not w263;
w265 <= not pi003 and w264;
w266 <= pi014 and not pi054;
w267 <= not pi016 and w63;
w268 <= w158 and w267;
w269 <= w212 and w268;
w270 <= not pi009 and pi013;
w271 <= w53 and w270;
w272 <= w224 and w271;
w273 <= w269 and w272;
w274 <= not w266 and not w273;
w275 <= not pi129 and not w274;
w276 <= not pi003 and w275;
w277 <= not pi041 and not pi043;
w278 <= w108 and w277;
w279 <= not pi045 and w93;
w280 <= w278 and w279;
w281 <= not pi046 and w97;
w282 <= w100 and w281;
w283 <= not pi015 and w282;
w284 <= w280 and w283;
w285 <= pi082 and not w284;
w286 <= not w88 and not w285;
w287 <= not pi070 and w286;
w288 <= not pi048 and w90;
w289 <= w279 and w288;
w290 <= w116 and w289;
w291 <= pi015 and not w290;
w292 <= not pi045 and w108;
w293 <= not pi002 and not pi020;
w294 <= not pi015 and not w293;
w295 <= w117 and w294;
w296 <= w93 and w295;
w297 <= w292 and w296;
w298 <= not w291 and not w297;
w299 <= pi082 and not w298;
w300 <= pi015 and w120;
w301 <= not w299 and not w300;
w302 <= not w287 and w301;
w303 <= not pi129 and not w302;
w304 <= pi016 and not pi054;
w305 <= pi006 and not pi012;
w306 <= not pi005 and w305;
w307 <= w54 and w306;
w308 <= w126 and w307;
w309 <= w143 and w308;
w310 <= not w304 and not w309;
w311 <= not pi129 and not w310;
w312 <= not pi003 and w311;
w313 <= pi017 and not pi054;
w314 <= not pi007 and w55;
w315 <= not pi025 and not pi028;
w316 <= not pi012 and w315;
w317 <= w314 and w316;
w318 <= w154 and w317;
w319 <= not pi016 and w60;
w320 <= w159 and w319;
w321 <= not pi011 and w20;
w322 <= not pi029 and pi059;
w323 <= w321 and w322;
w324 <= w320 and w323;
w325 <= w318 and w324;
w326 <= not w313 and not w325;
w327 <= not pi129 and not w326;
w328 <= not pi003 and w327;
w329 <= pi018 and not pi054;
w330 <= pi016 and pi054;
w331 <= w159 and w330;
w332 <= w65 and w331;
w333 <= w196 and w332;
w334 <= not w329 and not w333;
w335 <= not pi129 and not w334;
w336 <= not pi003 and w335;
w337 <= pi019 and not pi054;
w338 <= pi017 and w321;
w339 <= not pi004 and not pi018;
w340 <= not pi019 and w339;
w341 <= w157 and w340;
w342 <= w338 and w341;
w343 <= w196 and w342;
w344 <= not w337 and not w343;
w345 <= not pi129 and not w344;
w346 <= not pi003 and w345;
w347 <= w90 and w96;
w348 <= not pi024 and w89;
w349 <= w347 and w348;
w350 <= not pi040 and not pi042;
w351 <= w97 and w350;
w352 <= not pi044 and w110;
w353 <= w351 and w352;
w354 <= w349 and w353;
w355 <= pi082 and not w354;
w356 <= not w88 and not w355;
w357 <= not pi071 and w356;
w358 <= not pi050 and w112;
w359 <= not pi015 and not pi049;
w360 <= w99 and w359;
w361 <= w358 and w360;
w362 <= w349 and w361;
w363 <= pi020 and not w362;
w364 <= pi002 and w354;
w365 <= not w363 and not w364;
w366 <= pi082 and not w365;
w367 <= pi020 and w120;
w368 <= not w366 and not w367;
w369 <= not w357 and w368;
w370 <= not pi129 and not w369;
w371 <= pi021 and not pi054;
w372 <= w64 and w197;
w373 <= not pi021 and pi054;
w374 <= pi019 and w373;
w375 <= w8 and w374;
w376 <= w372 and w375;
w377 <= w196 and w376;
w378 <= not w371 and not w377;
w379 <= not pi129 and not w378;
w380 <= not pi003 and w379;
w381 <= pi022 and not pi054;
w382 <= not pi022 and w158;
w383 <= w157 and w382;
w384 <= w212 and w383;
w385 <= not pi009 and not pi010;
w386 <= w0 and w385;
w387 <= pi005 and not pi007;
w388 <= w188 and w387;
w389 <= w386 and w388;
w390 <= w384 and w389;
w391 <= not w381 and not w390;
w392 <= not pi129 and not w391;
w393 <= not pi003 and w392;
w394 <= not pi023 and pi055;
w395 <= not pi129 and not w394;
w396 <= pi061 and w395;
w397 <= not pi047 and w277;
w398 <= w89 and w397;
w399 <= w282 and w398;
w400 <= pi082 and not w399;
w401 <= w293 and w359;
w402 <= pi082 and not w401;
w403 <= w88 and not w402;
w404 <= not w400 and not w403;
w405 <= not pi024 and not w404;
w406 <= not pi002 and not pi045;
w407 <= w108 and w406;
w408 <= w110 and w407;
w409 <= w117 and w408;
w410 <= pi082 and not w409;
w411 <= not w88 and not w410;
w412 <= pi063 and w411;
w413 <= not pi043 and w96;
w414 <= w292 and w413;
w415 <= pi024 and pi082;
w416 <= w99 and w415;
w417 <= w358 and w416;
w418 <= w414 and w417;
w419 <= not pi129 and not w418;
w420 <= not w412 and w419;
w421 <= not w405 and w420;
w422 <= pi085 and pi116;
w423 <= not pi085 and not pi110;
w424 <= not pi096 and w423;
w425 <= not w422 and not w424;
w426 <= pi100 and not w425;
w427 <= pi025 and not pi116;
w428 <= pi085 and w427;
w429 <= not w426 and not w428;
w430 <= not pi026 and not w429;
w431 <= not pi051 and not pi052;
w432 <= not pi039 and w431;
w433 <= not pi095 and not pi100;
w434 <= not pi097 and w433;
w435 <= not pi110 and not w434;
w436 <= pi025 and not w435;
w437 <= pi026 and pi116;
w438 <= not w436 and not w437;
w439 <= not w432 and not w438;
w440 <= pi026 and w427;
w441 <= not w439 and not w440;
w442 <= not pi085 and not w441;
w443 <= not w430 and not w442;
w444 <= not pi027 and not w443;
w445 <= not pi039 and not pi052;
w446 <= not pi051 and w445;
w447 <= pi116 and w446;
w448 <= not w427 and not w447;
w449 <= pi027 and not w448;
w450 <= w432 and w436;
w451 <= not w449 and not w450;
w452 <= not pi026 and not pi085;
w453 <= not w451 and w452;
w454 <= not w444 and not w453;
w455 <= not pi053 and not w454;
w456 <= pi025 and not pi026;
w457 <= not pi116 and w456;
w458 <= pi053 and not pi085;
w459 <= not pi027 and w458;
w460 <= w457 and w459;
w461 <= not w455 and not w460;
w462 <= not pi058 and not w461;
w463 <= not pi027 and not pi085;
w464 <= not pi053 and pi058;
w465 <= w463 and w464;
w466 <= w457 and w465;
w467 <= not w462 and not w466;
w468 <= not pi129 and not w467;
w469 <= not pi003 and w468;
w470 <= pi085 and not pi116;
w471 <= not pi110 and not w470;
w472 <= not w437 and w471;
w473 <= not pi096 and w472;
w474 <= not pi026 and w422;
w475 <= not w473 and not w474;
w476 <= pi100 and not w475;
w477 <= not pi085 and not w447;
w478 <= pi026 and w477;
w479 <= not w476 and not w478;
w480 <= not pi129 and not w479;
w481 <= not pi003 and w480;
w482 <= not pi027 and not pi053;
w483 <= not pi058 and w482;
w484 <= w481 and w483;
w485 <= pi095 and not pi096;
w486 <= pi027 and pi116;
w487 <= w471 and not w486;
w488 <= w485 and w487;
w489 <= not pi027 and w422;
w490 <= not w488 and not w489;
w491 <= not pi100 and not w490;
w492 <= pi027 and w477;
w493 <= not w491 and not w492;
w494 <= not pi129 and not w493;
w495 <= not pi003 and w494;
w496 <= not pi053 and not pi058;
w497 <= not pi026 and w496;
w498 <= w495 and w497;
w499 <= not pi026 and not w432;
w500 <= not pi027 and w446;
w501 <= not w499 and not w500;
w502 <= not w435 and not w501;
w503 <= pi026 and not pi027;
w504 <= not pi026 and pi027;
w505 <= not w503 and not w504;
w506 <= not pi116 and not w505;
w507 <= not w502 and not w506;
w508 <= pi028 and not w507;
w509 <= not pi026 and not pi100;
w510 <= not pi110 and w509;
w511 <= w485 and w510;
w512 <= w437 and w446;
w513 <= not w511 and not w512;
w514 <= not pi027 and not w513;
w515 <= w486 and w499;
w516 <= not w514 and not w515;
w517 <= not w508 and w516;
w518 <= not pi085 and not w517;
w519 <= pi028 and not pi116;
w520 <= not pi100 and pi116;
w521 <= not w519 and not w520;
w522 <= pi085 and not w521;
w523 <= not pi026 and not pi027;
w524 <= w522 and w523;
w525 <= not w518 and not w524;
w526 <= not pi053 and not w525;
w527 <= not pi027 and pi028;
w528 <= not pi116 and w527;
w529 <= not pi026 and w458;
w530 <= w528 and w529;
w531 <= not w526 and not w530;
w532 <= not pi058 and not w531;
w533 <= w452 and w464;
w534 <= w528 and w533;
w535 <= not w532 and not w534;
w536 <= not pi129 and not w535;
w537 <= not pi003 and w536;
w538 <= pi029 and pi110;
w539 <= pi097 and not pi110;
w540 <= not pi096 and w539;
w541 <= pi029 and not pi097;
w542 <= not w540 and not w541;
w543 <= w433 and not w542;
w544 <= not w538 and not w543;
w545 <= not pi058 and not w544;
w546 <= pi097 and pi116;
w547 <= pi029 and not pi116;
w548 <= not w546 and not w547;
w549 <= pi058 and not w548;
w550 <= not w545 and not w549;
w551 <= not pi053 and not w550;
w552 <= pi053 and not pi058;
w553 <= w547 and w552;
w554 <= not w551 and not w553;
w555 <= not pi027 and not w554;
w556 <= pi027 and w547;
w557 <= w496 and w556;
w558 <= not w555 and not w557;
w559 <= not pi085 and not w558;
w560 <= pi085 and w483;
w561 <= w547 and w560;
w562 <= not w559 and not w561;
w563 <= not pi026 and not w562;
w564 <= w463 and w496;
w565 <= pi026 and w564;
w566 <= w547 and w565;
w567 <= not w563 and not w566;
w568 <= not pi129 and not w567;
w569 <= not pi003 and w568;
w570 <= pi030 and not pi109;
w571 <= pi060 and pi109;
w572 <= not w570 and not w571;
w573 <= not pi106 and not w572;
w574 <= pi088 and pi106;
w575 <= not w573 and not w574;
w576 <= not pi129 and not w575;
w577 <= pi089 and pi106;
w578 <= pi030 and pi109;
w579 <= pi031 and not pi109;
w580 <= not w578 and not w579;
w581 <= not pi106 and not w580;
w582 <= not w577 and not w581;
w583 <= not pi129 and not w582;
w584 <= pi099 and pi106;
w585 <= pi031 and pi109;
w586 <= pi032 and not pi109;
w587 <= not w585 and not w586;
w588 <= not pi106 and not w587;
w589 <= not w584 and not w588;
w590 <= not pi129 and not w589;
w591 <= pi090 and pi106;
w592 <= pi032 and pi109;
w593 <= pi033 and not pi109;
w594 <= not w592 and not w593;
w595 <= not pi106 and not w594;
w596 <= not w591 and not w595;
w597 <= not pi129 and not w596;
w598 <= pi091 and pi106;
w599 <= pi033 and pi109;
w600 <= pi034 and not pi109;
w601 <= not w599 and not w600;
w602 <= not pi106 and not w601;
w603 <= not w598 and not w602;
w604 <= not pi129 and not w603;
w605 <= pi092 and pi106;
w606 <= pi034 and pi109;
w607 <= pi035 and not pi109;
w608 <= not w606 and not w607;
w609 <= not pi106 and not w608;
w610 <= not w605 and not w609;
w611 <= not pi129 and not w610;
w612 <= pi098 and pi106;
w613 <= pi035 and pi109;
w614 <= pi036 and not pi109;
w615 <= not w613 and not w614;
w616 <= not pi106 and not w615;
w617 <= not w612 and not w616;
w618 <= not pi129 and not w617;
w619 <= pi093 and pi106;
w620 <= pi036 and pi109;
w621 <= pi037 and not pi109;
w622 <= not w620 and not w621;
w623 <= not pi106 and not w622;
w624 <= not w619 and not w623;
w625 <= not pi129 and not w624;
w626 <= pi082 and not w100;
w627 <= w115 and w288;
w628 <= w94 and w406;
w629 <= w627 and w628;
w630 <= pi082 and not w629;
w631 <= w88 and not w630;
w632 <= not w626 and not w631;
w633 <= not pi038 and not w632;
w634 <= not pi002 and not pi048;
w635 <= w107 and w634;
w636 <= w110 and w635;
w637 <= not pi050 and w100;
w638 <= w347 and w637;
w639 <= w636 and w638;
w640 <= pi082 and not w639;
w641 <= not w88 and not w640;
w642 <= pi074 and w641;
w643 <= not pi044 and pi082;
w644 <= pi038 and w350;
w645 <= w643 and w644;
w646 <= not pi129 and not w645;
w647 <= not w642 and w646;
w648 <= not w633 and w647;
w649 <= not pi051 and pi109;
w650 <= w445 and w649;
w651 <= not pi106 and not w650;
w652 <= pi109 and w431;
w653 <= pi039 and not w652;
w654 <= w651 and not w653;
w655 <= not pi129 and not w654;
w656 <= pi082 and not w99;
w657 <= w288 and w628;
w658 <= w98 and w657;
w659 <= pi082 and not w658;
w660 <= w88 and not w659;
w661 <= not w656 and not w660;
w662 <= not pi040 and not w661;
w663 <= w97 and w99;
w664 <= w347 and w663;
w665 <= w636 and w664;
w666 <= pi082 and not w665;
w667 <= not w88 and not w666;
w668 <= pi073 and w667;
w669 <= pi040 and pi082;
w670 <= w99 and w669;
w671 <= not pi129 and not w670;
w672 <= not w668 and w671;
w673 <= not w662 and w672;
w674 <= pi082 and not w282;
w675 <= pi082 and not w657;
w676 <= w88 and not w675;
w677 <= not w674 and not w676;
w678 <= not pi041 and not w677;
w679 <= w90 and w114;
w680 <= w113 and w679;
w681 <= w636 and w680;
w682 <= pi082 and not w681;
w683 <= not w88 and not w682;
w684 <= pi076 and w683;
w685 <= w112 and w114;
w686 <= pi041 and pi082;
w687 <= w99 and w686;
w688 <= w685 and w687;
w689 <= not pi129 and not w688;
w690 <= not w684 and w689;
w691 <= not w678 and w690;
w692 <= pi044 and pi082;
w693 <= w397 and w685;
w694 <= w636 and w693;
w695 <= pi082 and not w694;
w696 <= w88 and not w695;
w697 <= not w692 and not w696;
w698 <= not pi042 and not w697;
w699 <= not pi044 and w358;
w700 <= w347 and w699;
w701 <= w636 and w700;
w702 <= pi082 and not w701;
w703 <= not w88 and not w702;
w704 <= pi072 and w703;
w705 <= pi042 and w643;
w706 <= not pi129 and not w705;
w707 <= not w704 and w706;
w708 <= not w698 and w707;
w709 <= pi082 and not w116;
w710 <= w94 and w407;
w711 <= pi082 and not w710;
w712 <= w88 and not w711;
w713 <= not w709 and not w712;
w714 <= not pi043 and not w713;
w715 <= not pi047 and w116;
w716 <= w636 and w715;
w717 <= pi082 and not w716;
w718 <= not w88 and not w717;
w719 <= pi077 and w718;
w720 <= pi043 and w350;
w721 <= w643 and w720;
w722 <= w98 and w721;
w723 <= not pi129 and not w722;
w724 <= not w719 and w723;
w725 <= not w714 and w724;
w726 <= w347 and w351;
w727 <= w636 and w726;
w728 <= pi082 and not w727;
w729 <= pi067 and not w88;
w730 <= not pi044 and w88;
w731 <= not w729 and not w730;
w732 <= not w728 and not w731;
w733 <= not pi129 and not w692;
w734 <= not w732 and w733;
w735 <= w108 and w413;
w736 <= w97 and w100;
w737 <= w735 and w736;
w738 <= pi082 and not w737;
w739 <= not pi024 and w401;
w740 <= pi082 and not w739;
w741 <= w88 and not w740;
w742 <= not w738 and not w741;
w743 <= not pi045 and not w742;
w744 <= not pi002 and w108;
w745 <= w94 and w744;
w746 <= w117 and w745;
w747 <= pi082 and not w746;
w748 <= not w88 and not w747;
w749 <= pi068 and w748;
w750 <= not pi038 and w350;
w751 <= pi045 and w750;
w752 <= w643 and w751;
w753 <= w627 and w752;
w754 <= not pi129 and not w753;
w755 <= not w749 and w754;
w756 <= not w743 and w755;
w757 <= pi082 and not w736;
w758 <= w397 and w636;
w759 <= pi082 and not w758;
w760 <= w88 and not w759;
w761 <= not w757 and not w760;
w762 <= not pi046 and not w761;
w763 <= not pi050 and w113;
w764 <= w758 and w763;
w765 <= pi082 and not w764;
w766 <= not w88 and not w765;
w767 <= pi075 and w766;
w768 <= pi046 and pi082;
w769 <= w763 and w768;
w770 <= not pi129 and not w769;
w771 <= not w767 and w770;
w772 <= not w762 and w771;
w773 <= pi082 and not w117;
w774 <= pi082 and not w636;
w775 <= w88 and not w774;
w776 <= not w773 and not w775;
w777 <= not pi047 and not w776;
w778 <= w117 and w636;
w779 <= pi082 and not w778;
w780 <= not w88 and not w779;
w781 <= pi064 and w780;
w782 <= w277 and w281;
w783 <= pi047 and w350;
w784 <= w643 and w783;
w785 <= w782 and w784;
w786 <= not pi129 and not w785;
w787 <= not w781 and w786;
w788 <= not w777 and w787;
w789 <= w347 and w736;
w790 <= pi082 and not w789;
w791 <= pi082 and not w628;
w792 <= w88 and not w791;
w793 <= not w790 and not w792;
w794 <= not pi048 and not w793;
w795 <= not pi002 and not pi047;
w796 <= w107 and w110;
w797 <= w795 and w796;
w798 <= w117 and w797;
w799 <= pi082 and not w798;
w800 <= not w88 and not w799;
w801 <= pi062 and w800;
w802 <= w90 and w115;
w803 <= pi048 and w750;
w804 <= w643 and w803;
w805 <= w802 and w804;
w806 <= not pi129 and not w805;
w807 <= not w801 and w806;
w808 <= not w794 and w807;
w809 <= w93 and w763;
w810 <= w414 and w809;
w811 <= pi082 and not w810;
w812 <= not w88 and not w811;
w813 <= not pi069 and w812;
w814 <= not pi024 and not pi042;
w815 <= w699 and w814;
w816 <= w414 and w815;
w817 <= pi049 and not w816;
w818 <= not pi002 and w92;
w819 <= w809 and not w818;
w820 <= w347 and w819;
w821 <= w89 and w820;
w822 <= not w817 and not w821;
w823 <= pi082 and not w822;
w824 <= pi049 and w120;
w825 <= not w823 and not w824;
w826 <= not w813 and w825;
w827 <= not pi129 and not w826;
w828 <= pi082 and not w113;
w829 <= w413 and w744;
w830 <= w796 and w829;
w831 <= pi082 and not w830;
w832 <= w88 and not w831;
w833 <= not w828 and not w832;
w834 <= not pi050 and not w833;
w835 <= w113 and w347;
w836 <= w636 and w835;
w837 <= pi082 and not w836;
w838 <= not w88 and not w837;
w839 <= pi066 and w838;
w840 <= pi050 and w750;
w841 <= w643 and w840;
w842 <= not pi129 and not w841;
w843 <= not w839 and w842;
w844 <= not w834 and w843;
w845 <= pi051 and not pi109;
w846 <= not w649 and not w845;
w847 <= not pi106 and w846;
w848 <= not pi129 and not w847;
w849 <= pi052 and not w649;
w850 <= not pi106 and not w652;
w851 <= not w849 and w850;
w852 <= not pi129 and not w851;
w853 <= pi058 and pi116;
w854 <= not pi058 and not pi110;
w855 <= not pi096 and w854;
w856 <= w433 and w855;
w857 <= not w853 and not w856;
w858 <= not pi053 and not w857;
w859 <= pi097 and w858;
w860 <= not pi116 and w552;
w861 <= not w859 and not w860;
w862 <= not pi129 and not w861;
w863 <= not pi003 and w862;
w864 <= w463 and w863;
w865 <= not pi026 and w864;
w866 <= w117 and w710;
w867 <= pi082 and not w866;
w868 <= not w88 and not w867;
w869 <= not pi129 and not w868;
w870 <= not pi123 and not pi129;
w871 <= pi114 and not pi122;
w872 <= w870 and w871;
w873 <= not pi026 and pi058;
w874 <= pi026 and not pi058;
w875 <= pi116 and w874;
w876 <= not w873 and not w875;
w877 <= pi094 and not w876;
w878 <= pi058 and not pi116;
w879 <= pi037 and not pi116;
w880 <= not w873 and not w879;
w881 <= not w878 and not w880;
w882 <= not w877 and not w881;
w883 <= not pi053 and not w882;
w884 <= not pi026 and pi037;
w885 <= not pi058 and w884;
w886 <= not w883 and not w885;
w887 <= not pi085 and not w886;
w888 <= w496 and w884;
w889 <= not w887 and not w888;
w890 <= not pi027 and not w889;
w891 <= not pi085 and w496;
w892 <= w884 and w891;
w893 <= not w890 and not w892;
w894 <= not pi129 and not w893;
w895 <= not pi003 and w894;
w896 <= not pi026 and not pi053;
w897 <= pi026 and pi053;
w898 <= not pi085 and not w897;
w899 <= not w896 and not w898;
w900 <= not pi058 and not w899;
w901 <= not pi085 and w896;
w902 <= not pi116 and w901;
w903 <= not w900 and not w902;
w904 <= pi057 and not w903;
w905 <= pi060 and w853;
w906 <= w901 and w905;
w907 <= not w904 and not w906;
w908 <= not pi027 and not w907;
w909 <= pi057 and not pi058;
w910 <= w901 and w909;
w911 <= not w908 and not w910;
w912 <= not pi129 and not w911;
w913 <= not pi003 and w912;
w914 <= w523 and w878;
w915 <= pi116 and not w505;
w916 <= not pi058 and w915;
w917 <= w446 and w916;
w918 <= not w914 and not w917;
w919 <= not pi129 and not w918;
w920 <= not pi003 and w919;
w921 <= not pi053 and w920;
w922 <= not pi085 and w921;
w923 <= not w464 and not w552;
w924 <= not pi116 and not w923;
w925 <= not w435 and w496;
w926 <= not w924 and not w925;
w927 <= pi059 and not w926;
w928 <= w435 and w496;
w929 <= pi096 and w928;
w930 <= not w927 and not w929;
w931 <= not pi085 and not w930;
w932 <= pi059 and not pi116;
w933 <= pi085 and w496;
w934 <= w932 and w933;
w935 <= not w931 and not w934;
w936 <= not pi027 and not w935;
w937 <= pi027 and w891;
w938 <= w932 and w937;
w939 <= not w936 and not w938;
w940 <= not pi026 and not w939;
w941 <= w565 and w932;
w942 <= not w940 and not w941;
w943 <= not pi129 and not w942;
w944 <= not pi003 and w943;
w945 <= not pi117 and not pi122;
w946 <= pi060 and not w945;
w947 <= pi123 and w945;
w948 <= not w946 and not w947;
w949 <= not pi114 and pi123;
w950 <= not pi122 and w949;
w951 <= not pi129 and w950;
w952 <= not pi137 and not pi138;
w953 <= pi136 and w952;
w954 <= pi132 and pi133;
w955 <= pi131 and w954;
w956 <= w953 and w955;
w957 <= pi062 and not w956;
w958 <= pi136 and not pi137;
w959 <= not pi140 and w958;
w960 <= not pi138 and w955;
w961 <= w959 and w960;
w962 <= not w957 and not w961;
w963 <= not pi129 and not w962;
w964 <= pi063 and not w956;
w965 <= not pi142 and w958;
w966 <= w960 and w965;
w967 <= not w964 and not w966;
w968 <= not pi129 and not w967;
w969 <= pi064 and not w956;
w970 <= not pi139 and w958;
w971 <= w960 and w970;
w972 <= not w969 and not w971;
w973 <= not pi129 and not w972;
w974 <= pi065 and not w956;
w975 <= not pi146 and w958;
w976 <= w960 and w975;
w977 <= not w974 and not w976;
w978 <= not pi129 and not w977;
w979 <= not pi136 and not pi137;
w980 <= w960 and w979;
w981 <= pi066 and not w980;
w982 <= not pi143 and w980;
w983 <= not w981 and not w982;
w984 <= not pi129 and not w983;
w985 <= pi067 and not w980;
w986 <= not pi139 and w980;
w987 <= not w985 and not w986;
w988 <= not pi129 and not w987;
w989 <= pi068 and not w956;
w990 <= not pi141 and w958;
w991 <= w960 and w990;
w992 <= not w989 and not w991;
w993 <= not pi129 and not w992;
w994 <= pi069 and not w956;
w995 <= not pi143 and w958;
w996 <= w960 and w995;
w997 <= not w994 and not w996;
w998 <= not pi129 and not w997;
w999 <= pi070 and not w956;
w1000 <= not pi144 and w958;
w1001 <= w960 and w1000;
w1002 <= not w999 and not w1001;
w1003 <= not pi129 and not w1002;
w1004 <= pi071 and not w956;
w1005 <= not pi145 and w958;
w1006 <= w960 and w1005;
w1007 <= not w1004 and not w1006;
w1008 <= not pi129 and not w1007;
w1009 <= pi072 and not w980;
w1010 <= not pi140 and w980;
w1011 <= not w1009 and not w1010;
w1012 <= not pi129 and not w1011;
w1013 <= pi073 and not w980;
w1014 <= not pi141 and w980;
w1015 <= not w1013 and not w1014;
w1016 <= not pi129 and not w1015;
w1017 <= pi074 and not w980;
w1018 <= not pi142 and w980;
w1019 <= not w1017 and not w1018;
w1020 <= not pi129 and not w1019;
w1021 <= pi075 and not w980;
w1022 <= not pi144 and w980;
w1023 <= not w1021 and not w1022;
w1024 <= not pi129 and not w1023;
w1025 <= pi076 and not w980;
w1026 <= not pi145 and w980;
w1027 <= not w1025 and not w1026;
w1028 <= not pi129 and not w1027;
w1029 <= pi077 and not w980;
w1030 <= not pi146 and w980;
w1031 <= not w1029 and not w1030;
w1032 <= not pi129 and not w1031;
w1033 <= not pi136 and pi137;
w1034 <= w960 and w1033;
w1035 <= pi078 and not w1034;
w1036 <= pi142 and w1034;
w1037 <= not w1035 and not w1036;
w1038 <= not pi129 and not w1037;
w1039 <= pi079 and not w1034;
w1040 <= pi143 and w1034;
w1041 <= not w1039 and not w1040;
w1042 <= not pi129 and not w1041;
w1043 <= pi080 and not w1034;
w1044 <= pi144 and w1034;
w1045 <= not w1043 and not w1044;
w1046 <= not pi129 and not w1045;
w1047 <= pi081 and not w1034;
w1048 <= pi145 and w1034;
w1049 <= not w1047 and not w1048;
w1050 <= not pi129 and not w1049;
w1051 <= pi082 and not w1034;
w1052 <= pi146 and w1034;
w1053 <= not w1051 and not w1052;
w1054 <= not pi129 and not w1053;
w1055 <= pi089 and pi138;
w1056 <= not pi062 and not pi138;
w1057 <= not w1055 and not w1056;
w1058 <= pi136 and not w1057;
w1059 <= pi119 and pi138;
w1060 <= not pi072 and not pi138;
w1061 <= not w1059 and not w1060;
w1062 <= not pi136 and not w1061;
w1063 <= not w1058 and not w1062;
w1064 <= not pi137 and not w1063;
w1065 <= not pi115 and pi138;
w1066 <= pi087 and not pi138;
w1067 <= not w1065 and not w1066;
w1068 <= not pi136 and not w1067;
w1069 <= pi136 and not pi138;
w1070 <= pi031 and w1069;
w1071 <= not w1068 and not w1070;
w1072 <= pi137 and not w1071;
w1073 <= not w1064 and not w1072;
w1074 <= pi084 and not w1034;
w1075 <= pi141 and w1034;
w1076 <= not w1074 and not w1075;
w1077 <= not pi129 and not w1076;
w1078 <= not pi085 and not w434;
w1079 <= not pi110 and w1078;
w1080 <= pi096 and w1079;
w1081 <= not w470 and not w1080;
w1082 <= not pi129 and not w1081;
w1083 <= not pi003 and w1082;
w1084 <= w483 and w1083;
w1085 <= not pi026 and w1084;
w1086 <= pi086 and not w1034;
w1087 <= pi139 and w1034;
w1088 <= not w1086 and not w1087;
w1089 <= not pi129 and not w1088;
w1090 <= pi087 and not w1034;
w1091 <= pi140 and w1034;
w1092 <= not w1090 and not w1091;
w1093 <= not pi129 and not w1092;
w1094 <= pi136 and pi137;
w1095 <= w960 and w1094;
w1096 <= pi088 and not w1095;
w1097 <= pi139 and w1095;
w1098 <= not w1096 and not w1097;
w1099 <= not pi129 and not w1098;
w1100 <= pi089 and not w1095;
w1101 <= pi140 and w1095;
w1102 <= not w1100 and not w1101;
w1103 <= not pi129 and not w1102;
w1104 <= pi090 and not w1095;
w1105 <= pi142 and w1095;
w1106 <= not w1104 and not w1105;
w1107 <= not pi129 and not w1106;
w1108 <= pi091 and not w1095;
w1109 <= pi143 and w1095;
w1110 <= not w1108 and not w1109;
w1111 <= not pi129 and not w1110;
w1112 <= pi092 and not w1095;
w1113 <= pi144 and w1095;
w1114 <= not w1112 and not w1113;
w1115 <= not pi129 and not w1114;
w1116 <= pi093 and not w1095;
w1117 <= pi146 and w1095;
w1118 <= not w1116 and not w1117;
w1119 <= not pi129 and not w1118;
w1120 <= pi082 and not pi137;
w1121 <= not pi136 and w1120;
w1122 <= pi138 and w955;
w1123 <= w1121 and w1122;
w1124 <= pi094 and not w1123;
w1125 <= pi142 and w1123;
w1126 <= not w1124 and not w1125;
w1127 <= not pi129 and not w1126;
w1128 <= not pi003 and not w955;
w1129 <= not pi110 and w1128;
w1130 <= pi138 and w1121;
w1131 <= w955 and not w1130;
w1132 <= not w1129 and not w1131;
w1133 <= pi095 and not w1132;
w1134 <= pi143 and w1123;
w1135 <= not w1133 and not w1134;
w1136 <= not pi129 and not w1135;
w1137 <= pi096 and not w1132;
w1138 <= pi146 and w1123;
w1139 <= not w1137 and not w1138;
w1140 <= not pi129 and not w1139;
w1141 <= pi097 and not w1132;
w1142 <= pi145 and w1123;
w1143 <= not w1141 and not w1142;
w1144 <= not pi129 and not w1143;
w1145 <= pi098 and not w1095;
w1146 <= pi145 and w1095;
w1147 <= not w1145 and not w1146;
w1148 <= not pi129 and not w1147;
w1149 <= pi099 and not w1095;
w1150 <= pi141 and w1095;
w1151 <= not w1149 and not w1150;
w1152 <= not pi129 and not w1151;
w1153 <= pi100 and not w1132;
w1154 <= pi144 and w1123;
w1155 <= not w1153 and not w1154;
w1156 <= not pi129 and not w1155;
w1157 <= pi124 and pi138;
w1158 <= not pi077 and not pi138;
w1159 <= not w1157 and not w1158;
w1160 <= not pi136 and not w1159;
w1161 <= not pi065 and not pi138;
w1162 <= pi093 and pi138;
w1163 <= not w1161 and not w1162;
w1164 <= pi136 and not w1163;
w1165 <= not w1160 and not w1164;
w1166 <= not pi137 and not w1165;
w1167 <= pi037 and w1069;
w1168 <= pi096 and pi138;
w1169 <= pi082 and not pi138;
w1170 <= not w1168 and not w1169;
w1171 <= not pi136 and not w1170;
w1172 <= not w1167 and not w1171;
w1173 <= pi137 and not w1172;
w1174 <= not w1166 and not w1173;
w1175 <= pi091 and w958;
w1176 <= pi095 and w1033;
w1177 <= not w1175 and not w1176;
w1178 <= pi138 and not w1177;
w1179 <= pi079 and not pi136;
w1180 <= pi034 and pi136;
w1181 <= not w1179 and not w1180;
w1182 <= pi137 and not w1181;
w1183 <= not pi069 and pi136;
w1184 <= not pi066 and not pi136;
w1185 <= not w1183 and not w1184;
w1186 <= not pi137 and not w1185;
w1187 <= not w1182 and not w1186;
w1188 <= not pi138 and not w1187;
w1189 <= not w1178 and not w1188;
w1190 <= pi090 and w958;
w1191 <= pi094 and w1033;
w1192 <= not w1190 and not w1191;
w1193 <= pi138 and not w1192;
w1194 <= pi078 and not pi136;
w1195 <= pi033 and pi136;
w1196 <= not w1194 and not w1195;
w1197 <= pi137 and not w1196;
w1198 <= not pi063 and pi136;
w1199 <= not pi074 and not pi136;
w1200 <= not w1198 and not w1199;
w1201 <= not pi137 and not w1200;
w1202 <= not w1197 and not w1201;
w1203 <= not pi138 and not w1202;
w1204 <= not w1193 and not w1203;
w1205 <= pi099 and w958;
w1206 <= not pi112 and w1033;
w1207 <= not w1205 and not w1206;
w1208 <= pi138 and not w1207;
w1209 <= not pi068 and pi136;
w1210 <= not pi073 and not pi136;
w1211 <= not w1209 and not w1210;
w1212 <= not pi137 and not w1211;
w1213 <= pi084 and not pi136;
w1214 <= pi032 and pi136;
w1215 <= not w1213 and not w1214;
w1216 <= pi137 and not w1215;
w1217 <= not w1212 and not w1216;
w1218 <= not pi138 and not w1217;
w1219 <= not w1208 and not w1218;
w1220 <= pi092 and pi138;
w1221 <= not pi070 and not pi138;
w1222 <= not w1220 and not w1221;
w1223 <= pi136 and not w1222;
w1224 <= pi125 and pi138;
w1225 <= not pi075 and not pi138;
w1226 <= not w1224 and not w1225;
w1227 <= not pi136 and not w1226;
w1228 <= not w1223 and not w1227;
w1229 <= not pi137 and not w1228;
w1230 <= pi080 and not pi138;
w1231 <= pi100 and pi138;
w1232 <= not w1230 and not w1231;
w1233 <= not pi136 and not w1232;
w1234 <= pi035 and w1069;
w1235 <= not w1233 and not w1234;
w1236 <= pi137 and not w1235;
w1237 <= not w1229 and not w1236;
w1238 <= w497 and w1079;
w1239 <= not pi027 and w1238;
w1240 <= not w422 and not w1239;
w1241 <= not pi129 and not w1240;
w1242 <= not pi003 and w1241;
w1243 <= pi098 and pi138;
w1244 <= not pi071 and not pi138;
w1245 <= not w1243 and not w1244;
w1246 <= pi136 and not w1245;
w1247 <= not pi076 and not pi138;
w1248 <= pi023 and pi138;
w1249 <= not w1247 and not w1248;
w1250 <= not pi136 and not w1249;
w1251 <= not w1246 and not w1250;
w1252 <= not pi137 and not w1251;
w1253 <= pi036 and w1069;
w1254 <= pi081 and not pi138;
w1255 <= pi097 and pi138;
w1256 <= not w1254 and not w1255;
w1257 <= not pi136 and not w1256;
w1258 <= not w1253 and not w1257;
w1259 <= pi137 and not w1258;
w1260 <= not w1252 and not w1259;
w1261 <= pi088 and pi138;
w1262 <= not pi064 and not pi138;
w1263 <= not w1261 and not w1262;
w1264 <= pi136 and not w1263;
w1265 <= pi120 and pi138;
w1266 <= not pi067 and not pi138;
w1267 <= not w1265 and not w1266;
w1268 <= not pi136 and not w1267;
w1269 <= not w1264 and not w1268;
w1270 <= not pi137 and not w1269;
w1271 <= pi086 and not pi138;
w1272 <= pi111 and pi138;
w1273 <= not w1271 and not w1272;
w1274 <= not pi136 and not w1273;
w1275 <= pi030 and w1069;
w1276 <= not w1274 and not w1275;
w1277 <= pi137 and not w1276;
w1278 <= not w1270 and not w1277;
w1279 <= not w446 and w504;
w1280 <= not w503 and not w1279;
w1281 <= not pi129 and not w1280;
w1282 <= not pi003 and w1281;
w1283 <= pi116 and w1282;
w1284 <= not pi097 and w464;
w1285 <= not w552 and not w1284;
w1286 <= not pi129 and not w1285;
w1287 <= not pi003 and w1286;
w1288 <= pi116 and w1287;
w1289 <= pi111 and not w1130;
w1290 <= not pi136 and pi139;
w1291 <= not pi137 and pi138;
w1292 <= pi082 and w1291;
w1293 <= w1290 and w1292;
w1294 <= not w1289 and not w1293;
w1295 <= w955 and not w1294;
w1296 <= not pi129 and w1295;
w1297 <= not pi136 and pi141;
w1298 <= w1292 and w1297;
w1299 <= not pi112 and not w1130;
w1300 <= not w1298 and not w1299;
w1301 <= w955 and not w1300;
w1302 <= not pi129 and w1301;
w1303 <= not pi054 and not pi113;
w1304 <= not pi011 and not pi022;
w1305 <= pi054 and not w1304;
w1306 <= not w1303 and not w1305;
w1307 <= not pi129 and not w1306;
w1308 <= not pi003 and w1307;
w1309 <= not pi136 and pi140;
w1310 <= w1292 and w1309;
w1311 <= not pi115 and not w1130;
w1312 <= not w1310 and not w1311;
w1313 <= w955 and not w1312;
w1314 <= not pi129 and w1313;
w1315 <= not pi004 and not pi012;
w1316 <= not pi007 and not pi009;
w1317 <= w1315 and w1316;
w1318 <= not pi129 and not w1317;
w1319 <= not pi003 and w1318;
w1320 <= pi054 and w1319;
w1321 <= pi122 and not pi129;
w1322 <= not pi054 and pi118;
w1323 <= pi054 and not pi059;
w1324 <= w258 and w1323;
w1325 <= not w1322 and not w1324;
w1326 <= not pi129 and not w1325;
w1327 <= not pi129 and not w433;
w1328 <= not pi110 and not pi120;
w1329 <= not pi003 and w1328;
w1330 <= not pi129 and not w1329;
w1331 <= not pi111 and w1330;
w1332 <= pi081 and pi120;
w1333 <= not pi129 and w1332;
w1334 <= not pi129 and not pi134;
w1335 <= not pi129 and not pi135;
w1336 <= pi057 and not pi129;
w1337 <= not pi096 and pi125;
w1338 <= not pi003 and not w1337;
w1339 <= not pi129 and not w1338;
w1340 <= not pi126 and pi132;
w1341 <= pi133 and w1340;
one <= '1';
po000 <= pi108;-- level 0
po001 <= pi083;-- level 0
po002 <= pi104;-- level 0
po003 <= pi103;-- level 0
po004 <= pi102;-- level 0
po005 <= pi105;-- level 0
po006 <= pi107;-- level 0
po007 <= pi101;-- level 0
po008 <= pi126;-- level 0
po009 <= pi121;-- level 0
po010 <= pi001;-- level 0
po011 <= pi000;-- level 0
po012 <= one;-- level 0
po013 <= pi130;-- level 0
po014 <= pi128;-- level 0
po015 <= not w49;-- level 20
po016 <= not w87;-- level 16
po017 <= w124;-- level 10
po018 <= w138;-- level 8
po019 <= w148;-- level 8
po020 <= w166;-- level 9
po021 <= w180;-- level 9
po022 <= w194;-- level 8
po023 <= w206;-- level 8
po024 <= w219;-- level 8
po025 <= w231;-- level 8
po026 <= w242;-- level 8
po027 <= w252;-- level 8
po028 <= w265;-- level 9
po029 <= w276;-- level 8
po030 <= w303;-- level 12
po031 <= w312;-- level 8
po032 <= w328;-- level 8
po033 <= w336;-- level 8
po034 <= w346;-- level 8
po035 <= w370;-- level 11
po036 <= w380;-- level 8
po037 <= w393;-- level 8
po038 <= w396;-- level 3
po039 <= w421;-- level 10
po040 <= w469;-- level 17
po041 <= w484;-- level 10
po042 <= w498;-- level 10
po043 <= w537;-- level 16
po044 <= w569;-- level 17
po045 <= w576;-- level 5
po046 <= w583;-- level 5
po047 <= w590;-- level 5
po048 <= w597;-- level 5
po049 <= w604;-- level 5
po050 <= w611;-- level 5
po051 <= w618;-- level 5
po052 <= w625;-- level 5
po053 <= w648;-- level 10
po054 <= w655;-- level 5
po055 <= w673;-- level 10
po056 <= w691;-- level 9
po057 <= w708;-- level 10
po058 <= w725;-- level 10
po059 <= w734;-- level 7
po060 <= w756;-- level 10
po061 <= w772;-- level 10
po062 <= w788;-- level 10
po063 <= w808;-- level 10
po064 <= w827;-- level 12
po065 <= w844;-- level 9
po066 <= w848;-- level 4
po067 <= w852;-- level 5
po068 <= w865;-- level 11
po069 <= not w869;-- level 8
po070 <= w872;-- level 2
po071 <= w895;-- level 13
po072 <= w913;-- level 11
po073 <= w922;-- level 10
po074 <= w944;-- level 15
po075 <= not w948;-- level 3
po076 <= w951;-- level 3
po077 <= not w963;-- level 6
po078 <= not w968;-- level 6
po079 <= not w973;-- level 6
po080 <= not w978;-- level 6
po081 <= not w984;-- level 7
po082 <= not w988;-- level 7
po083 <= not w993;-- level 6
po084 <= not w998;-- level 6
po085 <= not w1003;-- level 6
po086 <= not w1008;-- level 6
po087 <= not w1012;-- level 7
po088 <= not w1016;-- level 7
po089 <= not w1020;-- level 7
po090 <= not w1024;-- level 7
po091 <= not w1028;-- level 7
po092 <= not w1032;-- level 7
po093 <= w1038;-- level 7
po094 <= w1042;-- level 7
po095 <= w1046;-- level 7
po096 <= w1050;-- level 7
po097 <= w1054;-- level 7
po098 <= not w1073;-- level 6
po099 <= w1077;-- level 7
po100 <= w1085;-- level 10
po101 <= w1089;-- level 7
po102 <= w1093;-- level 7
po103 <= w1099;-- level 7
po104 <= w1103;-- level 7
po105 <= w1107;-- level 7
po106 <= w1111;-- level 7
po107 <= w1115;-- level 7
po108 <= w1119;-- level 7
po109 <= w1127;-- level 7
po110 <= w1136;-- level 8
po111 <= w1140;-- level 8
po112 <= w1144;-- level 8
po113 <= w1148;-- level 7
po114 <= w1152;-- level 7
po115 <= w1156;-- level 8
po116 <= not w1174;-- level 6
po117 <= not w1189;-- level 6
po118 <= not w1204;-- level 6
po119 <= not w1219;-- level 6
po120 <= not w1237;-- level 6
po121 <= w1242;-- level 9
po122 <= not w1260;-- level 6
po123 <= not w1278;-- level 6
po124 <= w1283;-- level 7
po125 <= w1288;-- level 6
po126 <= w1296;-- level 7
po127 <= w1302;-- level 7
po128 <= w1308;-- level 5
po129 <= not w870;-- level 1
po130 <= w1314;-- level 7
po131 <= w1320;-- level 5
po132 <= not w1321;-- level 1
po133 <= w1326;-- level 5
po134 <= w1327;-- level 2
po135 <= w1331;-- level 4
po136 <= w1333;-- level 2
po137 <= not w1334;-- level 1
po138 <= not w1335;-- level 1
po139 <= w1336;-- level 1
po140 <= w1339;-- level 3
po141 <= w1341;-- level 2
end Behavioral;