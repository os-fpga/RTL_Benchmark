// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_dsp (
    core_clk,
    core_reset_n,
    dsp_instr_valid,
    dsp_operand_ctrl,
    dsp_function_ctrl,
    dsp_result_ctrl,
    dsp_overflow_ctrl,
    dsp_data_src1,
    dsp_data_src2,
    dsp_data_src3,
    dsp_data_src4,
    dsp_stage2_pipe_en,
    dsp_stage3_pipe_en,
    dsp_stage1_result,
    dsp_stage1_ovf_set,
    dsp_stage2_result,
    dsp_stage2_ovf_set,
    dsp_stage3_result,
    dsp_stage3_ovf_set
);
localparam DSP_OCTRL_WIDTH = 44;
localparam DSP_FCTRL_WIDTH = 151;
localparam DSP_RCTRL_WIDTH = 70;
localparam SHIFT_AMT_MSB = 4;
input core_clk;
input core_reset_n;
input dsp_instr_valid;
input [DSP_OCTRL_WIDTH - 1:0] dsp_operand_ctrl;
input [DSP_FCTRL_WIDTH - 1:0] dsp_function_ctrl;
input [DSP_RCTRL_WIDTH - 1:0] dsp_result_ctrl;
input dsp_overflow_ctrl;
input [31:0] dsp_data_src1;
input [31:0] dsp_data_src2;
input [31:0] dsp_data_src3;
input [31:0] dsp_data_src4;
input dsp_stage2_pipe_en;
input dsp_stage3_pipe_en;
output [63:0] dsp_stage1_result;
output dsp_stage1_ovf_set;
output [63:0] dsp_stage2_result;
output dsp_stage2_ovf_set;
output [63:0] dsp_stage3_result;
output dsp_stage3_ovf_set;


integer i;
wire operand_simd_op16;
wire operand_simd_cross_op16;
wire operand_simd_clip_op16;
wire operand_simd_op8;
wire operand_simd_clip_op8;
wire operand_simd_cross_op8;
wire operand_psimd_op32;
wire operand_psimd_opxlen;
wire operand_psimd_op16b_op16b;
wire operand_psimd_op16b_op16t;
wire operand_psimd_op16t_op16b;
wire operand_psimd_op16t_op16t;
wire operand_psimd_clip_op32;
wire operand_psimd_op64;
wire operand_psimd_op32_op16b;
wire operand_psimd_op32_op16t;
wire operand_psimd_op16;
wire operand_psimd_cross_op16;
wire operand_psimd_reverse_op16;
wire operand_psimd_smal_op16;
wire operand_psimd_op8;
wire operand_psimd_cross_op8;
wire operand_64p_opxlen;
wire operand_64p_op16b_op16b;
wire operand_64p_op16b_op16t;
wire operand_64p_op16t_op16t;
wire operand_64p_op16;
wire operand_64p_cross_op16;
wire operand_64p_reverse_op16;
wire operand_nsimd_s_op32_sexlen;
wire operand_nsimd_u_op32_sexlen;
wire operand_nsimd_op16b_op16b;
wire operand_nsimd_op16b_op16t;
wire operand_nsimd_op16t_op16t;
wire operand_nsimd_op32;
wire operand_nsimd_opxlen;
wire operand_simd_op32;
wire operand_simd_cross_op32;
wire operand_psimd_op32b_op32b;
wire operand_psimd_op32b_op32t;
wire operand_psimd_op32t_op32t;
wire operand_psimd_cross_op32;
wire operand_psimd_reverse_op32;
wire operand_psimd_op32t_op32b;
wire function_simd_s_add16;
wire function_simd_u_add16;
wire function_simd_s_sub16;
wire function_simd_u_sub16;
wire function_simd_s_as16;
wire function_simd_u_as16;
wire function_simd_s_sa16;
wire function_simd_u_sa16;
wire function_simd_s_sra16;
wire function_simd_u_srl16;
wire function_simd_s_sll16;
wire function_simd_s_slra16;
wire function_simd_s_cmpeq16;
wire function_simd_s_cmplt16;
wire function_simd_u_cmplt16;
wire function_simd_s_cmple16;
wire function_simd_u_cmple16;
wire function_simd_s_min16;
wire function_simd_u_min16;
wire function_simd_s_max16;
wire function_simd_u_max16;
wire function_simd_s_abs16;
wire function_simd_s_clip16;
wire function_simd_s_mul16;
wire function_simd_s_swap16;
wire function_simd_s_clz16;
wire function_simd_s_clo16;
wire function_simd_s_clrs16;
wire function_simd_s_add8;
wire function_simd_u_add8;
wire function_simd_s_sub8;
wire function_simd_u_sub8;
wire function_simd_s_sra8;
wire function_simd_u_srl8;
wire function_simd_s_sll8;
wire function_simd_s_slra8;
wire function_simd_s_cmpeq8;
wire function_simd_s_cmplt8;
wire function_simd_u_cmplt8;
wire function_simd_s_cmple8;
wire function_simd_u_cmple8;
wire function_simd_s_min8;
wire function_simd_u_min8;
wire function_simd_s_max8;
wire function_simd_u_max8;
wire function_simd_s_abs8;
wire function_simd_s_clip8;
wire function_simd_s_mul8;
wire function_simd_s_swap8;
wire function_simd_s_clz8;
wire function_simd_s_clo8;
wire function_simd_s_clrs8;
wire function_simd_s_unpk8_10;
wire function_simd_s_unpk8_20;
wire function_simd_s_unpk8_30;
wire function_simd_s_unpk8_31;
wire function_simd_s_unpk8_32;
wire function_psimd_s_add32;
wire function_psimd_u_add32;
wire function_psimd_s_sub32;
wire function_psimd_u_sub32;
wire function_psimd_s_sraxlen;
wire function_psimd_s_sll32;
wire function_psimd_s_pk16;
wire function_psimd_s_clip32;
wire function_psimd_u_bitrevxlen;
wire function_psimd_s_wext32;
wire function_psimd_s_bpickxlen;
wire function_psimd_s_insbxlen;
wire function_psimd_s_min32;
wire function_psimd_s_max32;
wire function_psimd_s_abs32;
wire function_psimd_s_clz32;
wire function_psimd_s_clo32;
wire function_psimd_s_clrs32;
wire function_psimd_s_mul32x32_acc32_func0;
wire function_psimd_s_mul32x32_acc32_func1;
wire function_psimd_s_mul32x32_acc32_func2;
wire function_psimd_s_mul32x32_acc32_func3;
wire function_psimd_s_mul32x32_acc32_func4;
wire function_psimd_s_mul32x32_acc32_func5;
wire function_psimd_s_mul32x16_acc32_func0;
wire function_psimd_s_mul32x16_acc32_func1;
wire function_psimd_s_mul32x16_acc32_func2;
wire function_psimd_s_mul32x16_acc32_func3;
wire function_psimd_s_mul16x16_acc32_func0;
wire function_psimd_s_mul16x16_acc32_func1;
wire function_psimd_s_mul16x16_acc32_func2;
wire function_psimd_s_mul16x16_acc32_func3;
wire function_psimd_s_mul16x16_acc32_func4;
wire function_psimd_s_mul16x16_acc32_func5;
wire function_psimd_s_mul16x16_acc32_func6;
wire function_psimd_s_mul16x16_acc64_func0;
wire function_psimd_s_mul8x8_acc32_func0;
wire function_psimd_s_mul8x8_acc32_func1;
wire function_psimd_s_mul8x8_acc32_func2;
wire function_psimd_u_abs8_accxlen_func0;
wire function_psimd_u_abs8_accxlen_func1;
wire function_psimd_s_mul16x16_out64;
wire function_psimd_u_mul16x16_out64;
wire function_psimd_s_mul8x8_out64;
wire function_psimd_u_mul8x8_out64;
wire function_psimd_u_mul32x32_out64;
wire function_psimd_s_mul32x32_out64;
wire function_64p_s_add64;
wire function_64p_u_add64;
wire function_64p_s_sub64;
wire function_64p_u_sub64;
wire function_64p_s_mul32x32_acc64_func0;
wire function_64p_u_mul32x32_acc64_func0;
wire function_64p_s_mul32x32_acc64_func1;
wire function_64p_u_mul32x32_acc64_func1;
wire function_64p_s_mul16x16_acc64_func0;
wire function_64p_s_mul16x16_acc64_func1;
wire function_64p_s_mul16x16_acc64_func2;
wire function_64p_s_mul16x16_acc64_func3;
wire function_nsimd_s_addxlen;
wire function_nsimd_u_addxlen;
wire function_nsimd_s_subxlen;
wire function_nsimd_u_subxlen;
wire function_nsimd_s_mul16x16;
wire function_nsimd_s_mul16x16_double32;
wire function_nsimd_s_slra32;
wire function_nsimd_s_mul16x16_double32_acc32;
wire function_nsimd_s_avexlen;
wire function_simd_s_add32;
wire function_simd_u_add32;
wire function_simd_s_sub32;
wire function_simd_u_sub32;
wire function_simd_s_as32;
wire function_simd_u_as32;
wire function_simd_s_sa32;
wire function_simd_u_sa32;
wire function_simd_s_sra32;
wire function_simd_u_srl32;
wire function_simd_s_sll32;
wire function_simd_s_slra32;
wire function_simd_s_min32;
wire function_simd_u_min32;
wire function_simd_s_max32;
wire function_simd_u_max32;
wire function_simd_s_abs32;
wire function_nsimd_s_sra32;
wire function_psimd_s_mul32x32_acc64_func0;
wire function_psimd_s_mul32x32_acc64_func1;
wire function_psimd_s_mul32x32_acc64_func2;
wire function_psimd_s_mul32x32_acc64_func3;
wire function_psimd_s_mul32x32_acc64_func4;
wire function_psimd_s_mul32x32_acc64_func5;
wire function_psimd_s_mul32x32_acc64_func6;
wire function_psimd_s_pk32;
wire result_simd_s_wrap16;
wire result_simd_s_halve16;
wire result_simd_u_halve16;
wire result_simd_s_sat16;
wire result_simd_u_sat16;
wire result_simd_s_rnd16;
wire result_simd_s_rndsat16;
wire result_simd_s_wrap8;
wire result_simd_s_halve8;
wire result_simd_u_halve8;
wire result_simd_s_sat8;
wire result_simd_u_sat8;
wire result_simd_s_rnd8;
wire result_simd_s_rndsat8;
wire result_simd_s_unpk8;
wire result_psimd_s_halve32_sexlen;
wire result_psimd_u_halve32_sexlen;
wire result_psimd_s_rndxlen;
wire result_psimd_s_sat32_sexlen;
wire result_psimd_s_bypass32_sexlen;
wire result_psimd_s_cmpsel32_sexlen;
wire result_simd_s_bypass32;
wire result_simd_s_rnd32;
wire result_simd_s_sat32;
wire result_simd_s_rnd32_sat32;
wire result_psimd_s_sat32;
wire result_64p_s_wrap64;
wire result_64p_s_halve64;
wire result_64p_u_halve64;
wire result_64p_s_sat64;
wire result_64p_u_sat64;
wire result_nsimd_s_sat16_sexlen;
wire result_nsimd_u_sat16_sexlen;
wire result_nsimd_s_sat32_sexlen;
wire result_nsimd_u_sat32_sexlen;
wire result_nsimd_s_rndsat32_sexlen;
wire result_nsimd_s_halvexlen;
wire result_simd_s_wrap32;
wire result_simd_s_halve32;
wire result_simd_u_halve32;
wire result_simd_u_sat32;
wire result_simd_s_rndsat32;
wire result_nsimd_s_rnd32_se64;
wire result_psimd_s_sat64;
wire result_nsimd_s_sat16_se32;
wire result_nsimd_s_sat32;
wire [63:0] dsp_src1_64b_sxlen;
wire [63:0] dsp_src2_64b_sxlen;
wire [63:0] dsp_src1_64b_simd;
wire [63:0] dsp_src2_64b_simd;
wire [63:0] dsp_src3_64b_simd;
wire [63:0] dsp_src1_64b_pair;
wire [63:0] dsp_src2_64b_pair;
wire [63:0] dsp_src3_64b_pair;
wire [31:0] dsp_src1_W1;
wire [31:0] dsp_src1_W0;
wire [31:0] dsp_src2_W1;
wire [31:0] dsp_src2_W0;
wire [15:0] dsp_src1_H3;
wire [15:0] dsp_src1_H2;
wire [15:0] dsp_src1_H1;
wire [15:0] dsp_src1_H0;
wire [15:0] dsp_src2_H3;
wire [15:0] dsp_src2_H2;
wire [15:0] dsp_src2_H1;
wire [15:0] dsp_src2_H0;
wire [7:0] dsp_src1_B7;
wire [7:0] dsp_src1_B6;
wire [7:0] dsp_src1_B5;
wire [7:0] dsp_src1_B4;
wire [7:0] dsp_src1_B3;
wire [7:0] dsp_src1_B2;
wire [7:0] dsp_src1_B1;
wire [7:0] dsp_src1_B0;
wire [7:0] dsp_src2_B7;
wire [7:0] dsp_src2_B6;
wire [7:0] dsp_src2_B5;
wire [7:0] dsp_src2_B4;
wire [7:0] dsp_src2_B3;
wire [7:0] dsp_src2_B2;
wire [7:0] dsp_src2_B1;
wire [7:0] dsp_src2_B0;
wire [7:0] dsp_src3_B7;
wire [7:0] dsp_src3_B6;
wire [7:0] dsp_src3_B5;
wire [7:0] dsp_src3_B4;
wire [7:0] dsp_src3_B3;
wire [7:0] dsp_src3_B2;
wire [7:0] dsp_src3_B1;
wire [7:0] dsp_src3_B0;
wire [31:0] dsp_clipmin_W;
wire [15:0] dsp_clipmin_H;
wire [7:0] dsp_clipmin_B;
wire [31:0] dsp_clipmax_W;
wire [15:0] dsp_clipmax_H;
wire [7:0] dsp_clipmax_B;
wire simd16_op1_bottom16_sel;
wire simd16_op1_top16_sel;
wire simd16_op1_smal_sel;
wire simd16_op2_bottom16_sel;
wire simd16_op2_top16_sel;
wire simd16_op2_clipmin_sel_H0;
wire simd16_op2_clipmax_sel_H0;
wire simd16_op2_clipmin_sel_H1;
wire simd16_op2_clipmax_sel_H1;
wire simd16_op2_clipmin_sel_H2;
wire simd16_op2_clipmax_sel_H2;
wire simd16_op2_clipmin_sel_H3;
wire simd16_op2_clipmax_sel_H3;
wire [15:0] simd16_op1_H0;
wire [15:0] simd16_op2_H0;
wire [15:0] simd16_op1_H1;
wire [15:0] simd16_op2_H1;
wire [15:0] simd16_op1_H2;
wire [15:0] simd16_op2_H2;
wire [15:0] simd16_op1_H3;
wire [15:0] simd16_op2_H3;
wire [15:0] simd16_mul_op1_H0;
wire [15:0] simd16_mul_op2_H0;
wire [15:0] simd16_mul_op1_H1;
wire [15:0] simd16_mul_op2_H1;
wire [15:0] simd16_mul_op1_H2;
wire [15:0] simd16_mul_op2_H2;
wire [15:0] simd16_mul_op1_H3;
wire [15:0] simd16_mul_op2_H3;
wire simd16_addcmp_se1_H0;
wire simd16_addcmp_se1_H1;
wire simd16_addcmp_se1_H2;
wire simd16_addcmp_se1_H3;
wire simd16_addcmp_se2_H0;
wire simd16_addcmp_se2_H1;
wire simd16_addcmp_se2_H2;
wire simd16_addcmp_se2_H3;
wire simd16_addcmp_neg1_H0;
wire simd16_addcmp_neg1_H1;
wire simd16_addcmp_neg1_H2;
wire simd16_addcmp_neg1_H3;
wire simd16_addcmp_neg2_H0;
wire simd16_addcmp_neg2_H1;
wire simd16_addcmp_neg2_H2;
wire simd16_addcmp_neg2_H3;
wire [17:0] simd16_addcmp_out_H0;
wire [17:0] simd16_addcmp_out_H1;
wire [17:0] simd16_addcmp_out_H2;
wire [17:0] simd16_addcmp_out_H3;
wire simd16_addcmp_wrap;
wire simd16_addcmp_halve;
wire simd16_addcmp_s_sat;
wire simd16_addcmp_u_sat;
wire [16:0] simd16_addcmp_result_H0;
wire [16:0] simd16_addcmp_result_H1;
wire [16:0] simd16_addcmp_result_H2;
wire [16:0] simd16_addcmp_result_H3;
wire [63:0] simd16_addcmp_result_64b;
wire simd16_addcmp_ovf_set;
wire [16:0] simd16_shift_result_H0;
wire [16:0] simd16_shift_result_H1;
wire [16:0] simd16_shift_result_H2;
wire [16:0] simd16_shift_result_H3;
wire [63:0] simd16_shift_result_64b;
wire simd16_shift_ovf_set;
wire simd16_mul_se1_H0;
wire simd16_mul_se1_H1;
wire simd16_mul_se1_H2;
wire simd16_mul_se1_H3;
wire simd16_mul_se2_H0;
wire simd16_mul_se2_H1;
wire simd16_mul_se2_H2;
wire simd16_mul_se2_H3;
wire [31:0] simd16_mul_out_H0;
wire [31:0] simd16_mul_out_H1;
wire [31:0] simd16_mul_out_H2;
wire [31:0] simd16_mul_out_H3;
wire simd16_mul_s_sat;
wire [16:0] simd16_mul_result_H0;
wire [16:0] simd16_mul_result_H1;
wire [16:0] simd16_mul_result_H2;
wire [16:0] simd16_mul_result_H3;
wire [63:0] simd16_mul_result_64b;
wire simd16_mul_ovf_set;
wire [63:0] simd16_swap_result_64b;
wire simd16_swap_ovf_set;
wire [15:0] simd16_clz_result_H0;
wire [15:0] simd16_clz_result_H1;
wire [15:0] simd16_clz_result_H2;
wire [15:0] simd16_clz_result_H3;
wire [63:0] simd16_clz_result_64b;
wire simd16_clz_ovf_set;
wire simd16_result_addcmp_sel;
wire simd16_result_shift_sel;
wire simd16_result_mul_sel;
wire simd16_result_swap_sel;
wire simd16_result_clz_sel;
wire [63:0] stage1_simd16_final_result_64b;
wire stage1_simd16_final_ovf_set;
wire simd8_op1_base_sel;
wire simd8_op2_base_sel;
wire simd8_op2_cross_sel;
wire simd8_op2_clipmin_sel_B0;
wire simd8_op2_clipmax_sel_B0;
wire simd8_op2_clipmin_sel_B1;
wire simd8_op2_clipmax_sel_B1;
wire simd8_op2_clipmin_sel_B2;
wire simd8_op2_clipmax_sel_B2;
wire simd8_op2_clipmin_sel_B3;
wire simd8_op2_clipmax_sel_B3;
wire simd8_op2_clipmin_sel_B4;
wire simd8_op2_clipmax_sel_B4;
wire simd8_op2_clipmin_sel_B5;
wire simd8_op2_clipmax_sel_B5;
wire simd8_op2_clipmin_sel_B6;
wire simd8_op2_clipmax_sel_B6;
wire simd8_op2_clipmin_sel_B7;
wire simd8_op2_clipmax_sel_B7;
wire [7:0] simd8_op1_B0;
wire [7:0] simd8_op2_B0;
wire [7:0] simd8_op1_B1;
wire [7:0] simd8_op2_B1;
wire [7:0] simd8_op1_B2;
wire [7:0] simd8_op2_B2;
wire [7:0] simd8_op1_B3;
wire [7:0] simd8_op2_B3;
wire [7:0] simd8_op1_B4;
wire [7:0] simd8_op2_B4;
wire [7:0] simd8_op1_B5;
wire [7:0] simd8_op2_B5;
wire [7:0] simd8_op1_B6;
wire [7:0] simd8_op2_B6;
wire [7:0] simd8_op1_B7;
wire [7:0] simd8_op2_B7;
wire simd8_addcmp_se1_B0;
wire simd8_addcmp_se1_B1;
wire simd8_addcmp_se1_B2;
wire simd8_addcmp_se1_B3;
wire simd8_addcmp_se1_B4;
wire simd8_addcmp_se1_B5;
wire simd8_addcmp_se1_B6;
wire simd8_addcmp_se1_B7;
wire simd8_addcmp_se2_B0;
wire simd8_addcmp_se2_B1;
wire simd8_addcmp_se2_B2;
wire simd8_addcmp_se2_B3;
wire simd8_addcmp_se2_B4;
wire simd8_addcmp_se2_B5;
wire simd8_addcmp_se2_B6;
wire simd8_addcmp_se2_B7;
wire simd8_addcmp_neg1_B0;
wire simd8_addcmp_neg1_B1;
wire simd8_addcmp_neg1_B2;
wire simd8_addcmp_neg1_B3;
wire simd8_addcmp_neg1_B4;
wire simd8_addcmp_neg1_B5;
wire simd8_addcmp_neg1_B6;
wire simd8_addcmp_neg1_B7;
wire simd8_addcmp_neg2_B0;
wire simd8_addcmp_neg2_B1;
wire simd8_addcmp_neg2_B2;
wire simd8_addcmp_neg2_B3;
wire simd8_addcmp_neg2_B4;
wire simd8_addcmp_neg2_B5;
wire simd8_addcmp_neg2_B6;
wire simd8_addcmp_neg2_B7;
wire [9:0] simd8_addcmp_out_B0;
wire [9:0] simd8_addcmp_out_B1;
wire [9:0] simd8_addcmp_out_B2;
wire [9:0] simd8_addcmp_out_B3;
wire [9:0] simd8_addcmp_out_B4;
wire [9:0] simd8_addcmp_out_B5;
wire [9:0] simd8_addcmp_out_B6;
wire [9:0] simd8_addcmp_out_B7;
wire simd8_addcmp_wrap;
wire simd8_addcmp_halve;
wire simd8_addcmp_s_sat;
wire simd8_addcmp_u_sat;
wire [8:0] simd8_addcmp_result_B0;
wire [8:0] simd8_addcmp_result_B1;
wire [8:0] simd8_addcmp_result_B2;
wire [8:0] simd8_addcmp_result_B3;
wire [8:0] simd8_addcmp_result_B4;
wire [8:0] simd8_addcmp_result_B5;
wire [8:0] simd8_addcmp_result_B6;
wire [8:0] simd8_addcmp_result_B7;
wire [63:0] simd8_addcmp_result_64b;
wire simd8_addcmp_ovf_set;
wire [8:0] simd8_shift_result_B0;
wire [8:0] simd8_shift_result_B1;
wire [8:0] simd8_shift_result_B2;
wire [8:0] simd8_shift_result_B3;
wire [8:0] simd8_shift_result_B4;
wire [8:0] simd8_shift_result_B5;
wire [8:0] simd8_shift_result_B6;
wire [8:0] simd8_shift_result_B7;
wire [63:0] simd8_shift_result_64b;
wire simd8_shift_ovf_set;
wire simd8_mul_se1_B0;
wire simd8_mul_se1_B1;
wire simd8_mul_se1_B2;
wire simd8_mul_se1_B3;
wire simd8_mul_se1_B4;
wire simd8_mul_se1_B5;
wire simd8_mul_se1_B6;
wire simd8_mul_se1_B7;
wire simd8_mul_se2_B0;
wire simd8_mul_se2_B1;
wire simd8_mul_se2_B2;
wire simd8_mul_se2_B3;
wire simd8_mul_se2_B4;
wire simd8_mul_se2_B5;
wire simd8_mul_se2_B6;
wire simd8_mul_se2_B7;
wire [17:0] simd8_mul_out_B0;
wire [17:0] simd8_mul_out_B1;
wire [17:0] simd8_mul_out_B2;
wire [17:0] simd8_mul_out_B3;
wire [17:0] simd8_mul_out_B4;
wire [17:0] simd8_mul_out_B5;
wire [17:0] simd8_mul_out_B6;
wire [17:0] simd8_mul_out_B7;
wire simd8_mul_s_sat;
wire [8:0] simd8_mul_result_B0;
wire [8:0] simd8_mul_result_B1;
wire [8:0] simd8_mul_result_B2;
wire [8:0] simd8_mul_result_B3;
wire [8:0] simd8_mul_result_B4;
wire [8:0] simd8_mul_result_B5;
wire [8:0] simd8_mul_result_B6;
wire [8:0] simd8_mul_result_B7;
wire [63:0] simd8_mul_result_64b;
wire simd8_mul_ovf_set;
wire [63:0] simd8_swap_result_64b;
wire simd8_swap_ovf_set;
wire [7:0] simd8_clz_result_B0;
wire [7:0] simd8_clz_result_B1;
wire [7:0] simd8_clz_result_B2;
wire [7:0] simd8_clz_result_B3;
wire [7:0] simd8_clz_result_B4;
wire [7:0] simd8_clz_result_B5;
wire [7:0] simd8_clz_result_B6;
wire [7:0] simd8_clz_result_B7;
wire [63:0] simd8_clz_result_64b;
wire simd8_clz_ovf_set;
wire simd8_unpack_en1_H0;
wire simd8_unpack_en2_H0;
wire simd8_unpack_en3_H0;
wire simd8_unpack_en1_H1;
wire simd8_unpack_en2_H1;
wire simd8_unpack_en3_H1;
wire simd8_unpack_en1_H2;
wire simd8_unpack_en2_H2;
wire simd8_unpack_en3_H2;
wire simd8_unpack_en1_H3;
wire simd8_unpack_en2_H3;
wire simd8_unpack_en3_H3;
wire [15:0] simd8_unpack_result_H0;
wire [15:0] simd8_unpack_result_H1;
wire [15:0] simd8_unpack_result_H2;
wire [15:0] simd8_unpack_result_H3;
wire [63:0] simd8_unpack_result_64b;
wire simd8_unpack_ovf_set;
wire simd8_result_addcmp_sel;
wire simd8_result_shift_sel;
wire simd8_result_mul_sel;
wire simd8_result_swap_sel;
wire simd8_result_clz_sel;
wire simd8_result_unpack_sel;
wire [63:0] stage1_simd8_final_result_64b;
wire stage1_simd8_final_ovf_set;
wire psimd32_op1_base_sel;
wire psimd32_op1_top32_sel;
wire psimd32_op2_base_sel;
wire psimd32_op2_top32_sel;
wire psimd32_op2_clipmin_sel_W0;
wire psimd32_op2_clipmax_sel_W0;
wire psimd32_op2_clipmin_sel_W1;
wire psimd32_op2_clipmax_sel_W1;
wire psimd32_op2_bottom16_sel;
wire psimd32_op2_top16_sel;
wire [31:0] psimd32_op1_W0;
wire [31:0] psimd32_op2_W0;
wire [31:0] psimd32_op1_W1;
wire [31:0] psimd32_op2_W1;
wire [63:0] psimd32_pack_result_64b;
wire psimd32_pack_ovf_set;
wire psimd32_addcmp_se1_W0;
wire psimd32_addcmp_se1_W1;
wire psimd32_addcmp_se2_W0;
wire psimd32_addcmp_se2_W1;
wire psimd32_addcmp_neg1_W0;
wire psimd32_addcmp_neg1_W1;
wire psimd32_addcmp_neg2_W0;
wire psimd32_addcmp_neg2_W1;
wire [33:0] psimd32_addcmp_out_W0;
wire [33:0] psimd32_addcmp_out_W1;
wire psimd32_addcmp_min;
wire psimd32_addcmp_max;
wire psimd32_addcmp_clip;
wire psimd32_addcmp_wrap;
wire psimd32_addcmp_halve;
wire psimd32_addcmp_s_sat;
wire psimd32_addcmp_u_sat;
wire [32:0] psimd32_addcmp_result_W0;
wire [32:0] psimd32_addcmp_result_W1;
wire psimd32_addcmp_result32sexlen;
wire [63:0] psimd32_addcmp_result_64b;
wire psimd32_addcmp_ovf_set;
wire [31:0] psimd32_clz_result_W0;
wire [31:0] psimd32_clz_result_W1;
wire [63:0] psimd32_clz_result_64b;
wire psimd32_clz_ovf_set;
wire psimd32_mul_se1_W0;
wire psimd32_mul_se2_W0;
wire psimd32_mul_se1_W1;
wire psimd32_mul_se2_W1;
wire psimd32_mul_32x16;
wire psimd32_mul_no_opovf;
wire [66:0] psimd32_mul_lv1_wt_sum_W0;
wire [66:0] psimd32_mul_lv1_wt_cout_W0;
wire [134:0] psimd32_mul_lv1_out_W0;
wire [66:0] psimd32_mul_lv1_wt_sum_W1;
wire [66:0] psimd32_mul_lv1_wt_cout_W1;
wire [134:0] psimd32_mul_lv1_out_W1;
wire stage2_psimd32_mul_data_en;
wire [16:0] stage2_psimd32_mul_fctrl_nx;
wire [4:0] stage2_psimd32_mul_rctrl_nx;
reg [16:0] stage2_psimd32_mul_fctrl;
reg [4:0] stage2_psimd32_mul_rctrl;
wire [64:0] stage2_psimd32_mul_result_W0;
wire [64:0] stage2_psimd32_mul_result_W1;
wire [175:0] stage2_psimd32_mul_lv1_result_W0_nx;
wire [175:0] stage2_psimd32_mul_lv1_result_W1_nx;
reg [175:0] stage2_psimd32_mul_lv1_result_W0;
reg [175:0] stage2_psimd32_mul_lv1_result_W1;
wire stage2_psimd32_mul_result32sexlen;
wire stage2_psimd32_mul_resultout64;
wire [63:0] stage2_psimd32_mul_result_64b;
wire stage2_psimd32_mul_ovf_set;
wire stage3_psimd32_mul_data_en;
wire [5:0] stage3_psimd32_mul_fctrl_nx;
wire [1:0] stage3_psimd32_mul_rctrl_nx;
wire [66:0] stage3_psimd32_mul_out1_nx;
wire [66:0] stage3_psimd32_mul_out2_nx;
reg [5:0] stage3_psimd32_mul_fctrl;
reg [1:0] stage3_psimd32_mul_rctrl;
reg [66:0] stage3_psimd32_mul_out1;
reg [66:0] stage3_psimd32_mul_out2;
wire [63:0] stage3_psimd32_mul_result_64b;
wire stage3_psimd32_mul_ovf_set;
wire psimd32_result_addcmp_sel;
wire psimd32_result_clz_sel;
wire psimd32_result_pack_sel;
wire stage2_psimd32_result_mul_sel;
wire stage3_psimd32_result_mul_sel;
wire [63:0] stage1_psimd32_final_result_64b;
wire stage1_psimd32_final_ovf_set;
wire [63:0] stage2_psimd32_final_result_64b;
wire stage2_psimd32_final_ovf_set;
wire [63:0] stage3_psimd32_final_result_64b;
wire stage3_psimd32_final_ovf_set;
wire psimdxlen_op1_base_sel;
wire psimdxlen_op1_pair_sel;
wire psimdxlen_op2_base_sel;
wire psimdxlen_op2_pair_sel;
wire psimdxlen_op3_base_sel;
wire [63:0] psimdxlen_op1_64b;
wire [63:0] psimdxlen_op2_64b;
wire [63:0] psimdxlen_op3_64b;
wire psimdxlen_shift_s_rnd;
wire psimdxlen_shift_s_sat;
wire [64:0] psimdxlen_shift_result_W0XLEN;
wire [64:0] psimdxlen_shift_result_W1;
wire psimdxlen_shift_result32;
wire [63:0] psimdxlen_shift_result_64b;
wire psimdxlen_shift_ovf_set;
reg [63:0] psimdxlen_bpick_result_64b;
wire psimdxlen_bpick_ovf_set;
wire [7:0] psimdxlen_insb_byte_sel;
wire [7:0] psimdxlen_insb_result_B0;
wire [7:0] psimdxlen_insb_result_B1;
wire [7:0] psimdxlen_insb_result_B2;
wire [7:0] psimdxlen_insb_result_B3;
wire [7:0] psimdxlen_insb_result_B4;
wire [7:0] psimdxlen_insb_result_B5;
wire [7:0] psimdxlen_insb_result_B6;
wire [7:0] psimdxlen_insb_result_B7;
wire [63:0] psimdxlen_insb_result_64b;
wire psimdxlen_insb_ovf_set;
wire psimdxlen_result_shift_sel;
wire psimdxlen_result_bpick_sel;
wire psimdxlen_result_insb_sel;
wire [63:0] stage1_psimdxlen_final_result_64b;
wire stage1_psimdxlen_final_ovf_set;
wire psimd16_op1_bottom_sel;
wire psimd16_op1_top_sel;
wire psimd16_op2_bottom_sel;
wire psimd16_op2_top_sel;
wire [15:0] psimd16_op1_H0;
wire [15:0] psimd16_op2_H0;
wire [15:0] psimd16_op1_H2;
wire [15:0] psimd16_op2_H2;
wire [63:0] psimd16_pack_result_64b;
wire psimd16_pack_ovf_set;
wire psimd16_result_pack_sel;
wire [31:0] stage1_psimd16_mul_out_H0;
wire [31:0] stage1_psimd16_mul_out_H1;
wire [31:0] stage1_psimd16_mul_out_H2;
wire [31:0] stage1_psimd16_mul_out_H3;
wire stage1_is_mul16x16_out64;
wire [63:0] stage1_psimd16_mul_result_64b;
wire stage1_psimd16_mul_ovf_set;
wire stage2_psimd16_mul_data_en;
wire [10:0] stage2_psimd16_mul_fctrl_nx;
wire [1:0] stage2_psimd16_mul_rctrl_nx;
wire [31:0] stage2_psimd16_mul_out_H0_nx;
wire [31:0] stage2_psimd16_mul_out_H1_nx;
wire [31:0] stage2_psimd16_mul_out_H2_nx;
wire [31:0] stage2_psimd16_mul_out_H3_nx;
wire stage2_psimd16_opovf_H0_nx;
wire stage2_psimd16_opovf_H2_nx;
reg [10:0] stage2_psimd16_mul_fctrl;
reg [1:0] stage2_psimd16_mul_rctrl;
reg [31:0] stage2_psimd16_mul_out_H0;
reg [31:0] stage2_psimd16_mul_out_H1;
reg [31:0] stage2_psimd16_mul_out_H2;
reg [31:0] stage2_psimd16_mul_out_H3;
reg stage2_psimd16_opovf_H0;
reg stage2_psimd16_opovf_H2;
wire [34:0] stage2_psimd16_mul_result_W0;
wire [34:0] stage2_psimd16_mul_result_W1;
wire stage2_psimd16_mul_result32sexlen;
wire [63:0] stage2_psimd16_mul_result_64b;
wire stage2_psimd16_mul_ovf_set;
wire stage3_psimd16_mul_data_en;
wire [3:0] stage3_psimd16_mul_fctrl_nx;
wire stage3_psimd16_mul_rctrl_nx;
wire [33:0] stage3_psimd16_mul_out_W0_nx;
wire [33:0] stage3_psimd16_mul_out_W1_nx;
reg [3:0] stage3_psimd16_mul_fctrl;
reg stage3_psimd16_mul_rctrl;
reg [33:0] stage3_psimd16_mul_out_W0;
reg [33:0] stage3_psimd16_mul_out_W1;
wire [63:0] stage3_psimd16_mul_result_64b;
wire stage3_psimd16_mul_ovf_set;
wire stage1_psimd16_result_mul_sel;
wire stage2_psimd16_result_mul_sel;
wire stage3_psimd16_result_mul_sel;
wire [63:0] stage1_psimd16_final_result_64b;
wire stage1_psimd16_final_ovf_set;
wire [63:0] stage2_psimd16_final_result_64b;
wire stage2_psimd16_final_ovf_set;
wire [63:0] stage3_psimd16_final_result_64b;
wire stage3_psimd16_final_ovf_set;
wire function_psimd_s_mul8x8_acc32;
wire [39:0] stage1_psimd8_mul_out_W0;
wire [39:0] stage1_psimd8_mul_out_W1;
wire [63:0] stage1_psimd8_mul_result_64b;
wire stage1_psimd8_mul_ovf_set;
wire [23:0] stage1_psimd8_pbsad_out_W0;
wire [23:0] stage1_psimd8_pbsad_out_W1;
wire [23:0] stage1_psimd8_pbsad_out_64b;
wire stage2_psimd8_pbsad_data_en;
wire [1:0] stage2_psimd8_pbsad_fctrl_nx;
wire [23:0] stage2_psimd8_pbsad_out_nx;
reg [1:0] stage2_psimd8_pbsad_fctrl;
reg [23:0] stage2_psimd8_pbsad_out;
wire [31:0] stage2_psimd8_pbsad_out_xlen;
wire [63:0] stage2_psimd8_pbsad_result_64b;
wire stage1_psimd8_result_mul_sel;
wire [63:0] stage1_psimd8_final_result_64b;
wire stage1_psimd8_final_ovf_set;
wire stage2_psimd8_pbsad_ovf_set;
wire stage2_psimd8_result_pbsad_sel;
wire [63:0] stage2_psimd8_final_result_64b;
wire stage2_psimd8_final_ovf_set;
wire profile64_op1_base_sel;
wire profile64_op2_base_sel;
wire profile64_op1_sxlen_sel;
wire profile64_op2_sxlen_sel;
wire profile64_op1_s32_sel;
wire profile64_op2_s32_sel;
wire profile64_op1_u32_sel;
wire profile64_op2_u32_sel;
wire [63:0] profile64_op1_64b;
wire [63:0] profile64_op2_64b;
wire profile64_add_se1_64b;
wire profile64_add_se2_64b;
wire profile64_add_neg1_64b;
wire profile64_add_neg2_64b;
wire [64:0] profile64_add_out_64b;
wire [7:0] profile64_add_rctrl;
wire [63:0] profile64_add_result_64b;
wire profile64_add_ovf_set;
wire profile64_result_add_sel;
wire [66:0] stage2_profile64_mul_csa_out1;
wire [66:0] stage2_profile64_mul_csa_out2;
wire stage3_profile64_msr64;
wire stage3_profile64_s_sat64;
wire stage3_profile64_u_sat64;
wire [63:0] stage3_profile64_mul_result_64b;
wire stage3_profile64_mul_ovf_set;
wire [63:0] stage1_profile64_final_result_64b;
wire stage1_profile64_final_ovf_set;
wire nsimd16_mul_s_sat16;
wire nsimd16_mul_s_sat32;
wire [32:0] nsimd16_mul_result_H0;
wire [32:0] nsimd16_mul_result_H2;
wire nsimd16_mul_resultsexlen;
wire [63:0] stage1_nsimd16_mul_result_64b;
wire stage1_nsimd16_mul_ovf_set;
wire stage1_nsimd16_result_mul_sel;
wire [63:0] stage1_nsimd16_final_result_64b;
wire stage1_nsimd16_final_ovf_set;
wire stage2_dsp_ctrl_en;
wire stage3_dsp_ctrl_en;
wire stage1_dsp_ivalid;
reg stage2_dsp_ivalid;
wire stage1_dsp_ovfset;
reg stage2_dsp_ovfset;
reg stage3_dsp_ovfset;
wire acc_din_base_sel;
wire acc_din_smal_sel;
wire [31:0] stage1_acc_din_W0;
wire [31:0] stage1_acc_din_W1;
wire stage2_acc_din_en;
wire [31:0] stage2_acc_din_W0_nx;
wire [31:0] stage2_acc_din_W1_nx;
wire stage2_acc_din_sign_nx;
reg [31:0] stage2_acc_din_W0;
reg [31:0] stage2_acc_din_W1;
reg stage2_acc_din_sign;
wire [63:0] stage2_acc_din_64b;
wire stage3_acc_din_en;
wire [31:0] stage3_acc_din_W0_nx;
wire [31:0] stage3_acc_din_W1_nx;
reg [31:0] stage3_acc_din_W0;
reg [31:0] stage3_acc_din_W1;
wire stage1_xsimd16_result_mul_sel;
wire [63:0] stage1_xsimd16_mul_result_64b;
wire stage1_xsimd16_mul_ovf_set;
reg stage2_xsimd16_result_mul_sel;
reg [63:0] stage2_xsimd16_mul_result_64b;
reg stage2_xsimd16_mul_ovf_set;
wire [63:0] stage2_xsimd16_final_result_64b;
wire stage2_xsimd16_final_ovf_set;
wire stage2_xsimd16_mul_data_en;
assign operand_simd_op16 = dsp_operand_ctrl[0];
assign operand_simd_cross_op16 = dsp_operand_ctrl[1];
assign operand_simd_clip_op16 = dsp_operand_ctrl[2];
assign operand_simd_op8 = dsp_operand_ctrl[3];
assign operand_simd_clip_op8 = dsp_operand_ctrl[4];
assign operand_simd_cross_op8 = dsp_operand_ctrl[5];
assign operand_psimd_op32 = dsp_operand_ctrl[6];
assign operand_psimd_opxlen = dsp_operand_ctrl[7];
assign operand_psimd_op16b_op16b = dsp_operand_ctrl[8];
assign operand_psimd_op16b_op16t = dsp_operand_ctrl[9];
assign operand_psimd_op16t_op16b = dsp_operand_ctrl[10];
assign operand_psimd_op16t_op16t = dsp_operand_ctrl[11];
assign operand_psimd_clip_op32 = dsp_operand_ctrl[12];
assign operand_psimd_op64 = dsp_operand_ctrl[13];
assign operand_psimd_op32_op16b = dsp_operand_ctrl[14];
assign operand_psimd_op32_op16t = dsp_operand_ctrl[15];
assign operand_psimd_op16 = dsp_operand_ctrl[16];
assign operand_psimd_cross_op16 = dsp_operand_ctrl[17];
assign operand_psimd_reverse_op16 = dsp_operand_ctrl[18];
assign operand_psimd_smal_op16 = dsp_operand_ctrl[19];
assign operand_psimd_op8 = dsp_operand_ctrl[20];
assign operand_psimd_cross_op8 = dsp_operand_ctrl[21];
assign operand_64p_opxlen = dsp_operand_ctrl[22];
assign operand_64p_op16b_op16b = dsp_operand_ctrl[23];
assign operand_64p_op16b_op16t = dsp_operand_ctrl[24];
assign operand_64p_op16t_op16t = dsp_operand_ctrl[25];
assign operand_64p_op16 = dsp_operand_ctrl[26];
assign operand_64p_cross_op16 = dsp_operand_ctrl[27];
assign operand_64p_reverse_op16 = dsp_operand_ctrl[28];
assign operand_nsimd_s_op32_sexlen = dsp_operand_ctrl[29];
assign operand_nsimd_u_op32_sexlen = dsp_operand_ctrl[30];
assign operand_nsimd_op16b_op16b = dsp_operand_ctrl[31];
assign operand_nsimd_op16b_op16t = dsp_operand_ctrl[32];
assign operand_nsimd_op16t_op16t = dsp_operand_ctrl[33];
assign operand_nsimd_op32 = dsp_operand_ctrl[34];
assign operand_nsimd_opxlen = dsp_operand_ctrl[35];
assign operand_simd_op32 = dsp_operand_ctrl[36];
assign operand_simd_cross_op32 = dsp_operand_ctrl[37];
assign operand_psimd_op32b_op32b = dsp_operand_ctrl[38];
assign operand_psimd_op32b_op32t = dsp_operand_ctrl[39];
assign operand_psimd_op32t_op32t = dsp_operand_ctrl[40];
assign operand_psimd_cross_op32 = dsp_operand_ctrl[41];
assign operand_psimd_reverse_op32 = dsp_operand_ctrl[42];
assign operand_psimd_op32t_op32b = dsp_operand_ctrl[43];
assign function_simd_s_add16 = dsp_function_ctrl[0];
assign function_simd_u_add16 = dsp_function_ctrl[1];
assign function_simd_s_sub16 = dsp_function_ctrl[2];
assign function_simd_u_sub16 = dsp_function_ctrl[3];
assign function_simd_s_as16 = dsp_function_ctrl[4];
assign function_simd_u_as16 = dsp_function_ctrl[5];
assign function_simd_s_sa16 = dsp_function_ctrl[6];
assign function_simd_u_sa16 = dsp_function_ctrl[7];
assign function_simd_s_sra16 = dsp_function_ctrl[8];
assign function_simd_u_srl16 = dsp_function_ctrl[9];
assign function_simd_s_sll16 = dsp_function_ctrl[10];
assign function_simd_s_slra16 = dsp_function_ctrl[11];
assign function_simd_s_cmpeq16 = dsp_function_ctrl[12];
assign function_simd_s_cmplt16 = dsp_function_ctrl[13];
assign function_simd_u_cmplt16 = dsp_function_ctrl[14];
assign function_simd_s_cmple16 = dsp_function_ctrl[15];
assign function_simd_u_cmple16 = dsp_function_ctrl[16];
assign function_simd_s_min16 = dsp_function_ctrl[17];
assign function_simd_u_min16 = dsp_function_ctrl[18];
assign function_simd_s_max16 = dsp_function_ctrl[19];
assign function_simd_u_max16 = dsp_function_ctrl[20];
assign function_simd_s_abs16 = dsp_function_ctrl[21];
assign function_simd_s_clip16 = dsp_function_ctrl[22];
assign function_simd_s_mul16 = dsp_function_ctrl[23];
assign function_simd_s_swap16 = dsp_function_ctrl[24];
assign function_simd_s_clz16 = dsp_function_ctrl[25];
assign function_simd_s_clo16 = dsp_function_ctrl[26];
assign function_simd_s_clrs16 = dsp_function_ctrl[27];
assign function_simd_s_add8 = dsp_function_ctrl[28];
assign function_simd_u_add8 = dsp_function_ctrl[29];
assign function_simd_s_sub8 = dsp_function_ctrl[30];
assign function_simd_u_sub8 = dsp_function_ctrl[31];
assign function_simd_s_sra8 = dsp_function_ctrl[32];
assign function_simd_u_srl8 = dsp_function_ctrl[33];
assign function_simd_s_sll8 = dsp_function_ctrl[34];
assign function_simd_s_slra8 = dsp_function_ctrl[35];
assign function_simd_s_cmpeq8 = dsp_function_ctrl[36];
assign function_simd_s_cmplt8 = dsp_function_ctrl[37];
assign function_simd_u_cmplt8 = dsp_function_ctrl[38];
assign function_simd_s_cmple8 = dsp_function_ctrl[39];
assign function_simd_u_cmple8 = dsp_function_ctrl[40];
assign function_simd_s_min8 = dsp_function_ctrl[41];
assign function_simd_u_min8 = dsp_function_ctrl[42];
assign function_simd_s_max8 = dsp_function_ctrl[43];
assign function_simd_u_max8 = dsp_function_ctrl[44];
assign function_simd_s_abs8 = dsp_function_ctrl[45];
assign function_simd_s_clip8 = dsp_function_ctrl[46];
assign function_simd_s_mul8 = dsp_function_ctrl[47];
assign function_simd_s_swap8 = dsp_function_ctrl[48];
assign function_simd_s_clz8 = dsp_function_ctrl[49];
assign function_simd_s_clo8 = dsp_function_ctrl[50];
assign function_simd_s_clrs8 = dsp_function_ctrl[51];
assign function_simd_s_unpk8_10 = dsp_function_ctrl[52];
assign function_simd_s_unpk8_20 = dsp_function_ctrl[53];
assign function_simd_s_unpk8_30 = dsp_function_ctrl[54];
assign function_simd_s_unpk8_31 = dsp_function_ctrl[55];
assign function_simd_s_unpk8_32 = dsp_function_ctrl[56];
assign function_psimd_s_add32 = dsp_function_ctrl[57];
assign function_psimd_u_add32 = dsp_function_ctrl[58];
assign function_psimd_s_sub32 = dsp_function_ctrl[59];
assign function_psimd_u_sub32 = dsp_function_ctrl[60];
assign function_psimd_s_sraxlen = dsp_function_ctrl[61];
assign function_psimd_s_sll32 = dsp_function_ctrl[62];
assign function_psimd_s_pk16 = dsp_function_ctrl[63];
assign function_psimd_s_clip32 = dsp_function_ctrl[64];
assign function_psimd_u_bitrevxlen = dsp_function_ctrl[65];
assign function_psimd_s_wext32 = dsp_function_ctrl[66];
assign function_psimd_s_bpickxlen = dsp_function_ctrl[67];
assign function_psimd_s_insbxlen = dsp_function_ctrl[68];
assign function_psimd_s_min32 = dsp_function_ctrl[69];
assign function_psimd_s_max32 = dsp_function_ctrl[70];
assign function_psimd_s_abs32 = dsp_function_ctrl[71];
assign function_psimd_s_clz32 = dsp_function_ctrl[72];
assign function_psimd_s_clo32 = dsp_function_ctrl[73];
assign function_psimd_s_clrs32 = dsp_function_ctrl[74];
assign function_psimd_s_mul32x32_acc32_func0 = dsp_function_ctrl[75];
assign function_psimd_s_mul32x32_acc32_func1 = dsp_function_ctrl[76];
assign function_psimd_s_mul32x32_acc32_func2 = dsp_function_ctrl[77];
assign function_psimd_s_mul32x32_acc32_func3 = dsp_function_ctrl[78];
assign function_psimd_s_mul32x32_acc32_func4 = dsp_function_ctrl[79];
assign function_psimd_s_mul32x32_acc32_func5 = dsp_function_ctrl[80];
assign function_psimd_s_mul32x16_acc32_func0 = dsp_function_ctrl[81];
assign function_psimd_s_mul32x16_acc32_func1 = dsp_function_ctrl[82];
assign function_psimd_s_mul32x16_acc32_func2 = dsp_function_ctrl[83];
assign function_psimd_s_mul32x16_acc32_func3 = dsp_function_ctrl[84];
assign function_psimd_s_mul16x16_acc32_func0 = dsp_function_ctrl[85];
assign function_psimd_s_mul16x16_acc32_func1 = dsp_function_ctrl[86];
assign function_psimd_s_mul16x16_acc32_func2 = dsp_function_ctrl[87];
assign function_psimd_s_mul16x16_acc32_func3 = dsp_function_ctrl[88];
assign function_psimd_s_mul16x16_acc32_func4 = dsp_function_ctrl[89];
assign function_psimd_s_mul16x16_acc32_func5 = dsp_function_ctrl[90];
assign function_psimd_s_mul16x16_acc32_func6 = dsp_function_ctrl[91];
assign function_psimd_s_mul16x16_acc64_func0 = dsp_function_ctrl[92];
assign function_psimd_s_mul8x8_acc32_func0 = dsp_function_ctrl[93];
assign function_psimd_s_mul8x8_acc32_func1 = dsp_function_ctrl[94];
assign function_psimd_s_mul8x8_acc32_func2 = dsp_function_ctrl[95];
assign function_psimd_u_abs8_accxlen_func0 = dsp_function_ctrl[96];
assign function_psimd_u_abs8_accxlen_func1 = dsp_function_ctrl[97];
assign function_psimd_s_mul16x16_out64 = dsp_function_ctrl[98];
assign function_psimd_u_mul16x16_out64 = dsp_function_ctrl[99];
assign function_psimd_s_mul8x8_out64 = dsp_function_ctrl[100];
assign function_psimd_u_mul8x8_out64 = dsp_function_ctrl[101];
assign function_psimd_u_mul32x32_out64 = dsp_function_ctrl[102];
assign function_psimd_s_mul32x32_out64 = dsp_function_ctrl[103];
assign function_64p_s_add64 = dsp_function_ctrl[104];
assign function_64p_u_add64 = dsp_function_ctrl[105];
assign function_64p_s_sub64 = dsp_function_ctrl[106];
assign function_64p_u_sub64 = dsp_function_ctrl[107];
assign function_64p_s_mul32x32_acc64_func0 = dsp_function_ctrl[108];
assign function_64p_u_mul32x32_acc64_func0 = dsp_function_ctrl[109];
assign function_64p_s_mul32x32_acc64_func1 = dsp_function_ctrl[110];
assign function_64p_u_mul32x32_acc64_func1 = dsp_function_ctrl[111];
assign function_64p_s_mul16x16_acc64_func0 = dsp_function_ctrl[112];
assign function_64p_s_mul16x16_acc64_func1 = dsp_function_ctrl[113];
assign function_64p_s_mul16x16_acc64_func2 = dsp_function_ctrl[114];
assign function_64p_s_mul16x16_acc64_func3 = dsp_function_ctrl[115];
assign function_nsimd_s_addxlen = dsp_function_ctrl[116];
assign function_nsimd_u_addxlen = dsp_function_ctrl[117];
assign function_nsimd_s_subxlen = dsp_function_ctrl[118];
assign function_nsimd_u_subxlen = dsp_function_ctrl[119];
assign function_nsimd_s_mul16x16 = dsp_function_ctrl[120];
assign function_nsimd_s_mul16x16_double32 = dsp_function_ctrl[121];
assign function_nsimd_s_slra32 = dsp_function_ctrl[122];
assign function_nsimd_s_mul16x16_double32_acc32 = dsp_function_ctrl[123];
assign function_nsimd_s_avexlen = dsp_function_ctrl[124];
assign function_simd_s_add32 = dsp_function_ctrl[125];
assign function_simd_u_add32 = dsp_function_ctrl[126];
assign function_simd_s_sub32 = dsp_function_ctrl[127];
assign function_simd_u_sub32 = dsp_function_ctrl[128];
assign function_simd_s_as32 = dsp_function_ctrl[129];
assign function_simd_u_as32 = dsp_function_ctrl[130];
assign function_simd_s_sa32 = dsp_function_ctrl[131];
assign function_simd_u_sa32 = dsp_function_ctrl[132];
assign function_simd_s_sra32 = dsp_function_ctrl[133];
assign function_simd_u_srl32 = dsp_function_ctrl[134];
assign function_simd_s_sll32 = dsp_function_ctrl[135];
assign function_simd_s_slra32 = dsp_function_ctrl[136];
assign function_simd_s_min32 = dsp_function_ctrl[137];
assign function_simd_u_min32 = dsp_function_ctrl[138];
assign function_simd_s_max32 = dsp_function_ctrl[139];
assign function_simd_u_max32 = dsp_function_ctrl[140];
assign function_simd_s_abs32 = dsp_function_ctrl[141];
assign function_nsimd_s_sra32 = dsp_function_ctrl[142];
assign function_psimd_s_mul32x32_acc64_func0 = dsp_function_ctrl[143];
assign function_psimd_s_mul32x32_acc64_func1 = dsp_function_ctrl[144];
assign function_psimd_s_mul32x32_acc64_func2 = dsp_function_ctrl[145];
assign function_psimd_s_mul32x32_acc64_func3 = dsp_function_ctrl[146];
assign function_psimd_s_mul32x32_acc64_func4 = dsp_function_ctrl[147];
assign function_psimd_s_mul32x32_acc64_func5 = dsp_function_ctrl[148];
assign function_psimd_s_mul32x32_acc64_func6 = dsp_function_ctrl[149];
assign function_psimd_s_pk32 = dsp_function_ctrl[150];
assign result_simd_s_wrap16 = dsp_result_ctrl[0];
assign result_simd_s_halve16 = dsp_result_ctrl[1];
assign result_simd_u_halve16 = dsp_result_ctrl[2];
assign result_simd_s_sat16 = dsp_result_ctrl[3];
assign result_simd_u_sat16 = dsp_result_ctrl[4];
assign result_simd_s_rnd16 = dsp_result_ctrl[6];
assign result_simd_s_rndsat16 = dsp_result_ctrl[7];
assign result_simd_s_wrap8 = dsp_result_ctrl[13];
assign result_simd_s_halve8 = dsp_result_ctrl[14];
assign result_simd_u_halve8 = dsp_result_ctrl[15];
assign result_simd_s_sat8 = dsp_result_ctrl[16];
assign result_simd_u_sat8 = dsp_result_ctrl[17];
assign result_simd_s_rnd8 = dsp_result_ctrl[19];
assign result_simd_s_rndsat8 = dsp_result_ctrl[20];
assign result_simd_s_unpk8 = dsp_result_ctrl[26];
assign result_psimd_s_halve32_sexlen = dsp_result_ctrl[28];
assign result_psimd_u_halve32_sexlen = dsp_result_ctrl[29];
assign result_psimd_s_rndxlen = dsp_result_ctrl[30];
assign result_psimd_s_sat32_sexlen = dsp_result_ctrl[31];
assign result_psimd_s_bypass32_sexlen = dsp_result_ctrl[35];
assign result_psimd_s_cmpsel32_sexlen = dsp_result_ctrl[38];
assign result_simd_s_bypass32 = dsp_result_ctrl[40];
assign result_simd_s_rnd32 = dsp_result_ctrl[41];
assign result_simd_s_sat32 = dsp_result_ctrl[42];
assign result_simd_s_rnd32_sat32 = dsp_result_ctrl[43];
assign result_psimd_s_sat32 = dsp_result_ctrl[45];
assign result_64p_s_wrap64 = dsp_result_ctrl[47];
assign result_64p_s_halve64 = dsp_result_ctrl[48];
assign result_64p_u_halve64 = dsp_result_ctrl[49];
assign result_64p_s_sat64 = dsp_result_ctrl[50];
assign result_64p_u_sat64 = dsp_result_ctrl[51];
assign result_nsimd_s_sat16_sexlen = dsp_result_ctrl[53];
assign result_nsimd_u_sat16_sexlen = dsp_result_ctrl[54];
assign result_nsimd_s_sat32_sexlen = dsp_result_ctrl[55];
assign result_nsimd_u_sat32_sexlen = dsp_result_ctrl[56];
assign result_nsimd_s_rndsat32_sexlen = dsp_result_ctrl[57];
assign result_nsimd_s_halvexlen = dsp_result_ctrl[58];
assign result_simd_s_wrap32 = dsp_result_ctrl[59];
assign result_simd_s_halve32 = dsp_result_ctrl[60];
assign result_simd_u_halve32 = dsp_result_ctrl[61];
assign result_simd_u_sat32 = dsp_result_ctrl[62];
assign result_simd_s_rndsat32 = dsp_result_ctrl[63];
assign result_nsimd_s_rnd32_se64 = dsp_result_ctrl[65];
assign result_psimd_s_sat64 = dsp_result_ctrl[66];
assign result_nsimd_s_sat16_se32 = dsp_result_ctrl[67];
assign result_nsimd_s_sat32 = dsp_result_ctrl[68];
assign dsp_src1_64b_sxlen = {{32{dsp_data_src1[31]}},dsp_data_src1};
assign dsp_src2_64b_sxlen = {{32{dsp_data_src2[31]}},dsp_data_src2};
assign dsp_src1_64b_simd = {32'd0,dsp_data_src1};
assign dsp_src2_64b_simd = {32'd0,dsp_data_src2};
assign dsp_src3_64b_simd = {32'd0,dsp_data_src3};
assign dsp_src1_64b_pair = {dsp_data_src3,dsp_data_src1};
assign dsp_src2_64b_pair = {dsp_data_src4,dsp_data_src2};
assign dsp_src3_64b_pair = {dsp_data_src4,dsp_data_src3};
assign dsp_src1_W1 = dsp_src1_64b_simd[63:32];
assign dsp_src1_W0 = dsp_src1_64b_simd[31:0];
assign dsp_src2_W1 = dsp_src2_64b_simd[63:32];
assign dsp_src2_W0 = dsp_src2_64b_simd[31:0];
assign dsp_src1_H3 = dsp_src1_64b_simd[63:48];
assign dsp_src1_H2 = dsp_src1_64b_simd[47:32];
assign dsp_src1_H1 = dsp_src1_64b_simd[31:16];
assign dsp_src1_H0 = dsp_src1_64b_simd[15:0];
assign dsp_src2_H3 = dsp_src2_64b_simd[63:48];
assign dsp_src2_H2 = dsp_src2_64b_simd[47:32];
assign dsp_src2_H1 = dsp_src2_64b_simd[31:16];
assign dsp_src2_H0 = dsp_src2_64b_simd[15:0];
assign dsp_src1_B7 = dsp_src1_64b_simd[63:56];
assign dsp_src1_B6 = dsp_src1_64b_simd[55:48];
assign dsp_src1_B5 = dsp_src1_64b_simd[47:40];
assign dsp_src1_B4 = dsp_src1_64b_simd[39:32];
assign dsp_src1_B3 = dsp_src1_64b_simd[31:24];
assign dsp_src1_B2 = dsp_src1_64b_simd[23:16];
assign dsp_src1_B1 = dsp_src1_64b_simd[15:8];
assign dsp_src1_B0 = dsp_src1_64b_simd[7:0];
assign dsp_src2_B7 = dsp_src2_64b_simd[63:56];
assign dsp_src2_B6 = dsp_src2_64b_simd[55:48];
assign dsp_src2_B5 = dsp_src2_64b_simd[47:40];
assign dsp_src2_B4 = dsp_src2_64b_simd[39:32];
assign dsp_src2_B3 = dsp_src2_64b_simd[31:24];
assign dsp_src2_B2 = dsp_src2_64b_simd[23:16];
assign dsp_src2_B1 = dsp_src2_64b_simd[15:8];
assign dsp_src2_B0 = dsp_src2_64b_simd[7:0];
assign dsp_src3_B7 = dsp_src3_64b_simd[63:56];
assign dsp_src3_B6 = dsp_src3_64b_simd[55:48];
assign dsp_src3_B5 = dsp_src3_64b_simd[47:40];
assign dsp_src3_B4 = dsp_src3_64b_simd[39:32];
assign dsp_src3_B3 = dsp_src3_64b_simd[31:24];
assign dsp_src3_B2 = dsp_src3_64b_simd[23:16];
assign dsp_src3_B1 = dsp_src3_64b_simd[15:8];
assign dsp_src3_B0 = dsp_src3_64b_simd[7:0];
assign dsp_clipmin_W = dsp_data_src3[31:0];
assign dsp_clipmin_H = dsp_data_src3[15:0];
assign dsp_clipmin_B = dsp_data_src3[7:0];
assign dsp_clipmax_W = dsp_data_src4[31:0];
assign dsp_clipmax_H = dsp_data_src4[15:0];
assign dsp_clipmax_B = dsp_data_src4[7:0];
assign simd16_op1_bottom16_sel = operand_simd_op16 | operand_simd_clip_op16 | operand_simd_cross_op16 | operand_psimd_op16 | operand_psimd_cross_op16 | operand_psimd_op16b_op16b | operand_psimd_op16b_op16t | operand_64p_op16 | operand_64p_cross_op16 | operand_64p_op16b_op16b | operand_64p_op16b_op16t | operand_nsimd_op16b_op16b | operand_nsimd_op16b_op16t;
assign simd16_op1_top16_sel = operand_psimd_op16t_op16t | operand_psimd_op16t_op16b | operand_psimd_reverse_op16 | operand_64p_op16t_op16t | operand_64p_reverse_op16 | operand_nsimd_op16t_op16t;
assign simd16_op1_smal_sel = operand_psimd_smal_op16;
assign simd16_op2_bottom16_sel = operand_simd_op16 | operand_psimd_op16 | operand_psimd_op16b_op16b | operand_psimd_op16t_op16b | operand_psimd_smal_op16 | operand_64p_op16 | operand_64p_op16b_op16b | operand_nsimd_op16b_op16b;
assign simd16_op2_top16_sel = operand_simd_cross_op16 | operand_psimd_cross_op16 | operand_psimd_op16b_op16t | operand_psimd_op16t_op16t | operand_psimd_reverse_op16 | operand_64p_cross_op16 | operand_64p_op16b_op16t | operand_64p_op16t_op16t | operand_64p_reverse_op16 | operand_nsimd_op16b_op16t | operand_nsimd_op16t_op16t;
assign simd16_op2_clipmin_sel_H0 = operand_simd_clip_op16 & dsp_src1_H0[15];
assign simd16_op2_clipmax_sel_H0 = operand_simd_clip_op16 & !dsp_src1_H0[15];
assign simd16_op2_clipmin_sel_H1 = operand_simd_clip_op16 & dsp_src1_H1[15];
assign simd16_op2_clipmax_sel_H1 = operand_simd_clip_op16 & !dsp_src1_H1[15];
assign simd16_op2_clipmin_sel_H2 = operand_simd_clip_op16 & dsp_src1_H2[15];
assign simd16_op2_clipmax_sel_H2 = operand_simd_clip_op16 & !dsp_src1_H2[15];
assign simd16_op2_clipmin_sel_H3 = operand_simd_clip_op16 & dsp_src1_H3[15];
assign simd16_op2_clipmax_sel_H3 = operand_simd_clip_op16 & !dsp_src1_H3[15];
assign simd16_op1_H0 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H0) | ({16{simd16_op1_top16_sel}} & dsp_src1_H1) | ({16{simd16_op1_smal_sel}} & dsp_src2_H1);
assign simd16_op2_H0 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H0) | ({16{simd16_op2_top16_sel}} & dsp_src2_H1) | ({16{simd16_op2_clipmin_sel_H0}} & dsp_clipmin_H) | ({16{simd16_op2_clipmax_sel_H0}} & dsp_clipmax_H);
assign simd16_op1_H1 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H1) | ({16{simd16_op1_top16_sel}} & dsp_src1_H0);
assign simd16_op2_H1 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H1) | ({16{simd16_op2_top16_sel}} & dsp_src2_H0) | ({16{simd16_op2_clipmin_sel_H1}} & dsp_clipmin_H) | ({16{simd16_op2_clipmax_sel_H1}} & dsp_clipmax_H);
assign simd16_op1_H2 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H2) | ({16{simd16_op1_top16_sel}} & dsp_src1_H3) | ({16{simd16_op1_smal_sel}} & dsp_src2_H3);
assign simd16_op2_H2 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H2) | ({16{simd16_op2_top16_sel}} & dsp_src2_H3) | ({16{simd16_op2_clipmin_sel_H2}} & dsp_clipmin_H) | ({16{simd16_op2_clipmax_sel_H2}} & dsp_clipmax_H);
assign simd16_op1_H3 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H3) | ({16{simd16_op1_top16_sel}} & dsp_src1_H2);
assign simd16_op2_H3 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H3) | ({16{simd16_op2_top16_sel}} & dsp_src2_H2) | ({16{simd16_op2_clipmin_sel_H3}} & dsp_clipmin_H) | ({16{simd16_op2_clipmax_sel_H3}} & dsp_clipmax_H);
assign simd16_mul_op1_H0 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H0) | ({16{simd16_op1_top16_sel}} & dsp_src1_H1) | ({16{simd16_op1_smal_sel}} & dsp_src2_H1);
assign simd16_mul_op2_H0 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H0) | ({16{simd16_op2_top16_sel}} & dsp_src2_H1);
assign simd16_mul_op1_H1 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H1) | ({16{simd16_op1_top16_sel}} & dsp_src1_H0);
assign simd16_mul_op2_H1 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H1) | ({16{simd16_op2_top16_sel}} & dsp_src2_H0);
assign simd16_mul_op1_H2 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H2) | ({16{simd16_op1_top16_sel}} & dsp_src1_H3) | ({16{simd16_op1_smal_sel}} & dsp_src2_H3);
assign simd16_mul_op2_H2 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H2) | ({16{simd16_op2_top16_sel}} & dsp_src2_H3);
assign simd16_mul_op1_H3 = ({16{simd16_op1_bottom16_sel}} & dsp_src1_H3) | ({16{simd16_op1_top16_sel}} & dsp_src1_H2);
assign simd16_mul_op2_H3 = ({16{simd16_op2_bottom16_sel}} & dsp_src2_H3) | ({16{simd16_op2_top16_sel}} & dsp_src2_H2);
function  [17:0] simd16_addcmp_func;
input se1;
input se2;
input neg1;
input neg2;
input [15:0] op1;
input [15:0] op2;
reg [16:0] adder_in1;
reg [16:0] adder_in2;
reg adder_cin;
reg [16:0] adder_out;
reg cmpeq_out;
begin
    adder_in1 = {17{neg1}} ^ {(se1 & op1[15]),op1};
    adder_in2 = {17{neg2}} ^ {(se2 & op2[15]),op2};
    adder_cin = neg1 | neg2;
    adder_out = adder_in1 + adder_in2 + {16'd0,adder_cin};
    cmpeq_out = (op1 == op2);
    simd16_addcmp_func = {cmpeq_out,adder_out};
end
endfunction
function  [16:0] simd16_addcmp_result;
input is_func_sub;
input is_func_cmpeq;
input is_func_cmplt;
input is_func_cmple;
input is_func_min;
input is_func_max;
input is_func_clip;
input is_type_wrap;
input is_type_halve;
input is_type_s_sat;
input is_type_u_sat;
input [15:0] cmp_op1;
input [15:0] cmp_op2;
input [17:0] din;
reg [15:0] dout;
reg ovfout;
reg is_eq;
reg is_lt;
reg is_le;
reg is_gt;
reg exceed_clip_bound;
reg wrap_sel;
reg halve_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg u_ovf_sel;
reg u_udf_sel;
reg cmp_op1_sel;
reg cmp_op2_sel;
reg cmp_t_sel;
begin
    is_eq = din[17];
    is_lt = din[16];
    is_le = is_eq | is_lt;
    is_gt = !is_le;
    exceed_clip_bound = is_func_clip & ((!cmp_op1[15] & is_gt) | (cmp_op1[15] & is_lt));
    halve_sel = is_type_halve;
    s_ovf_sel = is_type_s_sat & (din[16:15] == 2'b01);
    s_udf_sel = is_type_s_sat & (din[16:15] == 2'b10);
    u_ovf_sel = is_type_u_sat & din[16] & !is_func_sub;
    u_udf_sel = is_type_u_sat & din[16] & is_func_sub;
    wrap_sel = is_type_wrap | (is_type_s_sat & !(s_ovf_sel | s_udf_sel)) | (is_type_u_sat & !(u_ovf_sel | u_udf_sel));
    cmp_t_sel = (is_func_cmpeq & is_eq) | (is_func_cmplt & is_lt) | (is_func_cmple & is_le);
    cmp_op1_sel = (is_func_min & din[16]) | (is_func_max & !din[16]) | (is_func_clip & !exceed_clip_bound);
    cmp_op2_sel = (is_func_min & !din[16]) | (is_func_max & din[16]) | (is_func_clip & exceed_clip_bound);
    dout = ({16{wrap_sel}} & din[15:0]) | ({16{halve_sel}} & din[16:1]) | ({16{s_ovf_sel}} & 16'h7fff) | ({16{s_udf_sel}} & 16'h8000) | ({16{u_ovf_sel}} & 16'hffff) | ({16{u_udf_sel}} & 16'h0000) | ({16{cmp_t_sel}} & 16'hffff) | ({16{cmp_op1_sel}} & cmp_op1) | ({16{cmp_op2_sel}} & cmp_op2);
    ovfout = s_ovf_sel | s_udf_sel | u_ovf_sel | u_udf_sel | exceed_clip_bound;
    simd16_addcmp_result = {ovfout,dout};
end
endfunction
assign simd16_addcmp_se1_H0 = function_simd_s_add16 | function_simd_s_sub16 | function_simd_s_as16 | function_simd_s_sa16 | function_simd_s_cmplt16 | function_simd_s_cmple16 | function_simd_s_min16 | function_simd_s_max16 | function_simd_s_abs16 | function_simd_s_clip16;
assign simd16_addcmp_se1_H1 = simd16_addcmp_se1_H0;
assign simd16_addcmp_se1_H2 = simd16_addcmp_se1_H0;
assign simd16_addcmp_se1_H3 = simd16_addcmp_se1_H0;
assign simd16_addcmp_se2_H0 = function_simd_s_add16 | function_simd_s_sub16 | function_simd_s_as16 | function_simd_s_sa16 | function_simd_s_cmplt16 | function_simd_s_cmple16 | function_simd_s_min16 | function_simd_s_max16 | function_simd_s_abs16 | function_simd_s_clip16;
assign simd16_addcmp_se2_H1 = simd16_addcmp_se2_H0;
assign simd16_addcmp_se2_H2 = simd16_addcmp_se2_H0;
assign simd16_addcmp_se2_H3 = simd16_addcmp_se2_H0;
assign simd16_addcmp_neg1_H0 = (function_simd_s_abs16 & simd16_op1_H0[15]);
assign simd16_addcmp_neg1_H1 = (function_simd_s_abs16 & simd16_op1_H1[15]);
assign simd16_addcmp_neg1_H2 = (function_simd_s_abs16 & simd16_op1_H2[15]);
assign simd16_addcmp_neg1_H3 = (function_simd_s_abs16 & simd16_op1_H3[15]);
assign simd16_addcmp_neg2_H0 = function_simd_s_sub16 | function_simd_u_sub16 | function_simd_s_as16 | function_simd_u_as16 | function_simd_s_cmplt16 | function_simd_u_cmplt16 | function_simd_s_cmple16 | function_simd_u_cmple16 | function_simd_s_min16 | function_simd_u_min16 | function_simd_s_max16 | function_simd_u_max16 | function_simd_s_clip16;
assign simd16_addcmp_neg2_H1 = function_simd_s_sub16 | function_simd_u_sub16 | function_simd_s_sa16 | function_simd_u_sa16 | function_simd_s_cmplt16 | function_simd_u_cmplt16 | function_simd_s_cmple16 | function_simd_u_cmple16 | function_simd_s_min16 | function_simd_u_min16 | function_simd_s_max16 | function_simd_u_max16 | function_simd_s_clip16;
assign simd16_addcmp_neg2_H2 = simd16_addcmp_neg2_H0;
assign simd16_addcmp_neg2_H3 = simd16_addcmp_neg2_H1;
assign simd16_addcmp_out_H0 = simd16_addcmp_func(simd16_addcmp_se1_H0, simd16_addcmp_se2_H0, simd16_addcmp_neg1_H0, simd16_addcmp_neg2_H0, simd16_op1_H0, simd16_op2_H0);
assign simd16_addcmp_out_H1 = simd16_addcmp_func(simd16_addcmp_se1_H1, simd16_addcmp_se2_H1, simd16_addcmp_neg1_H1, simd16_addcmp_neg2_H1, simd16_op1_H1, simd16_op2_H1);
assign simd16_addcmp_out_H2 = simd16_addcmp_func(simd16_addcmp_se1_H2, simd16_addcmp_se2_H2, simd16_addcmp_neg1_H2, simd16_addcmp_neg2_H2, simd16_op1_H2, simd16_op2_H2);
assign simd16_addcmp_out_H3 = simd16_addcmp_func(simd16_addcmp_se1_H3, simd16_addcmp_se2_H3, simd16_addcmp_neg1_H3, simd16_addcmp_neg2_H3, simd16_op1_H3, simd16_op2_H3);
assign simd16_addcmp_wrap = result_simd_s_wrap16;
assign simd16_addcmp_halve = result_simd_s_halve16 | result_simd_u_halve16;
assign simd16_addcmp_s_sat = result_simd_s_sat16;
assign simd16_addcmp_u_sat = result_simd_u_sat16;
assign simd16_addcmp_result_H0 = simd16_addcmp_result(simd16_addcmp_neg2_H0, function_simd_s_cmpeq16, (function_simd_s_cmplt16 | function_simd_u_cmplt16), (function_simd_s_cmple16 | function_simd_u_cmple16), (function_simd_s_min16 | function_simd_u_min16), (function_simd_s_max16 | function_simd_u_max16), function_simd_s_clip16, simd16_addcmp_wrap, simd16_addcmp_halve, simd16_addcmp_s_sat, simd16_addcmp_u_sat, simd16_op1_H0, simd16_op2_H0, simd16_addcmp_out_H0);
assign simd16_addcmp_result_H1 = simd16_addcmp_result(simd16_addcmp_neg2_H1, function_simd_s_cmpeq16, (function_simd_s_cmplt16 | function_simd_u_cmplt16), (function_simd_s_cmple16 | function_simd_u_cmple16), (function_simd_s_min16 | function_simd_u_min16), (function_simd_s_max16 | function_simd_u_max16), function_simd_s_clip16, simd16_addcmp_wrap, simd16_addcmp_halve, simd16_addcmp_s_sat, simd16_addcmp_u_sat, simd16_op1_H1, simd16_op2_H1, simd16_addcmp_out_H1);
assign simd16_addcmp_result_H2 = simd16_addcmp_result(simd16_addcmp_neg2_H2, function_simd_s_cmpeq16, (function_simd_s_cmplt16 | function_simd_u_cmplt16), (function_simd_s_cmple16 | function_simd_u_cmple16), (function_simd_s_min16 | function_simd_u_min16), (function_simd_s_max16 | function_simd_u_max16), function_simd_s_clip16, simd16_addcmp_wrap, simd16_addcmp_halve, simd16_addcmp_s_sat, simd16_addcmp_u_sat, simd16_op1_H2, simd16_op2_H2, simd16_addcmp_out_H2);
assign simd16_addcmp_result_H3 = simd16_addcmp_result(simd16_addcmp_neg2_H3, function_simd_s_cmpeq16, (function_simd_s_cmplt16 | function_simd_u_cmplt16), (function_simd_s_cmple16 | function_simd_u_cmple16), (function_simd_s_min16 | function_simd_u_min16), (function_simd_s_max16 | function_simd_u_max16), function_simd_s_clip16, simd16_addcmp_wrap, simd16_addcmp_halve, simd16_addcmp_s_sat, simd16_addcmp_u_sat, simd16_op1_H3, simd16_op2_H3, simd16_addcmp_out_H3);
assign simd16_addcmp_result_64b = {simd16_addcmp_result_H3[15:0],simd16_addcmp_result_H2[15:0],simd16_addcmp_result_H1[15:0],simd16_addcmp_result_H0[15:0]};
assign simd16_addcmp_ovf_set = simd16_addcmp_result_H0[16] | simd16_addcmp_result_H1[16] | simd16_addcmp_result_H2[16] | simd16_addcmp_result_H3[16];
function  [16:0] simd16_shift;
integer i;
input is_func_slra;
input is_func_sll;
input rnd;
input sat;
input se;
input [15:0] op1;
input [4:0] amt;
reg is_pos_amt;
reg is_neg_amt;
reg is_ovf_amt;
reg is_shift_l;
reg [3:0] shift_amt;
reg [31:0] shift_l_din;
reg [31:0] shift_r_din;
reg [31:0] shift_din;
reg signed [31:0] shift_r_dout;
reg [31:0] shift_l_dout;
reg [31:0] shift_dout;
reg is_type_s_rnd;
reg is_type_s_sat;
reg s_rnd_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg [16:0] rnd_dout;
reg [15:0] result;
reg ovfout;
begin
    is_pos_amt = is_func_slra & !amt[4];
    is_neg_amt = is_func_slra & amt[4];
    is_ovf_amt = is_func_slra & (amt[4:0] == 5'd16);
    is_shift_l = is_func_sll | is_pos_amt;
    shift_amt = is_ovf_amt ? 4'd15 : is_neg_amt ? (~amt[3:0] + 4'd1) : amt[3:0];
    shift_r_din = {{15{(se & op1[15])}},op1,1'b0};
    for (i = 0; i < 32; i = i + 1) begin:gen_shift_l_din
        shift_l_din[i] = shift_r_din[31 - i];
    end
    shift_din = is_shift_l ? shift_l_din : shift_r_din;
    shift_r_dout = $signed(shift_din) >>> shift_amt;
    for (i = 0; i < 32; i = i + 1) begin:gen_shift_l_dout
        shift_l_dout[i] = shift_r_dout[31 - i];
    end
    shift_dout = is_shift_l ? shift_l_dout : shift_r_dout;
    is_type_s_rnd = is_func_slra ? (rnd & is_neg_amt) : rnd;
    is_type_s_sat = is_func_slra ? (sat & is_pos_amt) : sat;
    s_ovf_sel = is_type_s_sat & !shift_dout[31] & (shift_dout[30:16] != 15'h0000);
    s_udf_sel = is_type_s_sat & shift_dout[31] & (shift_dout[30:16] != 15'h7fff);
    s_rnd_sel = !(s_ovf_sel | s_udf_sel);
    rnd_dout = shift_dout[16:0] + {16'd0,is_type_s_rnd};
    result = ({16{s_rnd_sel}} & rnd_dout[16:1]) | ({16{s_ovf_sel}} & 16'h7fff) | ({16{s_udf_sel}} & 16'h8000);
    ovfout = s_ovf_sel | s_udf_sel;
    simd16_shift = {ovfout,result};
end
endfunction
assign simd16_shift_result_H0 = simd16_shift(function_simd_s_slra16, function_simd_s_sll16, (result_simd_s_rnd16 | result_simd_s_rndsat16), (result_simd_s_sat16 | result_simd_s_rndsat16), !function_simd_u_srl16, simd16_op1_H0, dsp_data_src2[4:0]);
assign simd16_shift_result_H1 = simd16_shift(function_simd_s_slra16, function_simd_s_sll16, (result_simd_s_rnd16 | result_simd_s_rndsat16), (result_simd_s_sat16 | result_simd_s_rndsat16), !function_simd_u_srl16, simd16_op1_H1, dsp_data_src2[4:0]);
assign simd16_shift_result_H2 = simd16_shift(function_simd_s_slra16, function_simd_s_sll16, (result_simd_s_rnd16 | result_simd_s_rndsat16), (result_simd_s_sat16 | result_simd_s_rndsat16), !function_simd_u_srl16, simd16_op1_H2, dsp_data_src2[4:0]);
assign simd16_shift_result_H3 = simd16_shift(function_simd_s_slra16, function_simd_s_sll16, (result_simd_s_rnd16 | result_simd_s_rndsat16), (result_simd_s_sat16 | result_simd_s_rndsat16), !function_simd_u_srl16, simd16_op1_H3, dsp_data_src2[4:0]);
assign simd16_shift_result_64b = {simd16_shift_result_H3[15:0],simd16_shift_result_H2[15:0],simd16_shift_result_H1[15:0],simd16_shift_result_H0[15:0]};
assign simd16_shift_ovf_set = simd16_shift_result_H0[16] | simd16_shift_result_H1[16] | simd16_shift_result_H2[16] | simd16_shift_result_H3[16];
function  [31:0] simd16_mul_func;
input se1;
input se2;
input [15:0] op1;
input [15:0] op2;
reg [33:0] mul_in1;
reg [33:0] mul_in2;
reg signed [33:0] mul_out;
begin
    mul_in1 = {{18{(se1 & op1[15])}},op1};
    mul_in2 = {{18{(se2 & op2[15])}},op2};
    mul_out = $signed(mul_in1) * $signed(mul_in2);
    simd16_mul_func = mul_out[31:0];
end
endfunction
function  [16:0] simd16_mul_result;
input is_type_s_sat;
input [15:0] op1;
input [15:0] op2;
input [31:0] din;
reg [15:0] dout;
reg ovfout;
reg s_ovf_sel;
reg sra15_sel;
begin
    s_ovf_sel = is_type_s_sat & (op1 == 16'h8000) & (op2 == 16'h8000);
    sra15_sel = !s_ovf_sel;
    dout = ({16{sra15_sel}} & din[30:15]) | ({16{s_ovf_sel}} & 16'h7fff);
    ovfout = s_ovf_sel;
    simd16_mul_result = {ovfout,dout};
end
endfunction
assign simd16_mul_se1_H0 = function_simd_s_mul16 | function_psimd_s_mul16x16_acc32_func0 | function_psimd_s_mul16x16_acc32_func1 | function_psimd_s_mul16x16_acc32_func2 | function_psimd_s_mul16x16_acc32_func3 | function_psimd_s_mul16x16_acc32_func4 | function_psimd_s_mul16x16_acc32_func5 | function_psimd_s_mul16x16_acc32_func6 | function_psimd_s_mul16x16_acc64_func0 | function_psimd_s_mul16x16_out64 | function_64p_s_mul16x16_acc64_func0 | function_64p_s_mul16x16_acc64_func1 | function_64p_s_mul16x16_acc64_func2 | function_64p_s_mul16x16_acc64_func3 | function_nsimd_s_mul16x16 | function_nsimd_s_mul16x16_double32 | function_nsimd_s_mul16x16_double32_acc32;
assign simd16_mul_se1_H1 = simd16_mul_se1_H0;
assign simd16_mul_se1_H2 = simd16_mul_se1_H0;
assign simd16_mul_se1_H3 = simd16_mul_se1_H0;
assign simd16_mul_se2_H0 = function_simd_s_mul16 | function_psimd_s_mul16x16_acc32_func0 | function_psimd_s_mul16x16_acc32_func1 | function_psimd_s_mul16x16_acc32_func2 | function_psimd_s_mul16x16_acc32_func3 | function_psimd_s_mul16x16_acc32_func4 | function_psimd_s_mul16x16_acc32_func5 | function_psimd_s_mul16x16_acc32_func6 | function_psimd_s_mul16x16_acc64_func0 | function_psimd_s_mul16x16_out64 | function_64p_s_mul16x16_acc64_func0 | function_64p_s_mul16x16_acc64_func1 | function_64p_s_mul16x16_acc64_func2 | function_64p_s_mul16x16_acc64_func3 | function_nsimd_s_mul16x16 | function_nsimd_s_mul16x16_double32 | function_nsimd_s_mul16x16_double32_acc32;
assign simd16_mul_se2_H1 = simd16_mul_se2_H0;
assign simd16_mul_se2_H2 = simd16_mul_se2_H0;
assign simd16_mul_se2_H3 = simd16_mul_se2_H0;
assign simd16_mul_out_H0 = simd16_mul_func(simd16_mul_se1_H0, simd16_mul_se2_H0, simd16_op1_H0, simd16_op2_H0);
assign simd16_mul_out_H1 = simd16_mul_func(simd16_mul_se1_H1, simd16_mul_se2_H1, simd16_op1_H1, simd16_op2_H1);
assign simd16_mul_out_H2 = simd16_mul_func(simd16_mul_se1_H2, simd16_mul_se2_H2, simd16_op1_H2, simd16_op2_H2);
assign simd16_mul_out_H3 = simd16_mul_func(simd16_mul_se1_H3, simd16_mul_se2_H3, simd16_op1_H3, simd16_op2_H3);
assign simd16_mul_s_sat = result_simd_s_sat16;
assign simd16_mul_result_H0 = simd16_mul_result(simd16_mul_s_sat, simd16_mul_op1_H0, simd16_mul_op2_H0, simd16_mul_out_H0);
assign simd16_mul_result_H1 = simd16_mul_result(simd16_mul_s_sat, simd16_mul_op1_H1, simd16_mul_op2_H1, simd16_mul_out_H1);
assign simd16_mul_result_H2 = simd16_mul_result(simd16_mul_s_sat, simd16_mul_op1_H2, simd16_mul_op2_H2, simd16_mul_out_H2);
assign simd16_mul_result_H3 = simd16_mul_result(simd16_mul_s_sat, simd16_mul_op1_H3, simd16_mul_op2_H3, simd16_mul_out_H3);
assign simd16_mul_result_64b = {simd16_mul_result_H3[15:0],simd16_mul_result_H2[15:0],simd16_mul_result_H1[15:0],simd16_mul_result_H0[15:0]};
assign simd16_mul_ovf_set = simd16_mul_result_H0[16] | simd16_mul_result_H1[16] | simd16_mul_result_H2[16] | simd16_mul_result_H3[16];
assign simd16_swap_result_64b = {simd16_op1_H2[15:0],simd16_op1_H3[15:0],simd16_op1_H0[15:0],simd16_op1_H1[15:0]};
assign simd16_swap_ovf_set = 1'b0;
function  [15:0] simd16_clz;
input is_func_clz;
input is_func_clo;
input is_func_clrs;
input [15:0] op1;
reg [15:0] clz_in_16b;
reg [7:0] clz_in_8b;
reg [3:0] clz_in_4b;
reg [3:0] clz_out;
reg clz_in_eqz;
begin
    clz_in_16b = ({16{is_func_clz}} & op1) | ({16{is_func_clo}} & ~op1) | ({16{is_func_clrs}} & ({op1[14:0],!op1[15]} ^ {16{op1[15]}}));
    clz_out[3] = (clz_in_16b[15:8] == 8'd0);
    clz_in_8b = clz_out[3] ? clz_in_16b[7:0] : clz_in_16b[15:8];
    clz_out[2] = (clz_in_8b[7:4] == 4'd0);
    clz_in_4b = clz_out[2] ? clz_in_8b[3:0] : clz_in_8b[7:4];
    clz_out[1] = (clz_in_4b[3:2] == 2'd0);
    clz_out[0] = clz_out[1] ? !clz_in_4b[1] : !clz_in_4b[3];
    clz_in_eqz = (clz_in_16b == 16'd0);
    simd16_clz = clz_in_eqz ? 16'd16 : {12'd0,clz_out[3:0]};
end
endfunction
assign simd16_clz_result_H0 = simd16_clz(function_simd_s_clz16, function_simd_s_clo16, function_simd_s_clrs16, simd16_op1_H0);
assign simd16_clz_result_H1 = simd16_clz(function_simd_s_clz16, function_simd_s_clo16, function_simd_s_clrs16, simd16_op1_H1);
assign simd16_clz_result_H2 = simd16_clz(function_simd_s_clz16, function_simd_s_clo16, function_simd_s_clrs16, simd16_op1_H2);
assign simd16_clz_result_H3 = simd16_clz(function_simd_s_clz16, function_simd_s_clo16, function_simd_s_clrs16, simd16_op1_H3);
assign simd16_clz_result_64b = {simd16_clz_result_H3[15:0],simd16_clz_result_H2[15:0],simd16_clz_result_H1[15:0],simd16_clz_result_H0[15:0]};
assign simd16_clz_ovf_set = 1'b0;
assign simd16_result_addcmp_sel = function_simd_s_add16 | function_simd_u_add16 | function_simd_s_sub16 | function_simd_u_sub16 | function_simd_s_as16 | function_simd_u_as16 | function_simd_s_sa16 | function_simd_u_sa16 | function_simd_s_cmpeq16 | function_simd_s_cmplt16 | function_simd_u_cmplt16 | function_simd_s_cmple16 | function_simd_u_cmple16 | function_simd_s_min16 | function_simd_u_min16 | function_simd_s_max16 | function_simd_u_max16 | function_simd_s_abs16 | function_simd_s_clip16;
assign simd16_result_shift_sel = function_simd_s_sra16 | function_simd_u_srl16 | function_simd_s_sll16 | function_simd_s_slra16;
assign simd16_result_mul_sel = function_simd_s_mul16;
assign simd16_result_swap_sel = function_simd_s_swap16;
assign simd16_result_clz_sel = function_simd_s_clz16 | function_simd_s_clo16 | function_simd_s_clrs16;
assign stage1_simd16_final_result_64b = ({64{simd16_result_addcmp_sel}} & simd16_addcmp_result_64b) | ({64{simd16_result_shift_sel}} & simd16_shift_result_64b) | ({64{simd16_result_swap_sel}} & simd16_swap_result_64b) | ({64{simd16_result_clz_sel}} & simd16_clz_result_64b);
assign stage1_simd16_final_ovf_set = (simd16_result_addcmp_sel & simd16_addcmp_ovf_set) | (simd16_result_shift_sel & simd16_shift_ovf_set) | (simd16_result_swap_sel & simd16_swap_ovf_set) | (simd16_result_clz_sel & simd16_clz_ovf_set);
assign simd8_op1_base_sel = operand_simd_op8 | operand_simd_clip_op8 | operand_simd_cross_op8 | operand_psimd_op8 | operand_psimd_cross_op8;
assign simd8_op2_base_sel = operand_simd_op8 | operand_psimd_op8;
assign simd8_op2_cross_sel = operand_simd_cross_op8 | operand_psimd_cross_op8;
assign simd8_op2_clipmin_sel_B0 = operand_simd_clip_op8 & dsp_src1_B0[7];
assign simd8_op2_clipmax_sel_B0 = operand_simd_clip_op8 & !dsp_src1_B0[7];
assign simd8_op2_clipmin_sel_B1 = operand_simd_clip_op8 & dsp_src1_B1[7];
assign simd8_op2_clipmax_sel_B1 = operand_simd_clip_op8 & !dsp_src1_B1[7];
assign simd8_op2_clipmin_sel_B2 = operand_simd_clip_op8 & dsp_src1_B2[7];
assign simd8_op2_clipmax_sel_B2 = operand_simd_clip_op8 & !dsp_src1_B2[7];
assign simd8_op2_clipmin_sel_B3 = operand_simd_clip_op8 & dsp_src1_B3[7];
assign simd8_op2_clipmax_sel_B3 = operand_simd_clip_op8 & !dsp_src1_B3[7];
assign simd8_op2_clipmin_sel_B4 = operand_simd_clip_op8 & dsp_src1_B4[7];
assign simd8_op2_clipmax_sel_B4 = operand_simd_clip_op8 & !dsp_src1_B4[7];
assign simd8_op2_clipmin_sel_B5 = operand_simd_clip_op8 & dsp_src1_B5[7];
assign simd8_op2_clipmax_sel_B5 = operand_simd_clip_op8 & !dsp_src1_B5[7];
assign simd8_op2_clipmin_sel_B6 = operand_simd_clip_op8 & dsp_src1_B6[7];
assign simd8_op2_clipmax_sel_B6 = operand_simd_clip_op8 & !dsp_src1_B6[7];
assign simd8_op2_clipmin_sel_B7 = operand_simd_clip_op8 & dsp_src1_B7[7];
assign simd8_op2_clipmax_sel_B7 = operand_simd_clip_op8 & !dsp_src1_B7[7];
assign simd8_op1_B0 = ({8{simd8_op1_base_sel}} & dsp_src1_B0);
assign simd8_op2_B0 = ({8{simd8_op2_base_sel}} & dsp_src2_B0) | ({8{simd8_op2_cross_sel}} & dsp_src2_B1) | ({8{simd8_op2_clipmin_sel_B0}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B0}} & dsp_clipmax_B);
assign simd8_op1_B1 = ({8{simd8_op1_base_sel}} & dsp_src1_B1);
assign simd8_op2_B1 = ({8{simd8_op2_base_sel}} & dsp_src2_B1) | ({8{simd8_op2_cross_sel}} & dsp_src2_B0) | ({8{simd8_op2_clipmin_sel_B1}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B1}} & dsp_clipmax_B);
assign simd8_op1_B2 = ({8{simd8_op1_base_sel}} & dsp_src1_B2);
assign simd8_op2_B2 = ({8{simd8_op2_base_sel}} & dsp_src2_B2) | ({8{simd8_op2_cross_sel}} & dsp_src2_B3) | ({8{simd8_op2_clipmin_sel_B2}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B2}} & dsp_clipmax_B);
assign simd8_op1_B3 = ({8{simd8_op1_base_sel}} & dsp_src1_B3);
assign simd8_op2_B3 = ({8{simd8_op2_base_sel}} & dsp_src2_B3) | ({8{simd8_op2_cross_sel}} & dsp_src2_B2) | ({8{simd8_op2_clipmin_sel_B3}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B3}} & dsp_clipmax_B);
assign simd8_op1_B4 = ({8{simd8_op1_base_sel}} & dsp_src1_B4);
assign simd8_op2_B4 = ({8{simd8_op2_base_sel}} & dsp_src2_B4) | ({8{simd8_op2_cross_sel}} & dsp_src2_B5) | ({8{simd8_op2_clipmin_sel_B4}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B4}} & dsp_clipmax_B);
assign simd8_op1_B5 = ({8{simd8_op1_base_sel}} & dsp_src1_B5);
assign simd8_op2_B5 = ({8{simd8_op2_base_sel}} & dsp_src2_B5) | ({8{simd8_op2_cross_sel}} & dsp_src2_B4) | ({8{simd8_op2_clipmin_sel_B5}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B5}} & dsp_clipmax_B);
assign simd8_op1_B6 = ({8{simd8_op1_base_sel}} & dsp_src1_B6);
assign simd8_op2_B6 = ({8{simd8_op2_base_sel}} & dsp_src2_B6) | ({8{simd8_op2_cross_sel}} & dsp_src2_B7) | ({8{simd8_op2_clipmin_sel_B6}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B6}} & dsp_clipmax_B);
assign simd8_op1_B7 = ({8{simd8_op1_base_sel}} & dsp_src1_B7);
assign simd8_op2_B7 = ({8{simd8_op2_base_sel}} & dsp_src2_B7) | ({8{simd8_op2_cross_sel}} & dsp_src2_B6) | ({8{simd8_op2_clipmin_sel_B7}} & dsp_clipmin_B) | ({8{simd8_op2_clipmax_sel_B7}} & dsp_clipmax_B);
function  [9:0] simd8_addcmp_func;
input se1;
input se2;
input neg1;
input neg2;
input [7:0] op1;
input [7:0] op2;
reg [8:0] adder_in1;
reg [8:0] adder_in2;
reg adder_cin;
reg [8:0] adder_out;
reg cmpeq_out;
begin
    adder_in1 = {9{neg1}} ^ {(se1 & op1[7]),op1};
    adder_in2 = {9{neg2}} ^ {(se2 & op2[7]),op2};
    adder_cin = neg1 | neg2;
    adder_out = adder_in1 + adder_in2 + {8'd0,adder_cin};
    cmpeq_out = (op1 == op2);
    simd8_addcmp_func = {cmpeq_out,adder_out};
end
endfunction
function  [8:0] simd8_addcmp_result;
input is_func_sub;
input is_func_cmpeq;
input is_func_cmplt;
input is_func_cmple;
input is_func_min;
input is_func_max;
input is_func_clip;
input is_type_wrap;
input is_type_halve;
input is_type_s_sat;
input is_type_u_sat;
input [7:0] cmp_op1;
input [7:0] cmp_op2;
input [9:0] din;
reg [7:0] dout;
reg ovfout;
reg is_eq;
reg is_lt;
reg is_le;
reg is_gt;
reg exceed_clip_bound;
reg wrap_sel;
reg halve_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg u_ovf_sel;
reg u_udf_sel;
reg cmp_op1_sel;
reg cmp_op2_sel;
reg cmp_t_sel;
begin
    is_eq = din[9];
    is_lt = din[8];
    is_le = is_eq | is_lt;
    is_gt = !is_le;
    exceed_clip_bound = is_func_clip & ((!cmp_op1[7] & is_gt) | (cmp_op1[7] & is_lt));
    halve_sel = is_type_halve;
    s_ovf_sel = is_type_s_sat & (din[8:7] == 2'b01);
    s_udf_sel = is_type_s_sat & (din[8:7] == 2'b10);
    u_ovf_sel = is_type_u_sat & din[8] & !is_func_sub;
    u_udf_sel = is_type_u_sat & din[8] & is_func_sub;
    wrap_sel = is_type_wrap | (is_type_s_sat & !(s_ovf_sel | s_udf_sel)) | (is_type_u_sat & !(u_ovf_sel | u_udf_sel));
    cmp_t_sel = (is_func_cmpeq & is_eq) | (is_func_cmplt & is_lt) | (is_func_cmple & is_le);
    cmp_op1_sel = (is_func_min & din[8]) | (is_func_max & !din[8]) | (is_func_clip & !exceed_clip_bound);
    cmp_op2_sel = (is_func_min & !din[8]) | (is_func_max & din[8]) | (is_func_clip & exceed_clip_bound);
    dout = ({8{wrap_sel}} & din[7:0]) | ({8{halve_sel}} & din[8:1]) | ({8{s_ovf_sel}} & 8'h7f) | ({8{s_udf_sel}} & 8'h80) | ({8{u_ovf_sel}} & 8'hff) | ({8{u_udf_sel}} & 8'h00) | ({8{cmp_t_sel}} & 8'hff) | ({8{cmp_op1_sel}} & cmp_op1) | ({8{cmp_op2_sel}} & cmp_op2);
    ovfout = s_ovf_sel | s_udf_sel | u_ovf_sel | u_udf_sel | exceed_clip_bound;
    simd8_addcmp_result = {ovfout,dout};
end
endfunction
assign simd8_addcmp_se1_B0 = function_simd_s_add8 | function_simd_s_sub8 | function_simd_s_cmplt8 | function_simd_s_cmple8 | function_simd_s_min8 | function_simd_s_max8 | function_simd_s_abs8 | function_simd_s_clip8;
assign simd8_addcmp_se1_B1 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B2 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B3 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B4 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B5 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B6 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se1_B7 = simd8_addcmp_se1_B0;
assign simd8_addcmp_se2_B0 = function_simd_s_add8 | function_simd_s_sub8 | function_simd_s_cmplt8 | function_simd_s_cmple8 | function_simd_s_min8 | function_simd_s_max8 | function_simd_s_abs8 | function_simd_s_clip8;
assign simd8_addcmp_se2_B1 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B2 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B3 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B4 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B5 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B6 = simd8_addcmp_se2_B0;
assign simd8_addcmp_se2_B7 = simd8_addcmp_se2_B0;
assign simd8_addcmp_neg1_B0 = (function_simd_s_abs8 & simd8_op1_B0[7]);
assign simd8_addcmp_neg1_B1 = (function_simd_s_abs8 & simd8_op1_B1[7]);
assign simd8_addcmp_neg1_B2 = (function_simd_s_abs8 & simd8_op1_B2[7]);
assign simd8_addcmp_neg1_B3 = (function_simd_s_abs8 & simd8_op1_B3[7]);
assign simd8_addcmp_neg1_B4 = (function_simd_s_abs8 & simd8_op1_B4[7]);
assign simd8_addcmp_neg1_B5 = (function_simd_s_abs8 & simd8_op1_B5[7]);
assign simd8_addcmp_neg1_B6 = (function_simd_s_abs8 & simd8_op1_B6[7]);
assign simd8_addcmp_neg1_B7 = (function_simd_s_abs8 & simd8_op1_B7[7]);
assign simd8_addcmp_neg2_B0 = function_simd_s_sub8 | function_simd_u_sub8 | function_simd_s_cmplt8 | function_simd_u_cmplt8 | function_simd_s_cmple8 | function_simd_u_cmple8 | function_simd_s_min8 | function_simd_u_min8 | function_simd_s_max8 | function_simd_u_max8 | function_simd_s_clip8 | function_psimd_u_abs8_accxlen_func0 | function_psimd_u_abs8_accxlen_func1;
assign simd8_addcmp_neg2_B1 = function_simd_s_sub8 | function_simd_u_sub8 | function_simd_s_cmplt8 | function_simd_u_cmplt8 | function_simd_s_cmple8 | function_simd_u_cmple8 | function_simd_s_min8 | function_simd_u_min8 | function_simd_s_max8 | function_simd_u_max8 | function_simd_s_clip8 | function_psimd_u_abs8_accxlen_func0 | function_psimd_u_abs8_accxlen_func1;
assign simd8_addcmp_neg2_B2 = simd8_addcmp_neg2_B0;
assign simd8_addcmp_neg2_B3 = simd8_addcmp_neg2_B1;
assign simd8_addcmp_neg2_B4 = simd8_addcmp_neg2_B0;
assign simd8_addcmp_neg2_B5 = simd8_addcmp_neg2_B1;
assign simd8_addcmp_neg2_B6 = simd8_addcmp_neg2_B0;
assign simd8_addcmp_neg2_B7 = simd8_addcmp_neg2_B1;
assign simd8_addcmp_out_B0 = simd8_addcmp_func(simd8_addcmp_se1_B0, simd8_addcmp_se2_B0, simd8_addcmp_neg1_B0, simd8_addcmp_neg2_B0, simd8_op1_B0, simd8_op2_B0);
assign simd8_addcmp_out_B1 = simd8_addcmp_func(simd8_addcmp_se1_B1, simd8_addcmp_se2_B1, simd8_addcmp_neg1_B1, simd8_addcmp_neg2_B1, simd8_op1_B1, simd8_op2_B1);
assign simd8_addcmp_out_B2 = simd8_addcmp_func(simd8_addcmp_se1_B2, simd8_addcmp_se2_B2, simd8_addcmp_neg1_B2, simd8_addcmp_neg2_B2, simd8_op1_B2, simd8_op2_B2);
assign simd8_addcmp_out_B3 = simd8_addcmp_func(simd8_addcmp_se1_B3, simd8_addcmp_se2_B3, simd8_addcmp_neg1_B3, simd8_addcmp_neg2_B3, simd8_op1_B3, simd8_op2_B3);
assign simd8_addcmp_out_B4 = simd8_addcmp_func(simd8_addcmp_se1_B4, simd8_addcmp_se2_B4, simd8_addcmp_neg1_B4, simd8_addcmp_neg2_B4, simd8_op1_B4, simd8_op2_B4);
assign simd8_addcmp_out_B5 = simd8_addcmp_func(simd8_addcmp_se1_B5, simd8_addcmp_se2_B5, simd8_addcmp_neg1_B5, simd8_addcmp_neg2_B5, simd8_op1_B5, simd8_op2_B5);
assign simd8_addcmp_out_B6 = simd8_addcmp_func(simd8_addcmp_se1_B6, simd8_addcmp_se2_B6, simd8_addcmp_neg1_B6, simd8_addcmp_neg2_B6, simd8_op1_B6, simd8_op2_B6);
assign simd8_addcmp_out_B7 = simd8_addcmp_func(simd8_addcmp_se1_B7, simd8_addcmp_se2_B7, simd8_addcmp_neg1_B7, simd8_addcmp_neg2_B7, simd8_op1_B7, simd8_op2_B7);
assign simd8_addcmp_wrap = result_simd_s_wrap8;
assign simd8_addcmp_halve = result_simd_s_halve8 | result_simd_u_halve8;
assign simd8_addcmp_s_sat = result_simd_s_sat8;
assign simd8_addcmp_u_sat = result_simd_u_sat8;
assign simd8_addcmp_result_B0 = simd8_addcmp_result(simd8_addcmp_neg2_B0, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B0, simd8_op2_B0, simd8_addcmp_out_B0);
assign simd8_addcmp_result_B1 = simd8_addcmp_result(simd8_addcmp_neg2_B1, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B1, simd8_op2_B1, simd8_addcmp_out_B1);
assign simd8_addcmp_result_B2 = simd8_addcmp_result(simd8_addcmp_neg2_B2, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B2, simd8_op2_B2, simd8_addcmp_out_B2);
assign simd8_addcmp_result_B3 = simd8_addcmp_result(simd8_addcmp_neg2_B3, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B3, simd8_op2_B3, simd8_addcmp_out_B3);
assign simd8_addcmp_result_B4 = simd8_addcmp_result(simd8_addcmp_neg2_B4, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B4, simd8_op2_B4, simd8_addcmp_out_B4);
assign simd8_addcmp_result_B5 = simd8_addcmp_result(simd8_addcmp_neg2_B5, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B5, simd8_op2_B5, simd8_addcmp_out_B5);
assign simd8_addcmp_result_B6 = simd8_addcmp_result(simd8_addcmp_neg2_B6, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B6, simd8_op2_B6, simd8_addcmp_out_B6);
assign simd8_addcmp_result_B7 = simd8_addcmp_result(simd8_addcmp_neg2_B7, function_simd_s_cmpeq8, (function_simd_s_cmplt8 | function_simd_u_cmplt8), (function_simd_s_cmple8 | function_simd_u_cmple8), (function_simd_s_min8 | function_simd_u_min8), (function_simd_s_max8 | function_simd_u_max8), function_simd_s_clip8, simd8_addcmp_wrap, simd8_addcmp_halve, simd8_addcmp_s_sat, simd8_addcmp_u_sat, simd8_op1_B7, simd8_op2_B7, simd8_addcmp_out_B7);
assign simd8_addcmp_result_64b = {simd8_addcmp_result_B7[7:0],simd8_addcmp_result_B6[7:0],simd8_addcmp_result_B5[7:0],simd8_addcmp_result_B4[7:0],simd8_addcmp_result_B3[7:0],simd8_addcmp_result_B2[7:0],simd8_addcmp_result_B1[7:0],simd8_addcmp_result_B0[7:0]};
assign simd8_addcmp_ovf_set = simd8_addcmp_result_B0[8] | simd8_addcmp_result_B1[8] | simd8_addcmp_result_B2[8] | simd8_addcmp_result_B3[8] | simd8_addcmp_result_B4[8] | simd8_addcmp_result_B5[8] | simd8_addcmp_result_B6[8] | simd8_addcmp_result_B7[8];
function  [8:0] simd8_shift;
integer i;
input is_func_slra;
input is_func_sll;
input rnd;
input sat;
input se;
input [7:0] op1;
input [3:0] amt;
reg is_pos_amt;
reg is_neg_amt;
reg is_ovf_amt;
reg is_shift_l;
reg [2:0] shift_amt;
reg [15:0] shift_l_din;
reg [15:0] shift_r_din;
reg [15:0] shift_din;
reg signed [15:0] shift_r_dout;
reg [15:0] shift_l_dout;
reg [15:0] shift_dout;
reg is_type_s_rnd;
reg is_type_s_sat;
reg s_rnd_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg [8:0] rnd_dout;
reg [7:0] result;
reg ovfout;
begin
    is_pos_amt = is_func_slra & !amt[3];
    is_neg_amt = is_func_slra & amt[3];
    is_ovf_amt = is_func_slra & (amt[3:0] == 4'd8);
    is_shift_l = is_func_sll | is_pos_amt;
    shift_amt = is_ovf_amt ? 3'd7 : is_neg_amt ? (~amt[2:0] + 3'd1) : amt[2:0];
    shift_r_din = {{7{(se & op1[7])}},op1,1'b0};
    for (i = 0; i < 16; i = i + 1) begin:gen_shift_l_din
        shift_l_din[i] = shift_r_din[15 - i];
    end
    shift_din = is_shift_l ? shift_l_din : shift_r_din;
    shift_r_dout = $signed(shift_din) >>> shift_amt;
    for (i = 0; i < 16; i = i + 1) begin:gen_shift_l_dout
        shift_l_dout[i] = shift_r_dout[15 - i];
    end
    shift_dout = is_shift_l ? shift_l_dout : shift_r_dout;
    is_type_s_rnd = is_func_slra ? (rnd & is_neg_amt) : rnd;
    is_type_s_sat = is_func_slra ? (sat & is_pos_amt) : sat;
    s_ovf_sel = is_type_s_sat & !shift_dout[15] & (shift_dout[14:8] != 7'h00);
    s_udf_sel = is_type_s_sat & shift_dout[15] & (shift_dout[14:8] != 7'h7f);
    s_rnd_sel = !(s_ovf_sel | s_udf_sel);
    rnd_dout = shift_dout[8:0] + {8'd0,is_type_s_rnd};
    result = ({8{s_rnd_sel}} & rnd_dout[8:1]) | ({8{s_ovf_sel}} & 8'h7f) | ({8{s_udf_sel}} & 8'h80);
    ovfout = s_ovf_sel | s_udf_sel;
    simd8_shift = {ovfout,result};
end
endfunction
assign simd8_shift_result_B0 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B0, dsp_data_src2[3:0]);
assign simd8_shift_result_B1 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B1, dsp_data_src2[3:0]);
assign simd8_shift_result_B2 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B2, dsp_data_src2[3:0]);
assign simd8_shift_result_B3 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B3, dsp_data_src2[3:0]);
assign simd8_shift_result_B4 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B4, dsp_data_src2[3:0]);
assign simd8_shift_result_B5 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B5, dsp_data_src2[3:0]);
assign simd8_shift_result_B6 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B6, dsp_data_src2[3:0]);
assign simd8_shift_result_B7 = simd8_shift(function_simd_s_slra8, function_simd_s_sll8, (result_simd_s_rnd8 | result_simd_s_rndsat8), (result_simd_s_sat8 | result_simd_s_rndsat8), !function_simd_u_srl8, simd8_op1_B7, dsp_data_src2[3:0]);
assign simd8_shift_result_64b = {simd8_shift_result_B7[7:0],simd8_shift_result_B6[7:0],simd8_shift_result_B5[7:0],simd8_shift_result_B4[7:0],simd8_shift_result_B3[7:0],simd8_shift_result_B2[7:0],simd8_shift_result_B1[7:0],simd8_shift_result_B0[7:0]};
assign simd8_shift_ovf_set = simd8_shift_result_B0[8] | simd8_shift_result_B1[8] | simd8_shift_result_B2[8] | simd8_shift_result_B3[8] | simd8_shift_result_B4[8] | simd8_shift_result_B5[8] | simd8_shift_result_B6[8] | simd8_shift_result_B7[8];
function  [17:0] simd8_mul_func;
input se1;
input se2;
input [7:0] op1;
input [7:0] op2;
reg [17:0] mul_in1;
reg [17:0] mul_in2;
reg signed [17:0] mul_out;
begin
    mul_in1 = {{10{(se1 & op1[7])}},op1};
    mul_in2 = {{10{(se2 & op2[7])}},op2};
    mul_out = $signed(mul_in1) * $signed(mul_in2);
    simd8_mul_func = mul_out[17:0];
end
endfunction
function  [8:0] simd8_mul_result;
input is_type_s_sat;
input [7:0] op1;
input [7:0] op2;
input [15:0] din;
reg [7:0] dout;
reg ovfout;
reg s_ovf_sel;
reg sra7_sel;
begin
    s_ovf_sel = is_type_s_sat & (op1 == 8'h80) & (op2 == 8'h80);
    sra7_sel = !s_ovf_sel;
    dout = ({8{sra7_sel}} & din[14:7]) | ({8{s_ovf_sel}} & 8'h7f);
    ovfout = s_ovf_sel;
    simd8_mul_result = {ovfout,dout};
end
endfunction
assign simd8_mul_se1_B0 = function_simd_s_mul8 | function_psimd_s_mul8x8_acc32_func0 | function_psimd_s_mul8x8_acc32_func2 | function_psimd_s_mul8x8_out64;
assign simd8_mul_se1_B1 = simd8_mul_se1_B0;
assign simd8_mul_se1_B2 = simd8_mul_se1_B0;
assign simd8_mul_se1_B3 = simd8_mul_se1_B0;
assign simd8_mul_se1_B4 = simd8_mul_se1_B0;
assign simd8_mul_se1_B5 = simd8_mul_se1_B0;
assign simd8_mul_se1_B6 = simd8_mul_se1_B0;
assign simd8_mul_se1_B7 = simd8_mul_se1_B0;
assign simd8_mul_se2_B0 = function_simd_s_mul8 | function_psimd_s_mul8x8_acc32_func0 | function_psimd_s_mul8x8_out64;
assign simd8_mul_se2_B1 = simd8_mul_se2_B0;
assign simd8_mul_se2_B2 = simd8_mul_se2_B0;
assign simd8_mul_se2_B3 = simd8_mul_se2_B0;
assign simd8_mul_se2_B4 = simd8_mul_se2_B0;
assign simd8_mul_se2_B5 = simd8_mul_se2_B0;
assign simd8_mul_se2_B6 = simd8_mul_se2_B0;
assign simd8_mul_se2_B7 = simd8_mul_se2_B0;
assign simd8_mul_out_B0 = simd8_mul_func(simd8_mul_se1_B0, simd8_mul_se2_B0, simd8_op1_B0, simd8_op2_B0);
assign simd8_mul_out_B1 = simd8_mul_func(simd8_mul_se1_B1, simd8_mul_se2_B1, simd8_op1_B1, simd8_op2_B1);
assign simd8_mul_out_B2 = simd8_mul_func(simd8_mul_se1_B2, simd8_mul_se2_B2, simd8_op1_B2, simd8_op2_B2);
assign simd8_mul_out_B3 = simd8_mul_func(simd8_mul_se1_B3, simd8_mul_se2_B3, simd8_op1_B3, simd8_op2_B3);
assign simd8_mul_out_B4 = simd8_mul_func(simd8_mul_se1_B4, simd8_mul_se2_B4, simd8_op1_B4, simd8_op2_B4);
assign simd8_mul_out_B5 = simd8_mul_func(simd8_mul_se1_B5, simd8_mul_se2_B5, simd8_op1_B5, simd8_op2_B5);
assign simd8_mul_out_B6 = simd8_mul_func(simd8_mul_se1_B6, simd8_mul_se2_B6, simd8_op1_B6, simd8_op2_B6);
assign simd8_mul_out_B7 = simd8_mul_func(simd8_mul_se1_B7, simd8_mul_se2_B7, simd8_op1_B7, simd8_op2_B7);
assign simd8_mul_s_sat = result_simd_s_sat8;
assign simd8_mul_result_B0 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B0, simd8_op2_B0, simd8_mul_out_B0[15:0]);
assign simd8_mul_result_B1 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B1, simd8_op2_B1, simd8_mul_out_B1[15:0]);
assign simd8_mul_result_B2 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B2, simd8_op2_B2, simd8_mul_out_B2[15:0]);
assign simd8_mul_result_B3 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B3, simd8_op2_B3, simd8_mul_out_B3[15:0]);
assign simd8_mul_result_B4 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B4, simd8_op2_B4, simd8_mul_out_B4[15:0]);
assign simd8_mul_result_B5 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B5, simd8_op2_B5, simd8_mul_out_B5[15:0]);
assign simd8_mul_result_B6 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B6, simd8_op2_B6, simd8_mul_out_B6[15:0]);
assign simd8_mul_result_B7 = simd8_mul_result(simd8_mul_s_sat, simd8_op1_B7, simd8_op2_B7, simd8_mul_out_B7[15:0]);
assign simd8_mul_result_64b = {simd8_mul_result_B7[7:0],simd8_mul_result_B6[7:0],simd8_mul_result_B5[7:0],simd8_mul_result_B4[7:0],simd8_mul_result_B3[7:0],simd8_mul_result_B2[7:0],simd8_mul_result_B1[7:0],simd8_mul_result_B0[7:0]};
assign simd8_mul_ovf_set = simd8_mul_result_B0[8] | simd8_mul_result_B1[8] | simd8_mul_result_B2[8] | simd8_mul_result_B3[8] | simd8_mul_result_B4[8] | simd8_mul_result_B5[8] | simd8_mul_result_B6[8] | simd8_mul_result_B7[8];
assign simd8_swap_result_64b = {simd8_op1_B6[7:0],simd8_op1_B7[7:0],simd8_op1_B4[7:0],simd8_op1_B5[7:0],simd8_op1_B2[7:0],simd8_op1_B3[7:0],simd8_op1_B0[7:0],simd8_op1_B1[7:0]};
assign simd8_swap_ovf_set = 1'b0;
function  [7:0] simd8_clz;
input is_func_clz;
input is_func_clo;
input is_func_clrs;
input [7:0] op1;
reg [7:0] clz_in_8b;
reg [3:0] clz_in_4b;
reg [2:0] clz_out;
reg clz_in_eqz;
begin
    clz_in_8b = ({8{is_func_clz}} & op1) | ({8{is_func_clo}} & ~op1) | ({8{is_func_clrs}} & ({op1[6:0],!op1[7]} ^ {8{op1[7]}}));
    clz_out[2] = (clz_in_8b[7:4] == 4'd0);
    clz_in_4b = clz_out[2] ? clz_in_8b[3:0] : clz_in_8b[7:4];
    clz_out[1] = (clz_in_4b[3:2] == 2'd0);
    clz_out[0] = clz_out[1] ? !clz_in_4b[1] : !clz_in_4b[3];
    clz_in_eqz = (clz_in_8b == 8'd0);
    simd8_clz = clz_in_eqz ? 8'd8 : {5'd0,clz_out[2:0]};
end
endfunction
assign simd8_clz_result_B0 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B0);
assign simd8_clz_result_B1 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B1);
assign simd8_clz_result_B2 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B2);
assign simd8_clz_result_B3 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B3);
assign simd8_clz_result_B4 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B4);
assign simd8_clz_result_B5 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B5);
assign simd8_clz_result_B6 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B6);
assign simd8_clz_result_B7 = simd8_clz(function_simd_s_clz8, function_simd_s_clo8, function_simd_s_clrs8, simd8_op1_B7);
assign simd8_clz_result_64b = {simd8_clz_result_B7[7:0],simd8_clz_result_B6[7:0],simd8_clz_result_B5[7:0],simd8_clz_result_B4[7:0],simd8_clz_result_B3[7:0],simd8_clz_result_B2[7:0],simd8_clz_result_B1[7:0],simd8_clz_result_B0[7:0]};
assign simd8_clz_ovf_set = 1'b0;
function  [15:0] simd8_unpack;
input se;
input en1;
input en2;
input en3;
input [7:0] op1;
input [7:0] op2;
input [7:0] op3;
reg [7:0] result_8b;
reg [15:0] result_16b;
begin
    result_8b = ({8{en1}} & op1) | ({8{en2}} & op2) | ({8{en3}} & op3);
    result_16b = {{8{(se & result_8b[7])}},result_8b};
    simd8_unpack = result_16b;
end
endfunction
assign simd8_unpack_en1_H0 = function_simd_s_unpk8_10 | function_simd_s_unpk8_20 | function_simd_s_unpk8_30;
assign simd8_unpack_en2_H0 = function_simd_s_unpk8_31;
assign simd8_unpack_en3_H0 = function_simd_s_unpk8_32;
assign simd8_unpack_en1_H1 = function_simd_s_unpk8_10;
assign simd8_unpack_en2_H1 = function_simd_s_unpk8_20;
assign simd8_unpack_en3_H1 = function_simd_s_unpk8_30 | function_simd_s_unpk8_31 | function_simd_s_unpk8_32;
assign simd8_unpack_en1_H2 = simd8_unpack_en1_H0;
assign simd8_unpack_en2_H2 = simd8_unpack_en2_H0;
assign simd8_unpack_en3_H2 = simd8_unpack_en3_H0;
assign simd8_unpack_en1_H3 = simd8_unpack_en1_H1;
assign simd8_unpack_en2_H3 = simd8_unpack_en2_H1;
assign simd8_unpack_en3_H3 = simd8_unpack_en3_H1;
assign simd8_unpack_result_H0 = simd8_unpack(result_simd_s_unpk8, simd8_unpack_en1_H0, simd8_unpack_en2_H0, simd8_unpack_en3_H0, simd8_op1_B0, simd8_op1_B1, simd8_op1_B2);
assign simd8_unpack_result_H1 = simd8_unpack(result_simd_s_unpk8, simd8_unpack_en1_H1, simd8_unpack_en2_H1, simd8_unpack_en3_H1, simd8_op1_B1, simd8_op1_B2, simd8_op1_B3);
assign simd8_unpack_result_H2 = simd8_unpack(result_simd_s_unpk8, simd8_unpack_en1_H2, simd8_unpack_en2_H2, simd8_unpack_en3_H2, simd8_op1_B4, simd8_op1_B5, simd8_op1_B6);
assign simd8_unpack_result_H3 = simd8_unpack(result_simd_s_unpk8, simd8_unpack_en1_H3, simd8_unpack_en2_H3, simd8_unpack_en3_H3, simd8_op1_B5, simd8_op1_B6, simd8_op1_B7);
assign simd8_unpack_result_64b = {simd8_unpack_result_H3[15:0],simd8_unpack_result_H2[15:0],simd8_unpack_result_H1[15:0],simd8_unpack_result_H0[15:0]};
assign simd8_unpack_ovf_set = 1'b0;
assign simd8_result_addcmp_sel = function_simd_s_add8 | function_simd_u_add8 | function_simd_s_sub8 | function_simd_u_sub8 | function_simd_s_cmpeq8 | function_simd_s_cmplt8 | function_simd_u_cmplt8 | function_simd_s_cmple8 | function_simd_u_cmple8 | function_simd_s_min8 | function_simd_u_min8 | function_simd_s_max8 | function_simd_u_max8 | function_simd_s_abs8 | function_simd_s_clip8;
assign simd8_result_shift_sel = function_simd_s_sra8 | function_simd_u_srl8 | function_simd_s_sll8 | function_simd_s_slra8;
assign simd8_result_mul_sel = function_simd_s_mul8;
assign simd8_result_swap_sel = function_simd_s_swap8;
assign simd8_result_clz_sel = function_simd_s_clz8 | function_simd_s_clo8 | function_simd_s_clrs8;
assign simd8_result_unpack_sel = function_simd_s_unpk8_10 | function_simd_s_unpk8_20 | function_simd_s_unpk8_30 | function_simd_s_unpk8_31 | function_simd_s_unpk8_32;
assign stage1_simd8_final_result_64b = ({64{simd8_result_addcmp_sel}} & simd8_addcmp_result_64b) | ({64{simd8_result_shift_sel}} & simd8_shift_result_64b) | ({64{simd8_result_mul_sel}} & simd8_mul_result_64b) | ({64{simd8_result_swap_sel}} & simd8_swap_result_64b) | ({64{simd8_result_clz_sel}} & simd8_clz_result_64b) | ({64{simd8_result_unpack_sel}} & simd8_unpack_result_64b);
assign stage1_simd8_final_ovf_set = (simd8_result_addcmp_sel & simd8_addcmp_ovf_set) | (simd8_result_shift_sel & simd8_shift_ovf_set) | (simd8_result_mul_sel & simd8_mul_ovf_set) | (simd8_result_swap_sel & simd8_swap_ovf_set) | (simd8_result_clz_sel & simd8_clz_ovf_set) | (simd8_result_unpack_sel & simd8_unpack_ovf_set);
assign psimd32_op1_base_sel = operand_psimd_op32 | operand_psimd_clip_op32 | operand_psimd_op32_op16b | operand_psimd_op32_op16t | operand_64p_opxlen | operand_simd_op32 | operand_simd_cross_op32 | operand_psimd_op32b_op32b | operand_psimd_op32b_op32t | operand_psimd_cross_op32;
assign psimd32_op1_top32_sel = operand_psimd_op32t_op32t | operand_psimd_op32t_op32b | operand_psimd_reverse_op32;
assign psimd32_op2_base_sel = operand_psimd_op32 | operand_64p_opxlen | operand_simd_op32 | operand_psimd_op32b_op32b | operand_psimd_op32t_op32b;
assign psimd32_op2_top32_sel = operand_simd_cross_op32 | operand_psimd_op32b_op32t | operand_psimd_op32t_op32t | operand_psimd_cross_op32 | operand_psimd_reverse_op32;
assign psimd32_op2_clipmin_sel_W0 = operand_psimd_clip_op32 & dsp_src1_W0[31];
assign psimd32_op2_clipmax_sel_W0 = operand_psimd_clip_op32 & !dsp_src1_W0[31];
assign psimd32_op2_clipmin_sel_W1 = operand_psimd_clip_op32 & dsp_src1_W1[31];
assign psimd32_op2_clipmax_sel_W1 = operand_psimd_clip_op32 & !dsp_src1_W1[31];
assign psimd32_op2_bottom16_sel = operand_psimd_op32_op16b;
assign psimd32_op2_top16_sel = operand_psimd_op32_op16t;
assign psimd32_op1_W0 = ({32{psimd32_op1_base_sel}} & dsp_src1_W0) | ({32{psimd32_op1_top32_sel}} & dsp_src1_W1);
assign psimd32_op2_W0 = ({32{psimd32_op2_base_sel}} & dsp_src2_W0) | ({32{psimd32_op2_top32_sel}} & dsp_src2_W1) | ({32{psimd32_op2_clipmin_sel_W0}} & dsp_clipmin_W) | ({32{psimd32_op2_clipmax_sel_W0}} & dsp_clipmax_W) | ({32{psimd32_op2_bottom16_sel}} & {{16{dsp_src2_H0[15]}},dsp_src2_H0}) | ({32{psimd32_op2_top16_sel}} & {{16{dsp_src2_H1[15]}},dsp_src2_H1});
assign psimd32_op1_W1 = ({32{psimd32_op1_base_sel}} & dsp_src1_W1) | ({32{psimd32_op1_top32_sel}} & dsp_src1_W0);
assign psimd32_op2_W1 = ({32{psimd32_op2_base_sel}} & dsp_src2_W1) | ({32{psimd32_op2_top32_sel}} & dsp_src2_W0) | ({32{psimd32_op2_clipmin_sel_W1}} & dsp_clipmin_W) | ({32{psimd32_op2_clipmax_sel_W1}} & dsp_clipmax_W) | ({32{psimd32_op2_bottom16_sel}} & {{16{dsp_src2_H2[15]}},dsp_src2_H2}) | ({32{psimd32_op2_top16_sel}} & {{16{dsp_src2_H3[15]}},dsp_src2_H3});
assign psimd32_pack_result_64b = {psimd32_op1_W0[31:0],psimd32_op2_W0[31:0]};
assign psimd32_pack_ovf_set = 1'b0;
function  [33:0] psimd32_addcmp_func;
input se1;
input se2;
input neg1;
input neg2;
input [31:0] op1;
input [31:0] op2;
reg [32:0] adder_in1;
reg [32:0] adder_in2;
reg adder_cin;
reg [32:0] adder_out;
reg cmpeq_out;
begin
    adder_in1 = {33{neg1}} ^ {(se1 & op1[31]),op1};
    adder_in2 = {33{neg2}} ^ {(se2 & op2[31]),op2};
    adder_cin = neg1 | neg2;
    adder_out = adder_in1 + adder_in2 + {32'd0,adder_cin};
    cmpeq_out = (op1 == op2);
    psimd32_addcmp_func = {cmpeq_out,adder_out};
end
endfunction
function  [32:0] psimd32_addcmp_result;
input is_func_sub;
input is_func_min;
input is_func_max;
input is_func_clip;
input is_type_wrap;
input is_type_halve;
input is_type_s_sat;
input is_type_u_sat;
input [31:0] cmp_op1;
input [31:0] cmp_op2;
input [33:0] din;
reg [31:0] dout;
reg ovfout;
reg is_eq;
reg is_lt;
reg is_le;
reg is_gt;
reg exceed_clip_bound;
reg wrap_sel;
reg halve_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg u_ovf_sel;
reg u_udf_sel;
reg cmp_op1_sel;
reg cmp_op2_sel;
begin
    is_eq = din[33];
    is_lt = din[32];
    is_le = is_eq | is_lt;
    is_gt = !is_le;
    exceed_clip_bound = is_func_clip & ((!cmp_op1[31] & is_gt) | (cmp_op1[31] & is_lt));
    halve_sel = is_type_halve;
    s_ovf_sel = is_type_s_sat & (din[32:31] == 2'b01);
    s_udf_sel = is_type_s_sat & (din[32:31] == 2'b10);
    u_ovf_sel = is_type_u_sat & din[32] & !is_func_sub;
    u_udf_sel = is_type_u_sat & din[32] & is_func_sub;
    wrap_sel = is_type_wrap | (is_type_s_sat & !(s_ovf_sel | s_udf_sel)) | (is_type_u_sat & !(u_ovf_sel | u_udf_sel));
    cmp_op1_sel = (is_func_min & din[32]) | (is_func_max & !din[32]) | (is_func_clip & !exceed_clip_bound);
    cmp_op2_sel = (is_func_min & !din[32]) | (is_func_max & din[32]) | (is_func_clip & exceed_clip_bound);
    dout = ({32{wrap_sel}} & din[31:0]) | ({32{halve_sel}} & din[32:1]) | ({32{s_ovf_sel}} & 32'h7fffffff) | ({32{s_udf_sel}} & 32'h80000000) | ({32{u_ovf_sel}} & 32'hffffffff) | ({32{u_udf_sel}} & 32'h00000000) | ({32{cmp_op1_sel}} & cmp_op1) | ({32{cmp_op2_sel}} & cmp_op2);
    ovfout = s_ovf_sel | s_udf_sel | u_ovf_sel | u_udf_sel | exceed_clip_bound;
    psimd32_addcmp_result = {ovfout,dout};
end
endfunction
assign psimd32_addcmp_se1_W0 = function_psimd_s_add32 | function_psimd_s_sub32 | function_psimd_s_min32 | function_psimd_s_max32 | function_psimd_s_abs32 | function_psimd_s_clip32 | function_simd_s_add32 | function_simd_s_sub32 | function_simd_s_as32 | function_simd_s_sa32 | function_simd_s_min32 | function_simd_s_max32 | function_simd_s_abs32;
assign psimd32_addcmp_se1_W1 = psimd32_addcmp_se1_W0;
assign psimd32_addcmp_se2_W0 = function_psimd_s_add32 | function_psimd_s_sub32 | function_psimd_s_min32 | function_psimd_s_max32 | function_psimd_s_abs32 | function_psimd_s_clip32 | function_simd_s_add32 | function_simd_s_sub32 | function_simd_s_as32 | function_simd_s_sa32 | function_simd_s_min32 | function_simd_s_max32 | function_simd_s_abs32;
assign psimd32_addcmp_se2_W1 = psimd32_addcmp_se2_W0;
assign psimd32_addcmp_neg1_W0 = (function_psimd_s_abs32 & psimd32_op1_W0[31]) | (function_simd_s_abs32 & psimd32_op1_W0[31]);
assign psimd32_addcmp_neg1_W1 = (function_psimd_s_abs32 & psimd32_op1_W1[31]) | (function_simd_s_abs32 & psimd32_op1_W1[31]);
assign psimd32_addcmp_neg2_W0 = function_psimd_s_sub32 | function_psimd_u_sub32 | function_psimd_s_min32 | function_psimd_s_max32 | function_psimd_s_clip32 | function_simd_s_sub32 | function_simd_u_sub32 | function_simd_s_as32 | function_simd_u_as32 | function_simd_s_min32 | function_simd_u_min32 | function_simd_s_max32 | function_simd_u_max32;
assign psimd32_addcmp_neg2_W1 = function_psimd_s_sub32 | function_psimd_u_sub32 | function_psimd_s_min32 | function_psimd_s_max32 | function_psimd_s_clip32 | function_simd_s_sub32 | function_simd_u_sub32 | function_simd_s_sa32 | function_simd_u_sa32 | function_simd_s_min32 | function_simd_u_min32 | function_simd_s_max32 | function_simd_u_max32;
assign psimd32_addcmp_out_W0 = psimd32_addcmp_func(psimd32_addcmp_se1_W0, psimd32_addcmp_se2_W0, psimd32_addcmp_neg1_W0, psimd32_addcmp_neg2_W0, psimd32_op1_W0, psimd32_op2_W0);
assign psimd32_addcmp_out_W1 = psimd32_addcmp_func(psimd32_addcmp_se1_W1, psimd32_addcmp_se2_W1, psimd32_addcmp_neg1_W1, psimd32_addcmp_neg2_W1, psimd32_op1_W1, psimd32_op2_W1);
assign psimd32_addcmp_min = function_psimd_s_min32 | function_simd_s_min32 | function_simd_u_min32;
assign psimd32_addcmp_max = function_psimd_s_max32 | function_simd_s_max32 | function_simd_u_max32;
assign psimd32_addcmp_clip = function_psimd_s_clip32;
assign psimd32_addcmp_wrap = result_simd_s_wrap32;
assign psimd32_addcmp_halve = result_psimd_s_halve32_sexlen | result_psimd_u_halve32_sexlen | result_simd_s_halve32 | result_simd_u_halve32;
assign psimd32_addcmp_s_sat = result_psimd_s_sat32_sexlen | result_simd_s_sat32;
assign psimd32_addcmp_u_sat = result_simd_u_sat32;
assign psimd32_addcmp_result_W0 = psimd32_addcmp_result(psimd32_addcmp_neg2_W0, psimd32_addcmp_min, psimd32_addcmp_max, psimd32_addcmp_clip, psimd32_addcmp_wrap, psimd32_addcmp_halve, psimd32_addcmp_s_sat, psimd32_addcmp_u_sat, psimd32_op1_W0, psimd32_op2_W0, psimd32_addcmp_out_W0);
assign psimd32_addcmp_result_W1 = psimd32_addcmp_result(psimd32_addcmp_neg2_W1, psimd32_addcmp_min, psimd32_addcmp_max, psimd32_addcmp_clip, psimd32_addcmp_wrap, psimd32_addcmp_halve, psimd32_addcmp_s_sat, psimd32_addcmp_u_sat, psimd32_op1_W1, psimd32_op2_W1, psimd32_addcmp_out_W1);
assign psimd32_addcmp_result32sexlen = result_psimd_s_halve32_sexlen | result_psimd_u_halve32_sexlen | result_psimd_s_sat32_sexlen | result_psimd_s_cmpsel32_sexlen;
assign psimd32_addcmp_result_64b[63:32] = psimd32_addcmp_result32sexlen ? {32{psimd32_addcmp_result_W0[31]}} : psimd32_addcmp_result_W1[31:0];
assign psimd32_addcmp_result_64b[31:0] = psimd32_addcmp_result_W0[31:0];
assign psimd32_addcmp_ovf_set = psimd32_addcmp_result_W0[32] | (!psimd32_addcmp_result32sexlen & psimd32_addcmp_result_W1[32]);
function  [31:0] psimd32_clz;
input is_func_clz;
input is_func_clo;
input is_func_clrs;
input [31:0] op1;
reg [31:0] clz_in_32b;
reg [15:0] clz_in_16b;
reg [7:0] clz_in_8b;
reg [3:0] clz_in_4b;
reg [4:0] clz_out;
reg clz_in_eqz;
begin
    clz_in_32b = ({32{is_func_clz}} & op1) | ({32{is_func_clo}} & ~op1) | ({32{is_func_clrs}} & ({op1[30:0],!op1[31]} ^ {32{op1[31]}}));
    clz_out[4] = (clz_in_32b[31:16] == 16'd0);
    clz_in_16b = clz_out[4] ? clz_in_32b[15:0] : clz_in_32b[31:16];
    clz_out[3] = (clz_in_16b[15:8] == 8'd0);
    clz_in_8b = clz_out[3] ? clz_in_16b[7:0] : clz_in_16b[15:8];
    clz_out[2] = (clz_in_8b[7:4] == 4'd0);
    clz_in_4b = clz_out[2] ? clz_in_8b[3:0] : clz_in_8b[7:4];
    clz_out[1] = (clz_in_4b[3:2] == 2'd0);
    clz_out[0] = clz_out[1] ? !clz_in_4b[1] : !clz_in_4b[3];
    clz_in_eqz = (clz_in_32b == 32'd0);
    psimd32_clz = clz_in_eqz ? 32'd32 : {27'd0,clz_out[4:0]};
end
endfunction
assign psimd32_clz_result_W0 = psimd32_clz(function_psimd_s_clz32, function_psimd_s_clo32, function_psimd_s_clrs32, psimd32_op1_W0);
assign psimd32_clz_result_W1 = psimd32_clz(function_psimd_s_clz32, function_psimd_s_clo32, function_psimd_s_clrs32, psimd32_op1_W1);
assign psimd32_clz_result_64b = {psimd32_clz_result_W1[31:0],psimd32_clz_result_W0[31:0]};
assign psimd32_clz_ovf_set = 1'b0;
function  [134:0] psimd32_mul_func;
input is_func_32x16;
input no_opovf;
input se1;
input se2;
input [31:0] op1;
input [31:0] op2;
input [66:0] wt_sum;
input [66:0] wt_cout;
reg opovf;
begin
    opovf = (!no_opovf & !is_func_32x16 & ((op1 == 32'h80000000) & (op2 == 32'h80000000))) | (!no_opovf & is_func_32x16 & ((op1 == 32'h80000000) & (op2 == 32'hffff8000)));
    psimd32_mul_func[134] = opovf;
    psimd32_mul_func[66:0] = opovf ? 67'h0_000000007fffffff : wt_sum[66:0];
    psimd32_mul_func[133:67] = opovf ? 67'h0_0000000000000000 : wt_cout[66:0];
end
endfunction
function  [175:0] stage1_psimd32_mul_result;
input bypass;
input [10:0] fctrl;
input [1:0] rctrl;
input opovf;
input [66:0] mul_sum;
input [66:0] mul_cout;
input [31:0] acc_din;
reg is_func_smmul;
reg is_func_kmmac;
reg is_func_kmmsb;
reg is_func_kwmmul;
reg is_func_maddr32;
reg is_func_msubr32;
reg is_func_smmw;
reg is_func_kmmaw;
reg is_func_kmmw2;
reg is_func_kmmaw2;
reg is_func_mulr64;
reg is_double32x32;
reg is_non_double32x32;
reg is_double32x16;
reg is_non_double32x16;
reg is_r32;
reg is_acc;
reg is_sub;
reg is_double_with_ovf;
reg is_type_s_rnd;
reg [33:0] rndacc_din1;
reg [66:0] rndacc_din2;
reg [66:0] rndacc_din3;
begin
    is_func_smmul = fctrl[0];
    is_func_kmmac = fctrl[1];
    is_func_kmmsb = fctrl[2];
    is_func_kwmmul = fctrl[3];
    is_func_maddr32 = fctrl[4];
    is_func_msubr32 = fctrl[5];
    is_func_smmw = fctrl[6];
    is_func_kmmaw = fctrl[7];
    is_func_kmmw2 = fctrl[8];
    is_func_kmmaw2 = fctrl[9];
    is_func_mulr64 = fctrl[10];
    is_double32x32 = is_func_kwmmul;
    is_non_double32x32 = is_func_smmul | is_func_kmmac | is_func_kmmsb | is_func_mulr64;
    is_double32x16 = is_func_kmmw2 | is_func_kmmaw2;
    is_non_double32x16 = is_func_smmw | is_func_kmmaw;
    is_r32 = is_func_maddr32 | is_func_msubr32;
    is_acc = is_func_kmmac | is_func_kmmsb | is_func_maddr32 | is_func_msubr32 | is_func_kmmaw | is_func_kmmaw2;
    is_sub = is_func_kmmsb | is_func_msubr32;
    is_double_with_ovf = (is_double32x32 | is_double32x16) & opovf;
    is_type_s_rnd = rctrl[1] & !is_double_with_ovf;
    rndacc_din1 = ({34{is_acc}} & {acc_din[31],acc_din[31:0],1'b0}) + (({34{(!is_sub & !is_type_s_rnd)}} & {34'd0}) | ({34{(!is_sub & is_type_s_rnd)}} & {34'd1}) | ({34{(is_sub & !is_type_s_rnd)}} & {34'd2}) | ({34{(is_sub & is_type_s_rnd)}} & {34'd1}));
    rndacc_din2 = {67{(is_sub & !bypass)}} ^ mul_sum[66:0];
    rndacc_din3 = {67{(is_sub & !bypass)}} ^ mul_cout[66:0];
    stage1_psimd32_mul_result[0] = is_double32x32;
    stage1_psimd32_mul_result[1] = is_non_double32x32;
    stage1_psimd32_mul_result[2] = is_double32x16;
    stage1_psimd32_mul_result[3] = is_non_double32x16;
    stage1_psimd32_mul_result[4] = is_r32;
    stage1_psimd32_mul_result[5] = is_acc;
    stage1_psimd32_mul_result[6] = is_sub;
    stage1_psimd32_mul_result[7] = is_double_with_ovf;
    stage1_psimd32_mul_result[41:8] = rndacc_din1;
    stage1_psimd32_mul_result[108:42] = rndacc_din2;
    stage1_psimd32_mul_result[175:109] = rndacc_din3;
end
endfunction
function  [64:0] stage2_psimd32_mul_result;
input [7:0] fctrl;
input [1:0] rctrl;
input [33:0] din1;
input [65:0] din2;
input [65:0] din3;
reg is_double32x32;
reg is_non_double32x32;
reg is_double32x16;
reg is_non_double32x16;
reg is_double_with_ovf;
reg is_r32;
reg is_sub;
reg is_type_s_sat;
reg [66:0] rndacc_din1;
reg [66:0] rndacc_din2;
reg [66:0] rndacc_din3;
reg [66:0] rndacc_dout;
reg s_ovf_sel;
reg s_udf_sel;
reg s_rndacc_sel;
reg [63:0] dout;
reg ovfout;
begin
    is_double32x32 = fctrl[0];
    is_non_double32x32 = fctrl[1];
    is_double32x16 = fctrl[2];
    is_non_double32x16 = fctrl[3];
    is_r32 = fctrl[4];
    is_sub = fctrl[6];
    is_double_with_ovf = fctrl[7];
    is_type_s_sat = rctrl[0];
    rndacc_din1 = {din1[33],din1[33:0],32'd0};
    rndacc_din2 = (({67{is_double32x32}} & {din2[64:0],is_sub,1'b0}) | ({67{is_non_double32x32}} & {din2[65:0],is_sub}) | ({67{is_double32x16}} & {din2[48:0],is_sub,17'd0}) | ({67{is_non_double32x16}} & {din2[49:0],is_sub,16'd0}) | ({67{(is_r32 | is_double_with_ovf)}} & {din2[33:0],is_sub,32'd0}));
    rndacc_din3 = (({67{is_double32x32}} & {din3[64:0],is_sub,1'b0}) | ({67{is_non_double32x32}} & {din3[65:0],is_sub}) | ({67{is_double32x16}} & {din3[48:0],is_sub,17'd0}) | ({67{is_non_double32x16}} & {din3[49:0],is_sub,16'd0}) | ({67{(is_r32 | is_double_with_ovf)}} & {din3[33:0],is_sub,32'd0}));
    rndacc_dout = csa67_1_level_add67(rndacc_din1, rndacc_din2, rndacc_din3);
    s_ovf_sel = is_type_s_sat & !rndacc_dout[66] & (rndacc_dout[65:64] != 2'b00);
    s_udf_sel = is_type_s_sat & rndacc_dout[66] & (rndacc_dout[65:64] != 2'b11);
    s_rndacc_sel = !(s_ovf_sel | s_udf_sel);
    dout[63:32] = ({32{s_rndacc_sel}} & rndacc_dout[64:33]) | ({32{s_ovf_sel}} & 32'h7fffffff) | ({32{s_udf_sel}} & 32'h80000000);
    dout[31:0] = rndacc_dout[32:1];
    ovfout = s_ovf_sel | s_udf_sel | is_double_with_ovf;
    stage2_psimd32_mul_result = {ovfout,dout};
end
endfunction
assign psimd32_mul_se1_W0 = function_psimd_s_mul32x32_acc32_func0 | function_psimd_s_mul32x32_acc32_func1 | function_psimd_s_mul32x32_acc32_func2 | function_psimd_s_mul32x32_acc32_func3 | function_psimd_s_mul32x32_acc32_func4 | function_psimd_s_mul32x32_acc32_func5 | function_psimd_s_mul32x16_acc32_func0 | function_psimd_s_mul32x16_acc32_func1 | function_psimd_s_mul32x16_acc32_func2 | function_psimd_s_mul32x16_acc32_func3 | function_psimd_s_mul32x32_out64 | function_64p_s_mul32x32_acc64_func0 | function_64p_s_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func0 | function_psimd_s_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func2 | function_psimd_s_mul32x32_acc64_func3 | function_psimd_s_mul32x32_acc64_func4 | function_psimd_s_mul32x32_acc64_func5 | function_psimd_s_mul32x32_acc64_func6;
assign psimd32_mul_se2_W0 = function_psimd_s_mul32x32_acc32_func0 | function_psimd_s_mul32x32_acc32_func1 | function_psimd_s_mul32x32_acc32_func2 | function_psimd_s_mul32x32_acc32_func3 | function_psimd_s_mul32x32_acc32_func4 | function_psimd_s_mul32x32_acc32_func5 | function_psimd_s_mul32x16_acc32_func0 | function_psimd_s_mul32x16_acc32_func1 | function_psimd_s_mul32x16_acc32_func2 | function_psimd_s_mul32x16_acc32_func3 | function_psimd_s_mul32x32_out64 | function_64p_s_mul32x32_acc64_func0 | function_64p_s_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func0 | function_psimd_s_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func2 | function_psimd_s_mul32x32_acc64_func3 | function_psimd_s_mul32x32_acc64_func4 | function_psimd_s_mul32x32_acc64_func5 | function_psimd_s_mul32x32_acc64_func6;
assign psimd32_mul_se1_W1 = psimd32_mul_se1_W0;
assign psimd32_mul_se2_W1 = psimd32_mul_se2_W0;
assign psimd32_mul_32x16 = operand_psimd_op32_op16b | operand_psimd_op32_op16t;
assign psimd32_mul_no_opovf = function_psimd_s_mul32x32_out64 | function_psimd_u_mul32x32_out64 | function_64p_s_mul32x32_acc64_func0 | function_64p_s_mul32x32_acc64_func1 | function_64p_u_mul32x32_acc64_func0 | function_64p_u_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func0 | function_psimd_s_mul32x32_acc64_func1 | function_psimd_s_mul32x32_acc64_func2 | function_psimd_s_mul32x32_acc64_func3 | function_psimd_s_mul32x32_acc64_func4 | function_psimd_s_mul32x32_acc64_func5 | function_psimd_s_mul32x32_acc64_func6 | function_psimd_s_mul32x16_acc32_func0 | function_psimd_s_mul32x16_acc32_func1 | function_psimd_s_mul32x32_acc32_func0 | function_psimd_s_mul32x32_acc32_func1 | function_psimd_s_mul32x32_acc32_func2 | function_psimd_s_mul32x32_acc32_func4 | function_psimd_s_mul32x32_acc32_func5;
kv_dsp_mul32 mul32_lv1_W0(
    .mul_op1(psimd32_op1_W0),
    .mul_op2(psimd32_op2_W0),
    .mul_op1_sign(psimd32_mul_se1_W0),
    .mul_op2_sign(psimd32_mul_se2_W0),
    .mul_wt_sum(psimd32_mul_lv1_wt_sum_W0),
    .mul_wt_cout(psimd32_mul_lv1_wt_cout_W0)
);
kv_dsp_mul32 mul32_lv1_W1(
    .mul_op1(psimd32_op1_W1),
    .mul_op2(psimd32_op2_W1),
    .mul_op1_sign(psimd32_mul_se1_W1),
    .mul_op2_sign(psimd32_mul_se2_W1),
    .mul_wt_sum(psimd32_mul_lv1_wt_sum_W1),
    .mul_wt_cout(psimd32_mul_lv1_wt_cout_W1)
);
assign psimd32_mul_lv1_out_W0 = psimd32_mul_func(psimd32_mul_32x16, psimd32_mul_no_opovf, psimd32_mul_se1_W0, psimd32_mul_se2_W0, psimd32_op1_W0, psimd32_op2_W0, psimd32_mul_lv1_wt_sum_W0, psimd32_mul_lv1_wt_cout_W0);
assign psimd32_mul_lv1_out_W1 = psimd32_mul_func(psimd32_mul_32x16, psimd32_mul_no_opovf, psimd32_mul_se1_W1, psimd32_mul_se2_W1, psimd32_op1_W1, psimd32_op2_W1, psimd32_mul_lv1_wt_sum_W1, psimd32_mul_lv1_wt_cout_W1);
assign stage2_psimd32_mul_data_en = stage2_dsp_ctrl_en & stage1_dsp_ivalid & (|stage2_psimd32_mul_fctrl_nx);
assign stage2_psimd32_mul_fctrl_nx[0] = function_psimd_s_mul32x32_acc32_func0;
assign stage2_psimd32_mul_fctrl_nx[1] = function_psimd_s_mul32x32_acc32_func1;
assign stage2_psimd32_mul_fctrl_nx[2] = function_psimd_s_mul32x32_acc32_func2;
assign stage2_psimd32_mul_fctrl_nx[3] = function_psimd_s_mul32x32_acc32_func3;
assign stage2_psimd32_mul_fctrl_nx[4] = function_psimd_s_mul32x32_acc32_func4;
assign stage2_psimd32_mul_fctrl_nx[5] = function_psimd_s_mul32x32_acc32_func5;
assign stage2_psimd32_mul_fctrl_nx[6] = function_psimd_s_mul32x16_acc32_func0;
assign stage2_psimd32_mul_fctrl_nx[7] = function_psimd_s_mul32x16_acc32_func1;
assign stage2_psimd32_mul_fctrl_nx[8] = function_psimd_s_mul32x16_acc32_func2;
assign stage2_psimd32_mul_fctrl_nx[9] = function_psimd_s_mul32x16_acc32_func3;
assign stage2_psimd32_mul_fctrl_nx[10] = function_psimd_s_mul32x32_out64 | function_psimd_u_mul32x32_out64 | function_psimd_s_mul32x32_acc64_func0;
assign stage2_psimd32_mul_fctrl_nx[11] = function_psimd_s_mul32x32_acc64_func1;
assign stage2_psimd32_mul_fctrl_nx[12] = function_psimd_s_mul32x32_acc64_func2;
assign stage2_psimd32_mul_fctrl_nx[13] = function_psimd_s_mul32x32_acc64_func3;
assign stage2_psimd32_mul_fctrl_nx[14] = function_psimd_s_mul32x32_acc64_func4 | function_64p_s_mul32x32_acc64_func0 | function_64p_u_mul32x32_acc64_func0;
assign stage2_psimd32_mul_fctrl_nx[15] = function_psimd_s_mul32x32_acc64_func5;
assign stage2_psimd32_mul_fctrl_nx[16] = function_psimd_s_mul32x32_acc64_func6 | function_64p_s_mul32x32_acc64_func1 | function_64p_u_mul32x32_acc64_func1;
assign stage2_psimd32_mul_rctrl_nx[0] = result_simd_s_sat32 | result_simd_s_rnd32_sat32;
assign stage2_psimd32_mul_rctrl_nx[1] = result_simd_s_rnd32 | result_simd_s_rnd32_sat32;
assign stage2_psimd32_mul_rctrl_nx[2] = result_psimd_s_bypass32_sexlen;
assign stage2_psimd32_mul_rctrl_nx[3] = result_64p_s_sat64 | result_psimd_s_sat64;
assign stage2_psimd32_mul_rctrl_nx[4] = result_64p_u_sat64;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd32_mul_fctrl <= 17'd0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_psimd32_mul_fctrl <= stage2_psimd32_mul_fctrl_nx;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd32_mul_rctrl <= 5'd0;
    end
    else if (stage2_psimd32_mul_data_en) begin
        stage2_psimd32_mul_rctrl <= stage2_psimd32_mul_rctrl_nx;
    end
end

assign stage2_psimd32_mul_lv1_result_W0_nx = stage1_psimd32_mul_result((|stage2_psimd32_mul_fctrl_nx[16:11]), stage2_psimd32_mul_fctrl_nx[10:0], stage2_psimd32_mul_rctrl_nx[1:0], psimd32_mul_lv1_out_W0[134], psimd32_mul_lv1_out_W0[66:0], psimd32_mul_lv1_out_W0[133:67], stage1_acc_din_W0);
assign stage2_psimd32_mul_lv1_result_W1_nx = stage1_psimd32_mul_result((|stage2_psimd32_mul_fctrl_nx[16:11]), stage2_psimd32_mul_fctrl_nx[10:0], stage2_psimd32_mul_rctrl_nx[1:0], psimd32_mul_lv1_out_W1[134], psimd32_mul_lv1_out_W1[66:0], psimd32_mul_lv1_out_W1[133:67], stage1_acc_din_W1);
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd32_mul_lv1_result_W0 <= 176'd0;
        stage2_psimd32_mul_lv1_result_W1 <= 176'd0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_psimd32_mul_lv1_result_W0 <= stage2_psimd32_mul_lv1_result_W0_nx;
        stage2_psimd32_mul_lv1_result_W1 <= stage2_psimd32_mul_lv1_result_W1_nx;
    end
end

assign stage2_psimd32_mul_result_W0 = stage2_psimd32_mul_result(stage2_psimd32_mul_lv1_result_W0[7:0], stage2_psimd32_mul_rctrl[1:0], stage2_psimd32_mul_lv1_result_W0[41:8], stage2_psimd32_mul_lv1_result_W0[107:42], stage2_psimd32_mul_lv1_result_W0[174:109]);
assign stage2_psimd32_mul_result_W1 = stage2_psimd32_mul_result(stage2_psimd32_mul_lv1_result_W1[7:0], stage2_psimd32_mul_rctrl[1:0], stage2_psimd32_mul_lv1_result_W1[41:8], stage2_psimd32_mul_lv1_result_W1[107:42], stage2_psimd32_mul_lv1_result_W1[174:109]);
assign stage2_psimd32_mul_result32sexlen = stage2_psimd32_mul_rctrl[2];
assign stage2_psimd32_mul_resultout64 = stage2_psimd32_mul_fctrl[10];
assign stage2_psimd32_mul_result_64b[63:32] = stage2_psimd32_mul_result32sexlen ? {32{stage2_psimd32_mul_result_W0[63]}} : stage2_psimd32_mul_resultout64 ? stage2_psimd32_mul_result_W0[63:32] : stage2_psimd32_mul_result_W1[63:32];
assign stage2_psimd32_mul_result_64b[31:0] = stage2_psimd32_mul_resultout64 ? stage2_psimd32_mul_result_W0[31:0] : stage2_psimd32_mul_result_W0[63:32];
assign stage2_psimd32_mul_ovf_set = stage2_psimd32_mul_result32sexlen ? stage2_psimd32_mul_result_W0[64] : stage2_psimd32_mul_resultout64 ? 1'b0 : (stage2_psimd32_mul_result_W0[64] | stage2_psimd32_mul_result_W1[64]);
assign stage3_psimd32_mul_data_en = stage3_dsp_ctrl_en & stage2_dsp_ivalid & (|stage3_psimd32_mul_fctrl_nx);
assign stage3_psimd32_mul_fctrl_nx[5:0] = stage2_psimd32_mul_fctrl[16:11];
assign stage3_psimd32_mul_rctrl_nx[1:0] = stage2_psimd32_mul_rctrl[4:3];
assign stage3_psimd32_mul_out1_nx = stage2_profile64_mul_csa_out1;
assign stage3_psimd32_mul_out2_nx = stage2_profile64_mul_csa_out2;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_psimd32_mul_fctrl <= 6'd0;
    end
    else if (stage3_dsp_ctrl_en) begin
        stage3_psimd32_mul_fctrl <= stage3_psimd32_mul_fctrl_nx;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_psimd32_mul_rctrl <= 2'd0;
        stage3_psimd32_mul_out1 <= 67'd0;
        stage3_psimd32_mul_out2 <= 67'd0;
    end
    else if (stage3_psimd32_mul_data_en) begin
        stage3_psimd32_mul_rctrl <= stage3_psimd32_mul_rctrl_nx;
        stage3_psimd32_mul_out1 <= stage3_psimd32_mul_out1_nx;
        stage3_psimd32_mul_out2 <= stage3_psimd32_mul_out2_nx;
    end
end

assign stage3_psimd32_mul_result_64b = stage3_profile64_mul_result_64b;
assign stage3_psimd32_mul_ovf_set = stage3_profile64_mul_ovf_set;
assign psimd32_result_addcmp_sel = function_psimd_s_add32 | function_psimd_u_add32 | function_psimd_s_sub32 | function_psimd_u_sub32 | function_psimd_s_min32 | function_psimd_s_max32 | function_psimd_s_abs32 | function_psimd_s_clip32 | function_simd_s_add32 | function_simd_u_add32 | function_simd_s_sub32 | function_simd_u_sub32 | function_simd_s_as32 | function_simd_u_as32 | function_simd_s_sa32 | function_simd_u_sa32 | function_simd_s_min32 | function_simd_u_min32 | function_simd_s_max32 | function_simd_u_max32 | function_simd_s_abs32;
assign psimd32_result_clz_sel = function_psimd_s_clz32 | function_psimd_s_clo32 | function_psimd_s_clrs32;
assign psimd32_result_pack_sel = function_psimd_s_pk32;
assign stage1_psimd32_final_result_64b = ({64{psimd32_result_addcmp_sel}} & psimd32_addcmp_result_64b) | ({64{psimd32_result_clz_sel}} & psimd32_clz_result_64b) | ({64{psimd32_result_pack_sel}} & psimd32_pack_result_64b);
assign stage1_psimd32_final_ovf_set = (psimd32_result_addcmp_sel & psimd32_addcmp_ovf_set) | (psimd32_result_clz_sel & psimd32_clz_ovf_set) | (psimd32_result_pack_sel & psimd32_pack_ovf_set);
assign stage2_psimd32_result_mul_sel = (|stage2_psimd32_mul_fctrl[10:0]);
assign stage2_psimd32_final_result_64b = ({64{stage2_psimd32_result_mul_sel}} & stage2_psimd32_mul_result_64b);
assign stage2_psimd32_final_ovf_set = (stage2_psimd32_result_mul_sel & stage2_psimd32_mul_ovf_set);
assign stage3_psimd32_result_mul_sel = (|stage3_psimd32_mul_fctrl);
assign stage3_psimd32_final_result_64b = ({64{stage3_psimd32_result_mul_sel}} & stage3_psimd32_mul_result_64b);
assign stage3_psimd32_final_ovf_set = (stage3_psimd32_result_mul_sel & stage3_psimd32_mul_ovf_set);
assign psimdxlen_op1_base_sel = operand_psimd_opxlen | operand_nsimd_op32 | operand_simd_op32;
assign psimdxlen_op1_pair_sel = operand_psimd_op64;
assign psimdxlen_op2_base_sel = operand_psimd_opxlen | operand_nsimd_op32 | operand_simd_op32;
assign psimdxlen_op2_pair_sel = operand_psimd_op64;
assign psimdxlen_op3_base_sel = operand_psimd_opxlen;
assign psimdxlen_op1_64b = ({64{psimdxlen_op1_base_sel}} & dsp_src1_64b_simd) | ({64{psimdxlen_op1_pair_sel}} & dsp_src1_64b_pair);
assign psimdxlen_op2_64b = ({64{psimdxlen_op2_base_sel}} & dsp_src2_64b_simd) | ({64{psimdxlen_op2_pair_sel}} & dsp_src2_64b_pair);
assign psimdxlen_op3_64b = ({64{psimdxlen_op3_base_sel}} & dsp_src3_64b_simd);
function  [64:0] psimdxlen_shift;
integer i;
input is_func_sra;
input is_func_sll;
input is_func_bitrev;
input is_func_wext;
input is_func_slra32;
input is_func_sra32;
input is_func_srl32;
input is_func_sll32;
input rnd;
input sat;
input [63:0] op1;
input [5:0] amt;
reg is_slra32_sra;
reg is_slra32_sll;
reg is_shift_l;
reg is_se;
reg is_shift32;
reg slra32_sra_amt_sel;
reg bitrev_amt_sel;
reg [5:0] slra32_sra_shift_amt;
reg [SHIFT_AMT_MSB:0] bitrev_shift_amt;
reg [5:0] base_shift_amt;
reg [SHIFT_AMT_MSB:0] shift_amt;
reg bitrev32_din_sel;
reg shift32_din_sel;
reg [64:0] bitrev32_din;
reg [64:0] shift32_din;
reg [64:0] shift64_din;
reg [64:0] shift_r_din;
reg [64:0] shift_l_din;
reg [64:0] shift_din;
reg signed [64:0] shift_r_dout;
reg [64:0] shift_l_dout;
reg [64:0] shift_dout;
reg is_type_s_rnd;
reg is_type_s_sat;
reg s_rnd_sel;
reg s_shift32_sel;
reg u_bitrev_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg [63:0] shift32_dout;
reg [63:0] bitrev_dout;
reg [64:0] rnd_dout;
reg [63:0] result;
reg ovfout;
begin
    is_slra32_sra = is_func_slra32 & amt[5];
    is_slra32_sll = is_func_slra32 & !amt[5];
    is_shift_l = is_func_sll | is_slra32_sll | is_func_sll32;
    is_se = is_func_sll | is_func_sra | is_func_wext | is_func_slra32 | is_func_sll32 | is_func_sra32;
    is_shift32 = (is_func_sra32) | is_func_srl32 | is_func_sll32;
    slra32_sra_amt_sel = is_slra32_sra;
    bitrev_amt_sel = is_func_bitrev;
    slra32_sra_shift_amt = (amt[5:0] == 6'd32) ? 6'd31 : (~amt[5:0] + 6'd1);
    bitrev_shift_amt = {(SHIFT_AMT_MSB + 1){1'b1}} + ~amt[SHIFT_AMT_MSB:0] + {{SHIFT_AMT_MSB{1'b0}},1'b1};
    base_shift_amt = {(amt[5] & !is_shift32),amt[4:0]};
    shift_amt = slra32_sra_amt_sel ? slra32_sra_shift_amt[SHIFT_AMT_MSB:0] : bitrev_amt_sel ? bitrev_shift_amt[SHIFT_AMT_MSB:0] : base_shift_amt[SHIFT_AMT_MSB:0];
    bitrev32_din_sel = is_func_bitrev;
    shift32_din_sel = !is_func_wext | (is_shift_l & (|amt[4:0])) | is_func_slra32 | is_func_sra32 | is_func_srl32 | is_func_sll32;
    bitrev32_din = {op1[31:0],32'd0,1'b0};
    shift32_din = {{32{(is_se & op1[31])}},op1[31:0],1'b0};
    shift64_din = {op1[63:0],1'b0};
    shift_r_din = bitrev32_din_sel ? bitrev32_din : shift32_din_sel ? shift32_din : shift64_din;
    for (i = 0; i < 65; i = i + 1) begin:gen_shift_l_din
        shift_l_din[i] = shift_r_din[64 - i];
    end
    shift_din = (is_shift_l | is_func_bitrev) ? shift_l_din : shift_r_din;
    shift_r_dout = $signed(shift_din) >>> shift_amt;
    for (i = 0; i < 65; i = i + 1) begin:gen_shift_l_dout
        shift_l_dout[i] = shift_r_dout[64 - i];
    end
    shift_dout = is_shift_l ? shift_l_dout : shift_r_dout;
    is_type_s_rnd = is_func_slra32 ? (rnd & is_slra32_sra) : rnd;
    is_type_s_sat = is_func_slra32 ? (sat & is_slra32_sll) : (sat & (|shift_amt));
    s_ovf_sel = is_type_s_sat & !shift_dout[64] & (shift_dout[63:32] != 32'h00000000);
    s_udf_sel = is_type_s_sat & shift_dout[64] & (shift_dout[63:32] != 32'hffffffff);
    s_shift32_sel = (is_shift_l & (|{shift_amt,is_slra32_sll}) & !(s_ovf_sel | s_udf_sel)) | is_func_wext;
    u_bitrev_sel = is_func_bitrev;
    s_rnd_sel = is_type_s_rnd | !(is_type_s_sat | is_func_bitrev | is_func_wext);
    shift32_dout = {{32{shift_dout[32]}},shift_dout[32:1]};
    bitrev_dout = shift_dout[63:0];
    rnd_dout = shift_dout + {64'd0,is_type_s_rnd};
    result = ({64{s_rnd_sel}} & rnd_dout[64:1]) | ({64{s_shift32_sel}} & shift32_dout[63:0]) | ({64{u_bitrev_sel}} & bitrev_dout[63:0]) | ({64{s_ovf_sel}} & 64'h000000007fffffff) | ({64{s_udf_sel}} & 64'hffffffff80000000);
    ovfout = s_ovf_sel | s_udf_sel;
    psimdxlen_shift = {ovfout,result};
end
endfunction
assign psimdxlen_shift_s_rnd = result_psimd_s_rndxlen | result_nsimd_s_rnd32_se64 | result_nsimd_s_rndsat32_sexlen | result_simd_s_rnd32 | result_simd_s_rndsat32;
assign psimdxlen_shift_s_sat = result_psimd_s_sat32_sexlen | result_nsimd_s_sat32_sexlen | result_nsimd_s_rndsat32_sexlen | result_simd_s_sat32 | result_simd_s_rndsat32;
assign psimdxlen_shift_result_W0XLEN = psimdxlen_shift(function_psimd_s_sraxlen, 1'b0, function_psimd_u_bitrevxlen, function_psimd_s_wext32, (function_nsimd_s_slra32 | function_simd_s_slra32), (function_nsimd_s_sra32 | function_simd_s_sra32), function_simd_u_srl32, (function_psimd_s_sll32 | function_simd_s_sll32), psimdxlen_shift_s_rnd, psimdxlen_shift_s_sat, psimdxlen_op1_64b, dsp_data_src2[5:0]);
assign psimdxlen_shift_result_W1 = psimdxlen_shift(1'b0, 1'b0, 1'b0, 1'b0, function_simd_s_slra32, function_simd_s_sra32, function_simd_u_srl32, function_simd_s_sll32, psimdxlen_shift_s_rnd, psimdxlen_shift_s_sat, {32'd0,dsp_src1_W1}, dsp_data_src2[5:0]);
assign psimdxlen_shift_result32 = result_simd_s_bypass32 | result_simd_s_rnd32 | result_simd_s_sat32 | result_simd_s_rndsat32;
assign psimdxlen_shift_result_64b[63:32] = psimdxlen_shift_result32 ? psimdxlen_shift_result_W1[31:0] : psimdxlen_shift_result_W0XLEN[63:32];
assign psimdxlen_shift_result_64b[31:0] = psimdxlen_shift_result_W0XLEN[31:0];
assign psimdxlen_shift_ovf_set = psimdxlen_shift_result_W0XLEN[64] | (psimdxlen_shift_result32 & psimdxlen_shift_result_W1[64]);
always @* begin
    for (i = 0; i < 64; i = i + 1) begin
        psimdxlen_bpick_result_64b[i] = psimdxlen_op3_64b[i] ? psimdxlen_op1_64b[i] : psimdxlen_op2_64b[i];
    end
end

assign psimdxlen_bpick_ovf_set = 1'b0;
assign psimdxlen_insb_byte_sel = 8'd1 << {1'b0,dsp_data_src2[1:0]};
assign psimdxlen_insb_result_B0 = psimdxlen_insb_byte_sel[0] ? dsp_src1_B0 : dsp_src3_B0;
assign psimdxlen_insb_result_B1 = psimdxlen_insb_byte_sel[1] ? dsp_src1_B0 : dsp_src3_B1;
assign psimdxlen_insb_result_B2 = psimdxlen_insb_byte_sel[2] ? dsp_src1_B0 : dsp_src3_B2;
assign psimdxlen_insb_result_B3 = psimdxlen_insb_byte_sel[3] ? dsp_src1_B0 : dsp_src3_B3;
assign psimdxlen_insb_result_B4 = psimdxlen_insb_byte_sel[4] ? dsp_src1_B0 : dsp_src3_B4;
assign psimdxlen_insb_result_B5 = psimdxlen_insb_byte_sel[5] ? dsp_src1_B0 : dsp_src3_B5;
assign psimdxlen_insb_result_B6 = psimdxlen_insb_byte_sel[6] ? dsp_src1_B0 : dsp_src3_B6;
assign psimdxlen_insb_result_B7 = psimdxlen_insb_byte_sel[7] ? dsp_src1_B0 : dsp_src3_B7;
assign psimdxlen_insb_result_64b = {psimdxlen_insb_result_B7[7:0],psimdxlen_insb_result_B6[7:0],psimdxlen_insb_result_B5[7:0],psimdxlen_insb_result_B4[7:0],psimdxlen_insb_result_B3[7:0],psimdxlen_insb_result_B2[7:0],psimdxlen_insb_result_B1[7:0],psimdxlen_insb_result_B0[7:0]};
assign psimdxlen_insb_ovf_set = 1'b0;
assign psimdxlen_result_shift_sel = function_psimd_s_sraxlen | function_psimd_s_sll32 | function_psimd_u_bitrevxlen | function_psimd_s_wext32 | function_nsimd_s_sra32 | function_nsimd_s_slra32 | function_simd_s_slra32 | function_simd_s_sra32 | function_simd_u_srl32 | function_simd_s_sll32;
assign psimdxlen_result_bpick_sel = function_psimd_s_bpickxlen;
assign psimdxlen_result_insb_sel = function_psimd_s_insbxlen;
assign stage1_psimdxlen_final_result_64b = ({64{psimdxlen_result_shift_sel}} & psimdxlen_shift_result_64b) | ({64{psimdxlen_result_bpick_sel}} & psimdxlen_bpick_result_64b) | ({64{psimdxlen_result_insb_sel}} & psimdxlen_insb_result_64b);
assign stage1_psimdxlen_final_ovf_set = (psimdxlen_result_shift_sel & psimdxlen_shift_ovf_set) | (psimdxlen_result_bpick_sel & psimdxlen_bpick_ovf_set) | (psimdxlen_result_insb_sel & psimdxlen_insb_ovf_set);
assign psimd16_op1_bottom_sel = operand_psimd_op16 | operand_psimd_op16b_op16b | operand_psimd_op16b_op16t | operand_psimd_cross_op16;
assign psimd16_op1_top_sel = operand_psimd_op16 | operand_psimd_op16t_op16b | operand_psimd_op16t_op16t;
assign psimd16_op2_bottom_sel = operand_psimd_op16 | operand_psimd_op16b_op16b | operand_psimd_op16t_op16b;
assign psimd16_op2_top_sel = operand_psimd_op16 | operand_psimd_op16b_op16t | operand_psimd_op16t_op16t | operand_psimd_cross_op16;
assign psimd16_op1_H0 = ({16{psimd16_op1_bottom_sel}} & dsp_src1_H0) | ({16{psimd16_op1_top_sel}} & dsp_src1_H1);
assign psimd16_op2_H0 = ({16{psimd16_op2_bottom_sel}} & dsp_src2_H0) | ({16{psimd16_op2_top_sel}} & dsp_src2_H1);
assign psimd16_op1_H2 = ({16{psimd16_op1_bottom_sel}} & dsp_src1_H2) | ({16{psimd16_op1_top_sel}} & dsp_src1_H3);
assign psimd16_op2_H2 = ({16{psimd16_op2_bottom_sel}} & dsp_src2_H2) | ({16{psimd16_op2_top_sel}} & dsp_src2_H3);
assign psimd16_pack_result_64b = {psimd16_op1_H2[15:0],psimd16_op2_H2[15:0],psimd16_op1_H0[15:0],psimd16_op2_H0[15:0]};
assign psimd16_pack_ovf_set = 1'b0;
function  [33:0] csa34_2_level_add34;
integer i;
input [33:0] din1;
input [33:0] din2;
input [33:0] din3;
input [33:0] din4;
reg [33:0] lv1_csa1_din1;
reg [33:0] lv1_csa1_din2;
reg [33:0] lv1_csa1_din3;
reg [33:0] lv1_csa1_dout1;
reg [33:0] lv1_csa1_dout2;
reg [33:0] lv2_csa1_din1;
reg [33:0] lv2_csa1_din2;
reg [33:0] lv2_csa1_din3;
reg [33:0] lv2_csa1_dout1;
reg [33:0] lv2_csa1_dout2;
reg [33:0] add_dout;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 34; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    lv2_csa1_din1 = lv1_csa1_dout1;
    lv2_csa1_din2 = {lv1_csa1_dout2[32:0],1'b0};
    lv2_csa1_din3 = din4;
    for (i = 0; i < 34; i = i + 1) begin
        {lv2_csa1_dout2[i],lv2_csa1_dout1[i]} = {1'b0,lv2_csa1_din1[i]} + {1'b0,lv2_csa1_din2[i]} + {1'b0,lv2_csa1_din3[i]};
    end
    add_dout = {lv2_csa1_dout2[32:0],1'b0} + lv2_csa1_dout1[33:0];
    csa34_2_level_add34 = add_dout;
end
endfunction
function  [63:0] csa64_1_level_add64;
integer i;
input [63:0] din1;
input [63:0] din2;
input [63:0] din3;
reg [63:0] lv1_csa1_din1;
reg [63:0] lv1_csa1_din2;
reg [63:0] lv1_csa1_din3;
reg [63:0] lv1_csa1_dout1;
reg [63:0] lv1_csa1_dout2;
reg [63:0] add_dout;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 64; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    add_dout = {lv1_csa1_dout2[62:0],1'b0} + lv1_csa1_dout1[63:0];
    csa64_1_level_add64 = add_dout;
end
endfunction
function  [66:0] csa67_1_level_add67;
integer i;
input [66:0] din1;
input [66:0] din2;
input [66:0] din3;
reg [66:0] lv1_csa1_din1;
reg [66:0] lv1_csa1_din2;
reg [66:0] lv1_csa1_din3;
reg [66:0] lv1_csa1_dout1;
reg [66:0] lv1_csa1_dout2;
reg [66:0] add_dout;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 67; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    add_dout = {lv1_csa1_dout2[65:0],1'b0} + lv1_csa1_dout1[66:0];
    csa67_1_level_add67 = add_dout;
end
endfunction
function  [34:0] stage2_psimd16_mul_result;
input [10:0] fctrl;
input rctrl;
input opovf;
input [31:0] mul_din1;
input [31:0] mul_din2;
input [31:0] acc_din;
input acc_sign;
reg is_func_kmda;
reg is_func_smds;
reg is_func_kma;
reg is_func_kmada;
reg is_func_kmads;
reg is_func_kmsda;
reg is_func_kdma;
reg is_func_smal;
reg is_func_smalda;
reg is_func_smalds;
reg is_func_smslda;
reg is_type_s_sat;
reg acc_din1_en;
reg acc_din2_en;
reg acc_din3_en;
reg acc_din2_sub;
reg acc_din3_sub;
reg [33:0] acc_din1;
reg [33:0] acc_din2;
reg [33:0] acc_din3;
reg [33:0] acc_din4;
reg [33:0] acc_dout;
reg s_ovf_sel;
reg s_udf_sel;
reg s_acc_sel;
reg [33:0] dout;
reg ovfout;
begin
    is_func_kmda = fctrl[0];
    is_func_smds = fctrl[1];
    is_func_kma = fctrl[2];
    is_func_kmada = fctrl[3];
    is_func_kmads = fctrl[4];
    is_func_kmsda = fctrl[5];
    is_func_kdma = fctrl[6];
    is_func_smal = fctrl[7];
    is_func_smalda = fctrl[8];
    is_func_smalds = fctrl[9];
    is_func_smslda = fctrl[10];
    is_type_s_sat = rctrl;
    acc_din1_en = is_func_kma | is_func_kmada | is_func_kmads | is_func_kmsda | is_func_kdma;
    acc_din2_en = is_func_kmda | is_func_smds | is_func_kmada | is_func_kmads | is_func_kmsda | is_func_smalda | is_func_smalds | is_func_smslda;
    acc_din3_en = is_func_kmda | is_func_smds | is_func_kma | is_func_kmada | is_func_kmads | is_func_kmsda | is_func_smal | is_func_smalda | is_func_smalds | is_func_smslda | is_func_kdma;
    acc_din2_sub = is_func_kmsda | is_func_smslda;
    acc_din3_sub = is_func_smds | is_func_kmads | is_func_kmsda | is_func_smalds | is_func_smslda;
    acc_din1 = {34{acc_din1_en}} & {{2{(acc_sign & acc_din[31])}},acc_din[31:0]};
    acc_din2 = {34{acc_din2_sub}} ^ {34{acc_din2_en}} & {{2{mul_din1[31]}},mul_din1[31:0]};
    acc_din3 = {34{acc_din3_sub}} ^ {34{acc_din3_en}} & {{2{mul_din2[31]}},mul_din2[31:0]};
    acc_din4[33:0] = {32'd0,({1'b0,acc_din2_sub} + {1'b0,acc_din3_sub})};
    acc_dout = csa34_2_level_add34(acc_din1, acc_din2, acc_din3, acc_din4);
    s_ovf_sel = is_type_s_sat & !acc_dout[33] & (acc_dout[32:31] != 2'b00);
    s_udf_sel = is_type_s_sat & acc_dout[33] & (acc_dout[32:31] != 2'b11);
    s_acc_sel = !(s_ovf_sel | s_udf_sel);
    dout = ({34{s_acc_sel}} & acc_dout[33:0]) | ({34{s_ovf_sel}} & 34'h0_7fffffff) | ({34{s_udf_sel}} & 34'h3_80000000);
    ovfout = s_ovf_sel | s_udf_sel | opovf;
    stage2_psimd16_mul_result = {ovfout,dout};
end
endfunction
function  [63:0] stage3_psimd16_mul_result;
input [3:0] fctrl;
input rctrl;
input [33:0] mul_din1;
input [33:0] mul_din2;
input [63:0] acc_din;
reg is_func_smal;
reg is_func_smalda;
reg is_func_smalds;
reg is_func_smslda;
reg acc_din1_en;
reg acc_din2_en;
reg acc_din3_en;
reg [63:0] acc_din1;
reg [63:0] acc_din2;
reg [63:0] acc_din3;
reg [63:0] acc_dout;
reg s_acc_sel;
reg [63:0] dout;
begin
    is_func_smal = fctrl[0];
    is_func_smalda = fctrl[1];
    is_func_smalds = fctrl[2];
    is_func_smslda = fctrl[3];
    acc_din1_en = is_func_smal | is_func_smalda | is_func_smalds | is_func_smslda;
    acc_din2_en = is_func_smal | is_func_smalda | is_func_smalds | is_func_smslda;
    acc_din3_en = is_func_smal | is_func_smalda | is_func_smalds | is_func_smslda;
    acc_din1 = {64{acc_din1_en}} & {acc_din[63:0]};
    acc_din2 = {64{acc_din2_en}} & {{30{mul_din1[33]}},mul_din1[33:0]};
    acc_din3 = {64{acc_din3_en}} & {{30{mul_din2[33]}},mul_din2[33:0]};
    acc_dout = csa64_1_level_add64(acc_din1, acc_din2, acc_din3);
    s_acc_sel = !rctrl;
    dout = ({64{s_acc_sel}} & acc_dout[63:0]);
    stage3_psimd16_mul_result = dout;
end
endfunction
assign stage1_psimd16_mul_out_H0 = simd16_mul_out_H0;
assign stage1_psimd16_mul_out_H1 = simd16_mul_out_H1;
assign stage1_psimd16_mul_out_H2 = simd16_mul_out_H2;
assign stage1_psimd16_mul_out_H3 = simd16_mul_out_H3;
assign stage1_is_mul16x16_out64 = function_psimd_s_mul16x16_out64 | function_psimd_u_mul16x16_out64;
assign stage1_psimd16_mul_result_64b[63:32] = stage1_is_mul16x16_out64 ? stage1_psimd16_mul_out_H1 : stage1_psimd16_mul_out_H2;
assign stage1_psimd16_mul_result_64b[31:0] = stage1_psimd16_mul_out_H0;
assign stage1_psimd16_mul_ovf_set = 1'b0;
assign stage2_psimd16_mul_data_en = stage2_dsp_ctrl_en & stage1_dsp_ivalid & (|stage2_psimd16_mul_fctrl_nx);
assign stage2_psimd16_mul_fctrl_nx[0] = function_psimd_s_mul16x16_acc32_func1;
assign stage2_psimd16_mul_fctrl_nx[1] = function_psimd_s_mul16x16_acc32_func2;
assign stage2_psimd16_mul_fctrl_nx[2] = function_psimd_s_mul16x16_acc32_func3;
assign stage2_psimd16_mul_fctrl_nx[3] = function_psimd_s_mul16x16_acc32_func4 | function_psimd_s_mul8x8_acc32;
assign stage2_psimd16_mul_fctrl_nx[4] = function_psimd_s_mul16x16_acc32_func5;
assign stage2_psimd16_mul_fctrl_nx[5] = function_psimd_s_mul16x16_acc32_func6;
assign stage2_psimd16_mul_fctrl_nx[6] = function_nsimd_s_mul16x16_double32_acc32;
assign stage2_psimd16_mul_fctrl_nx[7] = function_psimd_s_mul16x16_acc64_func0 | function_64p_s_mul16x16_acc64_func0;
assign stage2_psimd16_mul_fctrl_nx[8] = function_64p_s_mul16x16_acc64_func1;
assign stage2_psimd16_mul_fctrl_nx[9] = function_64p_s_mul16x16_acc64_func2;
assign stage2_psimd16_mul_fctrl_nx[10] = function_64p_s_mul16x16_acc64_func3;
assign stage2_psimd16_mul_rctrl_nx[0] = result_psimd_s_sat32 | result_nsimd_s_sat32;
assign stage2_psimd16_mul_rctrl_nx[1] = result_nsimd_s_sat32_sexlen;
assign stage2_psimd16_mul_out_H0_nx = function_psimd_s_mul8x8_acc32 ? {{12{stage1_psimd8_mul_out_W0[19]}},stage1_psimd8_mul_out_W0[19:0]} : function_nsimd_s_mul16x16_double32_acc32 ? nsimd16_mul_result_H0[31:0] : stage1_psimd16_mul_out_H0;
assign stage2_psimd16_mul_out_H1_nx = function_psimd_s_mul8x8_acc32 ? {{12{stage1_psimd8_mul_out_W0[39]}},stage1_psimd8_mul_out_W0[39:20]} : stage1_psimd16_mul_out_H1;
assign stage2_psimd16_mul_out_H2_nx = function_psimd_s_mul8x8_acc32 ? {{12{stage1_psimd8_mul_out_W1[19]}},stage1_psimd8_mul_out_W1[19:0]} : function_nsimd_s_mul16x16_double32_acc32 ? nsimd16_mul_result_H2[31:0] : stage1_psimd16_mul_out_H2;
assign stage2_psimd16_mul_out_H3_nx = function_psimd_s_mul8x8_acc32 ? {{12{stage1_psimd8_mul_out_W1[39]}},stage1_psimd8_mul_out_W1[39:20]} : stage1_psimd16_mul_out_H3;
assign stage2_psimd16_opovf_H0_nx = nsimd16_mul_result_H0[32];
assign stage2_psimd16_opovf_H2_nx = nsimd16_mul_result_H2[32];
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd16_mul_fctrl <= 11'd0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_psimd16_mul_fctrl <= stage2_psimd16_mul_fctrl_nx;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd16_mul_rctrl <= 2'd0;
        stage2_psimd16_mul_out_H0 <= 32'd0;
        stage2_psimd16_mul_out_H1 <= 32'd0;
        stage2_psimd16_mul_out_H2 <= 32'd0;
        stage2_psimd16_mul_out_H3 <= 32'd0;
        stage2_psimd16_opovf_H0 <= 1'b0;
        stage2_psimd16_opovf_H2 <= 1'b0;
    end
    else if (stage2_psimd16_mul_data_en) begin
        stage2_psimd16_mul_rctrl <= stage2_psimd16_mul_rctrl_nx;
        stage2_psimd16_mul_out_H0 <= stage2_psimd16_mul_out_H0_nx;
        stage2_psimd16_mul_out_H1 <= stage2_psimd16_mul_out_H1_nx;
        stage2_psimd16_mul_out_H2 <= stage2_psimd16_mul_out_H2_nx;
        stage2_psimd16_mul_out_H3 <= stage2_psimd16_mul_out_H3_nx;
        stage2_psimd16_opovf_H0 <= stage2_psimd16_opovf_H0_nx;
        stage2_psimd16_opovf_H2 <= stage2_psimd16_opovf_H2_nx;
    end
end

assign stage2_psimd16_mul_result_W0 = stage2_psimd16_mul_result(stage2_psimd16_mul_fctrl, (|stage2_psimd16_mul_rctrl), stage2_psimd16_opovf_H0, stage2_psimd16_mul_out_H1, stage2_psimd16_mul_out_H0, stage2_acc_din_W0, stage2_acc_din_sign);
assign stage2_psimd16_mul_result_W1 = stage2_psimd16_mul_result(stage2_psimd16_mul_fctrl, (|stage2_psimd16_mul_rctrl), stage2_psimd16_opovf_H2, stage2_psimd16_mul_out_H3, stage2_psimd16_mul_out_H2, stage2_acc_din_W1, stage2_acc_din_sign);
assign stage2_psimd16_mul_result32sexlen = stage2_psimd16_mul_rctrl[1];
assign stage2_psimd16_mul_result_64b[63:32] = stage2_psimd16_mul_result32sexlen ? {32{stage2_psimd16_mul_result_W0[31]}} : stage2_psimd16_mul_result_W1[31:0];
assign stage2_psimd16_mul_result_64b[31:0] = stage2_psimd16_mul_result_W0[31:0];
assign stage2_psimd16_mul_ovf_set = stage2_psimd16_mul_result_W0[34] | (!stage2_psimd16_mul_result32sexlen & stage2_psimd16_mul_result_W1[34]);
assign stage3_psimd16_mul_data_en = stage3_dsp_ctrl_en & stage2_dsp_ivalid & (|stage3_psimd16_mul_fctrl_nx);
assign stage3_psimd16_mul_fctrl_nx = stage2_psimd16_mul_fctrl[10:7];
assign stage3_psimd16_mul_rctrl_nx = stage2_psimd16_mul_rctrl[0];
assign stage3_psimd16_mul_out_W0_nx = stage2_psimd16_mul_result_W0[33:0];
assign stage3_psimd16_mul_out_W1_nx = stage2_psimd16_mul_result_W1[33:0];
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_psimd16_mul_fctrl <= 4'd0;
    end
    else if (stage3_dsp_ctrl_en) begin
        stage3_psimd16_mul_fctrl <= stage3_psimd16_mul_fctrl_nx;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_psimd16_mul_rctrl <= 1'b0;
        stage3_psimd16_mul_out_W0 <= 34'd0;
        stage3_psimd16_mul_out_W1 <= 34'd0;
    end
    else if (stage3_psimd16_mul_data_en) begin
        stage3_psimd16_mul_rctrl <= stage3_psimd16_mul_rctrl_nx;
        stage3_psimd16_mul_out_W0 <= stage3_psimd16_mul_out_W0_nx;
        stage3_psimd16_mul_out_W1 <= stage3_psimd16_mul_out_W1_nx;
    end
end

assign stage3_psimd16_mul_result_64b = stage3_psimd16_mul_result(stage3_psimd16_mul_fctrl, stage3_psimd16_mul_rctrl, stage3_psimd16_mul_out_W0, stage3_psimd16_mul_out_W1, {stage3_acc_din_W1,stage3_acc_din_W0});
assign stage3_psimd16_mul_ovf_set = 1'b0;
assign psimd16_result_pack_sel = function_psimd_s_pk16;
assign stage1_psimd16_result_mul_sel = function_psimd_s_mul16x16_acc32_func0 | function_psimd_s_mul16x16_out64 | function_psimd_u_mul16x16_out64;
assign stage1_psimd16_final_result_64b = ({64{psimd16_result_pack_sel}} & psimd16_pack_result_64b);
assign stage1_psimd16_final_ovf_set = (psimd16_result_pack_sel & psimd16_pack_ovf_set);
assign stage2_psimd16_result_mul_sel = (|stage2_psimd16_mul_fctrl[6:0]);
assign stage2_psimd16_final_result_64b = ({64{stage2_psimd16_result_mul_sel}} & stage2_psimd16_mul_result_64b);
assign stage2_psimd16_final_ovf_set = (stage2_psimd16_result_mul_sel & stage2_psimd16_mul_ovf_set);
assign stage3_psimd16_result_mul_sel = (|stage3_psimd16_mul_fctrl);
assign stage3_psimd16_final_result_64b = ({64{stage3_psimd16_result_mul_sel}} & stage3_psimd16_mul_result_64b);
assign stage3_psimd16_final_ovf_set = (stage3_psimd16_result_mul_sel & stage3_psimd16_mul_ovf_set);
function  [39:0] csa20_2_level;
integer i;
input [17:0] din1;
input [17:0] din2;
input [17:0] din3;
input [17:0] din4;
reg [19:0] lv1_csa1_din1;
reg [19:0] lv1_csa1_din2;
reg [19:0] lv1_csa1_din3;
reg [19:0] lv1_csa1_dout1;
reg [19:0] lv1_csa1_dout2;
reg [19:0] lv2_csa1_din1;
reg [19:0] lv2_csa1_din2;
reg [19:0] lv2_csa1_din3;
reg [19:0] lv2_csa1_dout1;
reg [19:0] lv2_csa1_dout2;
begin
    lv1_csa1_din1 = {{2{din1[17]}},din1};
    lv1_csa1_din2 = {{2{din2[17]}},din2};
    lv1_csa1_din3 = {{2{din3[17]}},din3};
    for (i = 0; i < 20; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    lv2_csa1_din1 = lv1_csa1_dout1;
    lv2_csa1_din2 = {lv1_csa1_dout2[18:0],1'b0};
    lv2_csa1_din3 = {{2{din4[17]}},din4};
    for (i = 0; i < 20; i = i + 1) begin
        {lv2_csa1_dout2[i],lv2_csa1_dout1[i]} = {1'b0,lv2_csa1_din1[i]} + {1'b0,lv2_csa1_din2[i]} + {1'b0,lv2_csa1_din3[i]};
    end
    csa20_2_level = {{lv2_csa1_dout2[18:0],1'b0},lv2_csa1_dout1[19:0]};
end
endfunction
assign function_psimd_s_mul8x8_acc32 = function_psimd_s_mul8x8_acc32_func0 | function_psimd_s_mul8x8_acc32_func1 | function_psimd_s_mul8x8_acc32_func2;
assign stage1_psimd8_mul_out_W0 = csa20_2_level(simd8_mul_out_B0, simd8_mul_out_B1, simd8_mul_out_B2, simd8_mul_out_B3);
assign stage1_psimd8_mul_out_W1 = csa20_2_level(simd8_mul_out_B4, simd8_mul_out_B5, simd8_mul_out_B6, simd8_mul_out_B7);
assign stage1_psimd8_mul_result_64b[63:48] = simd8_mul_out_B3[15:0];
assign stage1_psimd8_mul_result_64b[47:32] = simd8_mul_out_B2[15:0];
assign stage1_psimd8_mul_result_64b[31:16] = simd8_mul_out_B1[15:0];
assign stage1_psimd8_mul_result_64b[15:0] = simd8_mul_out_B0[15:0];
assign stage1_psimd8_mul_ovf_set = 1'b0;
function  [11:0] psimd8_abs_se12;
input [8:0] abs_in;
reg [8:0] adder_in1;
reg [8:0] adder_in2;
reg adder_cin;
reg [8:0] adder_out;
begin
    adder_in1 = 9'd0;
    adder_in2 = {9{abs_in[8]}} ^ abs_in;
    adder_cin = abs_in[8];
    adder_out = adder_in1 + adder_in2 + {8'd0,adder_cin};
    psimd8_abs_se12 = {{3{adder_out[8]}},adder_out};
end
endfunction
function  [23:0] csa12_2_level;
integer i;
input [11:0] din1;
input [11:0] din2;
input [11:0] din3;
input [11:0] din4;
reg [11:0] lv1_csa1_din1;
reg [11:0] lv1_csa1_din2;
reg [11:0] lv1_csa1_din3;
reg [11:0] lv1_csa1_dout1;
reg [11:0] lv1_csa1_dout2;
reg [11:0] lv2_csa1_din1;
reg [11:0] lv2_csa1_din2;
reg [11:0] lv2_csa1_din3;
reg [11:0] lv2_csa1_dout1;
reg [11:0] lv2_csa1_dout2;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 12; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    lv2_csa1_din1 = lv1_csa1_dout1;
    lv2_csa1_din2 = {lv1_csa1_dout2[10:0],1'b0};
    lv2_csa1_din3 = din4;
    for (i = 0; i < 12; i = i + 1) begin
        {lv2_csa1_dout2[i],lv2_csa1_dout1[i]} = {1'b0,lv2_csa1_din1[i]} + {1'b0,lv2_csa1_din2[i]} + {1'b0,lv2_csa1_din3[i]};
    end
    csa12_2_level = {{lv2_csa1_dout2[10:0],1'b0},lv2_csa1_dout1[11:0]};
end
endfunction
function  [31:0] csaxlen_1_level_addxlen;
integer i;
input [31:0] din1;
input [31:0] din2;
input [31:0] din3;
reg [31:0] lv1_csa1_din1;
reg [31:0] lv1_csa1_din2;
reg [31:0] lv1_csa1_din3;
reg [31:0] lv1_csa1_dout1;
reg [31:0] lv1_csa1_dout2;
reg [31:0] add_dout;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 32; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    add_dout = {lv1_csa1_dout2[30:0],1'b0} + lv1_csa1_dout1[31:0];
    csaxlen_1_level_addxlen = add_dout;
end
endfunction
assign stage1_psimd8_pbsad_out_W0 = csa12_2_level(psimd8_abs_se12(simd8_addcmp_out_B0[8:0]), psimd8_abs_se12(simd8_addcmp_out_B1[8:0]), psimd8_abs_se12(simd8_addcmp_out_B2[8:0]), psimd8_abs_se12(simd8_addcmp_out_B3[8:0]));
assign stage1_psimd8_pbsad_out_W1 = csa12_2_level(psimd8_abs_se12(simd8_addcmp_out_B4[8:0]), psimd8_abs_se12(simd8_addcmp_out_B5[8:0]), psimd8_abs_se12(simd8_addcmp_out_B6[8:0]), psimd8_abs_se12(simd8_addcmp_out_B7[8:0]));
assign stage1_psimd8_pbsad_out_64b = csa12_2_level(stage1_psimd8_pbsad_out_W0[11:0], stage1_psimd8_pbsad_out_W0[23:12], stage1_psimd8_pbsad_out_W1[11:0], stage1_psimd8_pbsad_out_W1[23:12]);
assign stage2_psimd8_pbsad_data_en = stage2_dsp_ctrl_en & stage1_dsp_ivalid & (|stage2_psimd8_pbsad_fctrl_nx);
assign stage2_psimd8_pbsad_fctrl_nx[0] = function_psimd_u_abs8_accxlen_func0;
assign stage2_psimd8_pbsad_fctrl_nx[1] = function_psimd_u_abs8_accxlen_func1;
assign stage2_psimd8_pbsad_out_nx = stage1_psimd8_pbsad_out_64b;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd8_pbsad_fctrl <= 2'd0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_psimd8_pbsad_fctrl <= stage2_psimd8_pbsad_fctrl_nx;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_psimd8_pbsad_out <= 24'd0;
    end
    else if (stage2_psimd8_pbsad_data_en) begin
        stage2_psimd8_pbsad_out <= stage2_psimd8_pbsad_out_nx;
    end
end

assign stage2_psimd8_pbsad_out_xlen = csaxlen_1_level_addxlen({{20{stage2_psimd8_pbsad_out[11]}},stage2_psimd8_pbsad_out[11:0]}, {{20{stage2_psimd8_pbsad_out[23]}},stage2_psimd8_pbsad_out[23:12]}, ({32{stage2_psimd8_pbsad_fctrl[1]}} & stage2_acc_din_64b[31:0]));
assign stage2_psimd8_pbsad_result_64b = {32'd0,stage2_psimd8_pbsad_out_xlen};
assign stage2_psimd8_pbsad_ovf_set = 1'b0;
assign stage1_psimd8_result_mul_sel = function_psimd_s_mul8x8_out64 | function_psimd_u_mul8x8_out64;
assign stage1_psimd8_final_result_64b = ({64{stage1_psimd8_result_mul_sel}} & stage1_psimd8_mul_result_64b);
assign stage1_psimd8_final_ovf_set = (stage1_psimd8_result_mul_sel & stage1_psimd8_mul_ovf_set);
assign stage2_psimd8_result_pbsad_sel = (|stage2_psimd8_pbsad_fctrl);
assign stage2_psimd8_final_result_64b = ({64{stage2_psimd8_result_pbsad_sel}} & stage2_psimd8_pbsad_result_64b);
assign stage2_psimd8_final_ovf_set = (stage2_psimd8_result_pbsad_sel & stage2_psimd8_pbsad_ovf_set);
assign profile64_op1_base_sel = operand_64p_opxlen;
assign profile64_op2_base_sel = operand_64p_opxlen;
assign profile64_op1_sxlen_sel = operand_nsimd_opxlen;
assign profile64_op2_sxlen_sel = operand_nsimd_opxlen;
assign profile64_op1_s32_sel = operand_nsimd_s_op32_sexlen;
assign profile64_op2_s32_sel = operand_nsimd_s_op32_sexlen;
assign profile64_op1_u32_sel = operand_nsimd_u_op32_sexlen;
assign profile64_op2_u32_sel = operand_nsimd_u_op32_sexlen;
assign profile64_op1_64b = ({64{profile64_op1_base_sel}} & dsp_src1_64b_pair) | ({64{profile64_op1_sxlen_sel}} & dsp_src1_64b_sxlen) | ({64{profile64_op1_s32_sel}} & {{32{dsp_data_src1[31]}},dsp_data_src1[31:0]}) | ({64{profile64_op1_u32_sel}} & {{32{1'b0}},dsp_data_src1[31:0]});
assign profile64_op2_64b = ({64{profile64_op2_base_sel}} & dsp_src2_64b_pair) | ({64{profile64_op2_sxlen_sel}} & dsp_src2_64b_sxlen) | ({64{profile64_op2_s32_sel}} & {{32{dsp_data_src2[31]}},dsp_data_src2[31:0]}) | ({64{profile64_op2_u32_sel}} & {{32{1'b0}},dsp_data_src2[31:0]});
function  [64:0] profile64_add_func;
input is_func_ave;
input se1;
input se2;
input neg1;
input neg2;
input [63:0] op1;
input [63:0] op2;
reg [64:0] adder_in1;
reg [64:0] adder_in2;
reg adder_cin;
reg [64:0] adder_out;
begin
    adder_in1 = {65{neg1}} ^ {(se1 & op1[63]),op1};
    adder_in2 = {65{neg2}} ^ {(se2 & op2[63]),op2};
    adder_cin = neg1 | neg2 | is_func_ave;
    adder_out = adder_in1 + adder_in2 + {64'd0,adder_cin};
    profile64_add_func = adder_out;
end
endfunction
function  [64:0] profile64_add_result;
input is_func_sub;
input [7:0] rctrl;
input [64:0] din;
reg [63:0] dout;
reg ovfout;
reg is_type_wrap64;
reg is_type_halve64;
reg is_type_s_sat64;
reg is_type_u_sat64;
reg is_type_s_sat32;
reg is_type_u_sat32;
reg is_type_s_sat16;
reg is_type_u_sat16;
reg wrap64_sel;
reg halve64_sel;
reg l32se64_sel;
reg l16se64_sel;
reg s_ovf64_sel;
reg s_udf64_sel;
reg u_ovf64_sel;
reg u_udf64_sel;
reg s_ovf32_sel;
reg s_udf32_sel;
reg u_ovf32_sel;
reg u_udf32_sel;
reg s_ovf16_sel;
reg s_udf16_sel;
reg u_ovf16_sel;
reg u_udf16_sel;
begin
    is_type_wrap64 = rctrl[0];
    is_type_halve64 = rctrl[1];
    is_type_s_sat64 = rctrl[2];
    is_type_u_sat64 = rctrl[3];
    is_type_s_sat32 = rctrl[4];
    is_type_u_sat32 = rctrl[5];
    is_type_s_sat16 = rctrl[6];
    is_type_u_sat16 = rctrl[7];
    halve64_sel = is_type_halve64;
    s_ovf64_sel = is_type_s_sat64 & (din[64:63] == 2'b01);
    s_udf64_sel = is_type_s_sat64 & (din[64:63] == 2'b10);
    u_ovf64_sel = is_type_u_sat64 & din[64] & !is_func_sub;
    u_udf64_sel = is_type_u_sat64 & din[64] & is_func_sub;
    s_ovf32_sel = is_type_s_sat32 & !din[64] & (din[63:31] != 33'h0_00000000);
    s_udf32_sel = is_type_s_sat32 & din[64] & (din[63:31] != 33'h1_ffffffff);
    u_ovf32_sel = is_type_u_sat32 & (is_func_sub ? (!din[64] & (|din[63:32])) : (|din[64:32]));
    u_udf32_sel = is_type_u_sat32 & din[64] & is_func_sub;
    s_ovf16_sel = is_type_s_sat16 & !din[64] & (din[63:15] != 49'h0_000000000000);
    s_udf16_sel = is_type_s_sat16 & din[64] & (din[63:15] != 49'h1_ffffffffffff);
    u_ovf16_sel = is_type_u_sat16 & (is_func_sub ? (!din[64] & (|din[63:16])) : (|din[64:16]));
    u_udf16_sel = is_type_u_sat16 & din[64] & is_func_sub;
    wrap64_sel = is_type_wrap64 | (is_type_s_sat64 & !(s_ovf64_sel | s_udf64_sel)) | (is_type_u_sat64 & !(u_ovf64_sel | u_udf64_sel));
    l32se64_sel = (is_type_s_sat32 & !(s_ovf32_sel | s_udf32_sel)) | (is_type_u_sat32 & !(u_ovf32_sel | u_udf32_sel));
    l16se64_sel = (is_type_s_sat16 & !(s_ovf16_sel | s_udf16_sel)) | (is_type_u_sat16 & !(u_ovf16_sel | u_udf16_sel));
    dout = ({64{wrap64_sel}} & din[63:0]) | ({64{halve64_sel}} & din[64:1]) | ({64{l32se64_sel}} & {{32{din[31]}},din[31:0]}) | ({64{l16se64_sel}} & {{48{din[15]}},din[15:0]}) | ({64{s_ovf64_sel}} & 64'h7fffffffffffffff) | ({64{s_udf64_sel}} & 64'h8000000000000000) | ({64{u_ovf64_sel}} & 64'hffffffffffffffff) | ({64{u_udf64_sel}} & 64'h0000000000000000) | ({64{s_ovf32_sel}} & 64'h000000007fffffff) | ({64{s_udf32_sel}} & 64'hffffffff80000000) | ({64{u_ovf32_sel}} & 64'hffffffffffffffff) | ({64{u_udf32_sel}} & 64'h0000000000000000) | ({64{s_ovf16_sel}} & 64'h0000000000007fff) | ({64{s_udf16_sel}} & 64'hffffffffffff8000) | ({64{u_ovf16_sel}} & 64'hffffffffffffffff) | ({64{u_udf16_sel}} & 64'h0000000000000000);
    ovfout = s_ovf64_sel | s_udf64_sel | u_ovf64_sel | u_udf64_sel | s_ovf32_sel | s_udf32_sel | u_ovf32_sel | u_udf32_sel | s_ovf16_sel | s_udf16_sel | u_ovf16_sel | u_udf16_sel;
    profile64_add_result = {ovfout,dout};
end
endfunction
assign profile64_add_se1_64b = function_64p_s_add64 | function_64p_s_sub64 | function_nsimd_s_addxlen | function_nsimd_s_subxlen | function_nsimd_s_avexlen;
assign profile64_add_se2_64b = function_64p_s_add64 | function_64p_s_sub64 | function_nsimd_s_addxlen | function_nsimd_s_subxlen | function_nsimd_s_avexlen;
assign profile64_add_neg1_64b = 1'b0;
assign profile64_add_neg2_64b = function_64p_s_sub64 | function_64p_u_sub64 | function_nsimd_s_subxlen | function_nsimd_u_subxlen;
assign profile64_add_out_64b = profile64_add_func(function_nsimd_s_avexlen, profile64_add_se1_64b, profile64_add_se2_64b, profile64_add_neg1_64b, profile64_add_neg2_64b, profile64_op1_64b, profile64_op2_64b);
assign profile64_add_rctrl[0] = result_64p_s_wrap64;
assign profile64_add_rctrl[1] = result_64p_s_halve64 | result_64p_u_halve64 | result_nsimd_s_halvexlen;
assign profile64_add_rctrl[2] = result_64p_s_sat64;
assign profile64_add_rctrl[3] = result_64p_u_sat64;
assign profile64_add_rctrl[4] = result_nsimd_s_sat32_sexlen;
assign profile64_add_rctrl[5] = result_nsimd_u_sat32_sexlen;
assign profile64_add_rctrl[6] = result_nsimd_s_sat16_sexlen;
assign profile64_add_rctrl[7] = result_nsimd_u_sat16_sexlen;
assign {profile64_add_ovf_set,profile64_add_result_64b} = profile64_add_result(profile64_add_neg2_64b, profile64_add_rctrl, profile64_add_out_64b);
function  [133:0] csa67_1_level;
integer i;
input [66:0] din1;
input [66:0] din2;
input [66:0] din3;
reg [66:0] lv1_csa1_din1;
reg [66:0] lv1_csa1_din2;
reg [66:0] lv1_csa1_din3;
reg [66:0] lv1_csa1_dout1;
reg [66:0] lv1_csa1_dout2;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 67; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    csa67_1_level = {{lv1_csa1_dout2[65:0],1'b0},lv1_csa1_dout1[66:0]};
end
endfunction
function  [133:0] csa67_2_level;
integer i;
input [66:0] din1;
input [66:0] din2;
input [66:0] din3;
input [66:0] din4;
reg [66:0] lv1_csa1_din1;
reg [66:0] lv1_csa1_din2;
reg [66:0] lv1_csa1_din3;
reg [66:0] lv1_csa1_dout1;
reg [66:0] lv1_csa1_dout2;
reg [66:0] lv2_csa1_din1;
reg [66:0] lv2_csa1_din2;
reg [66:0] lv2_csa1_din3;
reg [66:0] lv2_csa1_dout1;
reg [66:0] lv2_csa1_dout2;
begin
    lv1_csa1_din1 = din1;
    lv1_csa1_din2 = din2;
    lv1_csa1_din3 = din3;
    for (i = 0; i < 67; i = i + 1) begin
        {lv1_csa1_dout2[i],lv1_csa1_dout1[i]} = {1'b0,lv1_csa1_din1[i]} + {1'b0,lv1_csa1_din2[i]} + {1'b0,lv1_csa1_din3[i]};
    end
    lv2_csa1_din1 = lv1_csa1_dout1;
    lv2_csa1_din2 = {lv1_csa1_dout2[65:0],1'b0};
    lv2_csa1_din3 = din4;
    for (i = 0; i < 67; i = i + 1) begin
        {lv2_csa1_dout2[i],lv2_csa1_dout1[i]} = {1'b0,lv2_csa1_din1[i]} + {1'b0,lv2_csa1_din2[i]} + {1'b0,lv2_csa1_din3[i]};
    end
    csa67_2_level = {{lv2_csa1_dout2[65:0],1'b0},lv2_csa1_dout1[66:0]};
end
endfunction
function  [133:0] stage2_mul32x32_acc64_out;
input [5:0] fctrl;
input [133:0] mul_din1;
input [133:0] mul_din2;
input [63:0] acc_din;
input acc_sign;
reg is_func_kmda;
reg is_func_smds;
reg is_func_kma;
reg is_func_kmada;
reg is_func_kmads;
reg is_func_kmsda;
reg acc_din1_en;
reg acc_din2_en;
reg acc_din3_en;
reg acc_din2_sub;
reg acc_din3_sub;
reg [66:0] acc_din1;
reg [66:0] acc_din2;
reg [66:0] acc_din3;
reg [66:0] acc_din4;
reg [66:0] acc_din5;
reg [66:0] acc_din6;
reg [66:0] acc_pp1;
reg [66:0] acc_pp2;
reg [66:0] acc_pp3;
reg [66:0] acc_pp4;
reg [66:0] acc_dout1;
reg [66:0] acc_dout2;
begin
    is_func_kmda = fctrl[0];
    is_func_smds = fctrl[1];
    is_func_kma = fctrl[2];
    is_func_kmada = fctrl[3];
    is_func_kmads = fctrl[4];
    is_func_kmsda = fctrl[5];
    acc_din1_en = is_func_kma | is_func_kmada | is_func_kmads | is_func_kmsda;
    acc_din2_en = is_func_kmda | is_func_smds | is_func_kmada | is_func_kmads | is_func_kmsda;
    acc_din3_en = is_func_kmda | is_func_smds | is_func_kma | is_func_kmada | is_func_kmads | is_func_kmsda;
    acc_din2_sub = is_func_kmsda;
    acc_din3_sub = is_func_smds | is_func_kmads | is_func_kmsda;
    acc_din1 = {67{acc_din1_en}} & {{3{(acc_sign & acc_din[63])}},acc_din[63:0]};
    acc_din4[66:0] = {64'd0,({1'b0,acc_din2_sub} + {1'b0,acc_din3_sub}),1'b0};
    acc_din2 = {67{acc_din2_sub}} ^ {67{acc_din2_en}} & {mul_din1[66:0]};
    acc_din3 = {67{acc_din3_sub}} ^ {67{acc_din3_en}} & {mul_din2[66:0]};
    acc_din5 = {67{acc_din2_sub}} ^ {67{acc_din2_en}} & {mul_din1[133:67]};
    acc_din6 = {67{acc_din3_sub}} ^ {67{acc_din3_en}} & {mul_din2[133:67]};
    {acc_pp2,acc_pp1} = csa67_1_level(acc_din1, acc_din2, acc_din3);
    {acc_pp4,acc_pp3} = csa67_1_level(acc_din4, acc_din5, acc_din6);
    {acc_dout2,acc_dout1} = csa67_2_level(acc_pp1, acc_pp2, acc_pp3, acc_pp4);
    stage2_mul32x32_acc64_out = {acc_dout2,acc_dout1};
end
endfunction
function  [64:0] stage3_mul32x32_acc64_out;
input is_func_sub;
input is_type_s_sat;
input is_type_u_sat;
input [66:0] din1;
input [66:0] din2;
reg [66:0] adder_out;
reg [63:0] dout;
reg ovfout;
reg wrap_sel;
reg s_ovf_sel;
reg s_udf_sel;
reg u_ovf_sel;
reg u_udf_sel;
begin
    adder_out = din1 + din2;
    s_ovf_sel = is_type_s_sat & !adder_out[66] & (adder_out[65:63] != 3'b000);
    s_udf_sel = is_type_s_sat & adder_out[66] & (adder_out[65:63] != 3'b111);
    u_ovf_sel = is_type_u_sat & (is_func_sub ? (!adder_out[66] & (|adder_out[65:64])) : (|adder_out[66:64]));
    u_udf_sel = is_type_u_sat & adder_out[66] & is_func_sub;
    wrap_sel = (!is_type_s_sat & !is_type_u_sat) | (is_type_s_sat & !(s_ovf_sel | s_udf_sel)) | (is_type_u_sat & !(u_ovf_sel | u_udf_sel));
    dout = ({64{wrap_sel}} & adder_out[63:0]) | ({64{s_ovf_sel}} & 64'h7fffffffffffffff) | ({64{s_udf_sel}} & 64'h8000000000000000) | ({64{u_ovf_sel}} & 64'hffffffffffffffff) | ({64{u_udf_sel}} & 64'h0000000000000000);
    ovfout = s_ovf_sel | s_udf_sel | u_ovf_sel | u_udf_sel;
    stage3_mul32x32_acc64_out = {ovfout,dout};
end
endfunction
assign {stage2_profile64_mul_csa_out2,stage2_profile64_mul_csa_out1} = stage2_mul32x32_acc64_out(stage2_psimd32_mul_fctrl[16:11], stage2_psimd32_mul_lv1_result_W1[175:42], stage2_psimd32_mul_lv1_result_W0[175:42], stage2_acc_din_64b, stage2_acc_din_sign);
assign stage3_profile64_msr64 = stage3_psimd32_mul_fctrl[5];
assign stage3_profile64_s_sat64 = stage3_psimd32_mul_rctrl[0];
assign stage3_profile64_u_sat64 = stage3_psimd32_mul_rctrl[1];
assign {stage3_profile64_mul_ovf_set,stage3_profile64_mul_result_64b} = stage3_mul32x32_acc64_out(stage3_profile64_msr64, stage3_profile64_s_sat64, stage3_profile64_u_sat64, stage3_psimd32_mul_out1, stage3_psimd32_mul_out2);
assign profile64_result_add_sel = function_64p_s_add64 | function_64p_u_add64 | function_64p_s_sub64 | function_64p_u_sub64 | function_nsimd_s_addxlen | function_nsimd_u_addxlen | function_nsimd_s_subxlen | function_nsimd_u_subxlen | function_nsimd_s_avexlen;
assign stage1_profile64_final_result_64b = ({64{profile64_result_add_sel}} & profile64_add_result_64b);
assign stage1_profile64_final_ovf_set = (profile64_result_add_sel & profile64_add_ovf_set);
function  [32:0] nsimd16_mul_result;
input is_type_s_sat16;
input is_type_s_sat32;
input [15:0] op1;
input [15:0] op2;
input [31:0] din;
reg [31:0] dout;
reg ovfout;
reg s_ovf16_sel;
reg s_ovf32_sel;
reg sra15_sel;
reg sll1_sel;
begin
    s_ovf16_sel = is_type_s_sat16 & (op1 == 16'h8000) & (op2 == 16'h8000);
    sra15_sel = is_type_s_sat16 & !s_ovf16_sel;
    s_ovf32_sel = is_type_s_sat32 & (op1 == 16'h8000) & (op2 == 16'h8000);
    sll1_sel = is_type_s_sat32 & !s_ovf32_sel;
    dout = ({32{sra15_sel}} & {{16{din[30]}},din[30:15]}) | ({32{s_ovf16_sel}} & 32'h00007fff) | ({32{sll1_sel}} & {din[30:0],1'b0}) | ({32{s_ovf32_sel}} & 32'h7fffffff);
    ovfout = s_ovf16_sel | s_ovf32_sel;
    nsimd16_mul_result = {ovfout,dout};
end
endfunction
assign nsimd16_mul_s_sat16 = result_nsimd_s_sat16_sexlen | result_nsimd_s_sat16_se32;
assign nsimd16_mul_s_sat32 = result_nsimd_s_sat32_sexlen | result_nsimd_s_sat32;
assign nsimd16_mul_result_H0 = nsimd16_mul_result(nsimd16_mul_s_sat16, nsimd16_mul_s_sat32, simd16_op1_H0, simd16_op2_H0, simd16_mul_out_H0);
assign nsimd16_mul_result_H2 = nsimd16_mul_result(nsimd16_mul_s_sat16, nsimd16_mul_s_sat32, simd16_op1_H2, simd16_op2_H2, simd16_mul_out_H2);
assign nsimd16_mul_resultsexlen = result_nsimd_s_sat16_sexlen | result_nsimd_s_sat32_sexlen;
assign stage1_nsimd16_mul_result_64b[63:32] = nsimd16_mul_resultsexlen ? {32{nsimd16_mul_result_H0[31]}} : nsimd16_mul_result_H2[31:0];
assign stage1_nsimd16_mul_result_64b[31:0] = nsimd16_mul_result_H0[31:0];
assign stage1_nsimd16_mul_ovf_set = nsimd16_mul_result_H0[32] | (!nsimd16_mul_resultsexlen & nsimd16_mul_result_H2[32]);
assign stage1_nsimd16_result_mul_sel = function_nsimd_s_mul16x16 | function_nsimd_s_mul16x16_double32;
assign stage1_nsimd16_final_result_64b = 64'd0;
assign stage1_nsimd16_final_ovf_set = 1'b0;
assign stage1_xsimd16_result_mul_sel = simd16_result_mul_sel | stage1_psimd16_result_mul_sel | stage1_nsimd16_result_mul_sel;
assign stage1_xsimd16_mul_result_64b = ({64{simd16_result_mul_sel}} & simd16_mul_result_64b) | ({64{stage1_psimd16_result_mul_sel}} & stage1_psimd16_mul_result_64b) | ({64{stage1_nsimd16_result_mul_sel}} & stage1_nsimd16_mul_result_64b);
assign stage1_xsimd16_mul_ovf_set = (simd16_result_mul_sel & simd16_mul_ovf_set) | (stage1_psimd16_result_mul_sel & stage1_psimd16_mul_ovf_set) | (stage1_nsimd16_result_mul_sel & stage1_nsimd16_mul_ovf_set);
assign stage2_xsimd16_mul_data_en = stage2_dsp_ctrl_en & stage1_dsp_ivalid & stage1_xsimd16_result_mul_sel;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_xsimd16_result_mul_sel <= 1'b0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_xsimd16_result_mul_sel <= stage1_xsimd16_result_mul_sel;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_xsimd16_mul_result_64b <= 64'd0;
        stage2_xsimd16_mul_ovf_set <= 1'b0;
    end
    else if (stage2_xsimd16_mul_data_en) begin
        stage2_xsimd16_mul_result_64b <= stage1_xsimd16_mul_result_64b;
        stage2_xsimd16_mul_ovf_set <= stage1_xsimd16_mul_ovf_set;
    end
end

assign stage2_xsimd16_final_result_64b = ({64{stage2_xsimd16_result_mul_sel}} & stage2_xsimd16_mul_result_64b);
assign stage2_xsimd16_final_ovf_set = (stage2_xsimd16_result_mul_sel & stage2_xsimd16_mul_ovf_set);
assign dsp_stage1_result = stage1_simd16_final_result_64b | stage1_simd8_final_result_64b | stage1_psimd32_final_result_64b | stage1_psimdxlen_final_result_64b | stage1_psimd16_final_result_64b | stage1_psimd8_final_result_64b | stage1_profile64_final_result_64b | stage1_nsimd16_final_result_64b;
assign dsp_stage1_ovf_set = stage1_dsp_ovfset & (stage1_simd16_final_ovf_set | stage1_simd8_final_ovf_set | stage1_psimd32_final_ovf_set | stage1_psimdxlen_final_ovf_set | stage1_psimd16_final_ovf_set | stage1_psimd8_final_ovf_set | stage1_profile64_final_ovf_set | stage1_nsimd16_final_ovf_set);
assign dsp_stage2_result = stage2_psimd32_final_result_64b | stage2_psimd16_final_result_64b | stage2_xsimd16_final_result_64b | stage2_psimd8_final_result_64b;
assign dsp_stage2_ovf_set = stage2_dsp_ovfset & (stage2_psimd32_final_ovf_set | stage2_psimd16_final_ovf_set | stage2_xsimd16_final_ovf_set | stage2_psimd8_final_ovf_set);
assign dsp_stage3_result = stage3_psimd32_final_result_64b | stage3_psimd16_final_result_64b;
assign dsp_stage3_ovf_set = stage3_dsp_ovfset & (stage3_psimd32_final_ovf_set | stage3_psimd16_final_ovf_set);
assign stage2_dsp_ctrl_en = dsp_stage2_pipe_en;
assign stage3_dsp_ctrl_en = dsp_stage3_pipe_en;
assign stage1_dsp_ivalid = dsp_instr_valid;
assign stage1_dsp_ovfset = dsp_overflow_ctrl;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_dsp_ivalid <= 1'b0;
        stage2_dsp_ovfset <= 1'b0;
    end
    else if (stage2_dsp_ctrl_en) begin
        stage2_dsp_ivalid <= stage1_dsp_ivalid;
        stage2_dsp_ovfset <= stage1_dsp_ovfset;
    end
end

always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_dsp_ovfset <= 1'b0;
    end
    else if (stage3_dsp_ctrl_en) begin
        stage3_dsp_ovfset <= stage2_dsp_ovfset;
    end
end

assign acc_din_smal_sel = operand_psimd_smal_op16;
assign acc_din_base_sel = !acc_din_smal_sel;
assign stage1_acc_din_W0 = ({32{acc_din_base_sel}} & dsp_src3_64b_pair[31:0]) | ({32{acc_din_smal_sel}} & dsp_src1_64b_pair[31:0]);
assign stage1_acc_din_W1 = ({32{acc_din_base_sel}} & dsp_src3_64b_pair[63:32]) | ({32{acc_din_smal_sel}} & dsp_src1_64b_pair[63:32]);
assign stage2_acc_din_en = stage2_dsp_ctrl_en & stage1_dsp_ivalid & (|{stage2_psimd32_mul_fctrl_nx,stage2_psimd16_mul_fctrl_nx,stage2_psimd8_pbsad_fctrl_nx});
assign stage2_acc_din_W0_nx = stage1_acc_din_W0;
assign stage2_acc_din_W1_nx = stage1_acc_din_W1;
assign stage2_acc_din_sign_nx = !(function_64p_u_mul32x32_acc64_func0 | function_64p_u_mul32x32_acc64_func1 | function_psimd_s_mul8x8_acc32_func1);
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage2_acc_din_W0 <= 32'd0;
        stage2_acc_din_W1 <= 32'd0;
        stage2_acc_din_sign <= 1'b0;
    end
    else if (stage2_acc_din_en) begin
        stage2_acc_din_W0 <= stage2_acc_din_W0_nx;
        stage2_acc_din_W1 <= stage2_acc_din_W1_nx;
        stage2_acc_din_sign <= stage2_acc_din_sign_nx;
    end
end

assign stage2_acc_din_64b = {stage2_acc_din_W1,stage2_acc_din_W0};
assign stage3_acc_din_en = stage3_dsp_ctrl_en & stage2_dsp_ivalid & (|stage3_psimd16_mul_fctrl_nx);
assign stage3_acc_din_W0_nx = stage2_acc_din_W0;
assign stage3_acc_din_W1_nx = stage2_acc_din_W1;
always @(posedge core_clk or negedge core_reset_n) begin
    if (!core_reset_n) begin
        stage3_acc_din_W0 <= 32'd0;
        stage3_acc_din_W1 <= 32'd0;
    end
    else if (stage3_acc_din_en) begin
        stage3_acc_din_W0 <= stage3_acc_din_W0_nx;
        stage3_acc_din_W1 <= stage3_acc_din_W1_nx;
    end
end

endmodule

