-------------------------------------------------------------------------------
--
-- SD/MMC Bootloader
--
-- $Id: card-c.vhd,v 1.1 2005-02-08 21:09:18 arniml Exp $
--
-------------------------------------------------------------------------------

configuration card_behav_c0 of card is

  for behav
  end for;

end card_behav_c0;
