// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_dsp_mul32 (
    mul_op1,
    mul_op2,
    mul_op1_sign,
    mul_op2_sign,
    mul_wt_sum,
    mul_wt_cout
);
parameter INLEN = 32;
parameter OUTLEN = 67;
localparam PPLEN = OUTLEN;
input [INLEN - 1:0] mul_op1;
input [INLEN - 1:0] mul_op2;
input mul_op1_sign;
input mul_op2_sign;
output [OUTLEN - 1:0] mul_wt_sum;
output [OUTLEN - 1:0] mul_wt_cout;


wire [INLEN:0] s0;
wire [INLEN:0] s1;
wire s2;
wire [PPLEN - 1:0] s3;
wire [PPLEN - 1:0] s4;
wire [PPLEN - 1:1] s5;
wire [PPLEN - 1:2] s6;
wire [PPLEN - 1:3] s7;
wire [PPLEN - 1:4] s8;
wire [PPLEN - 1:5] s9;
wire [PPLEN - 1:6] s10;
wire [PPLEN - 1:7] s11;
wire [PPLEN - 1:8] s12;
wire [PPLEN - 1:9] s13;
wire [PPLEN - 1:10] s14;
wire [PPLEN - 1:11] s15;
wire [PPLEN - 1:12] s16;
wire [PPLEN - 1:13] s17;
wire [PPLEN - 1:14] s18;
wire [PPLEN - 1:15] s19;
wire [PPLEN - 1:16] s20;
wire [PPLEN - 1:17] s21;
wire [PPLEN - 1:18] s22;
wire [PPLEN - 1:19] s23;
wire [PPLEN - 1:20] s24;
wire [PPLEN - 1:21] s25;
wire [PPLEN - 1:22] s26;
wire [PPLEN - 1:23] s27;
wire [PPLEN - 1:24] s28;
wire [PPLEN - 1:25] s29;
wire [PPLEN - 1:26] s30;
wire [PPLEN - 1:27] s31;
wire [PPLEN - 1:28] s32;
wire [PPLEN - 1:29] s33;
wire [PPLEN - 1:30] s34;
wire [PPLEN - 1:31] s35;
wire [PPLEN - 1:32] s36;
wire [PPLEN - 1:32] s37;
wire [PPLEN - 1:0] s38;
wire [PPLEN:1] s39;
wire [PPLEN - 1:3] s40;
wire [PPLEN:4] s41;
wire [PPLEN - 1:6] s42;
wire [PPLEN:7] s43;
wire [PPLEN - 1:9] s44;
wire [PPLEN:10] s45;
wire [PPLEN - 1:12] s46;
wire [PPLEN:13] s47;
wire [PPLEN - 1:15] s48;
wire [PPLEN:16] s49;
wire [PPLEN - 1:18] s50;
wire [PPLEN:19] s51;
wire [PPLEN - 1:21] s52;
wire [PPLEN:22] s53;
wire [PPLEN - 1:24] s54;
wire [PPLEN:25] s55;
wire [PPLEN - 1:27] s56;
wire [PPLEN:28] s57;
wire [PPLEN - 1:30] s58;
wire [PPLEN:31] s59;
wire [PPLEN - 1:32] s60;
wire [PPLEN - 1:0] s61;
wire [PPLEN:1] s62;
wire [PPLEN - 1:4] s63;
wire [PPLEN:5] s64;
wire [PPLEN - 1:9] s65;
wire [PPLEN:10] s66;
wire [PPLEN - 1:13] s67;
wire [PPLEN:14] s68;
wire [PPLEN - 1:18] s69;
wire [PPLEN:19] s70;
wire [PPLEN - 1:22] s71;
wire [PPLEN:23] s72;
wire [PPLEN - 1:27] s73;
wire [PPLEN:28] s74;
wire [PPLEN - 1:31] s75;
wire [PPLEN - 1:32] s76;
wire [PPLEN - 1:0] s77;
wire [PPLEN:1] s78;
wire [PPLEN - 1:5] s79;
wire [PPLEN:6] s80;
wire [PPLEN - 1:13] s81;
wire [PPLEN:14] s82;
wire [PPLEN - 1:19] s83;
wire [PPLEN:20] s84;
wire [PPLEN - 1:27] s85;
wire [PPLEN:28] s86;
wire [PPLEN - 1:32] s87;
wire [PPLEN - 1:0] s88;
wire [PPLEN:1] s89;
wire [PPLEN - 1:6] s90;
wire [PPLEN:7] s91;
wire [PPLEN - 1:19] s92;
wire [PPLEN:20] s93;
wire [PPLEN - 1:28] s94;
wire [PPLEN - 1:32] s95;
wire [PPLEN - 1:0] s96;
wire [PPLEN:1] s97;
wire [PPLEN - 1:7] s98;
wire [PPLEN:8] s99;
wire [PPLEN - 1:28] s100;
wire [PPLEN - 1:32] s101;
wire [PPLEN - 1:0] s102;
wire [PPLEN:1] s103;
wire [PPLEN - 1:8] s104;
wire [PPLEN:9] s105;
wire [PPLEN - 1:0] s106;
wire [PPLEN:1] s107;
wire [PPLEN - 1:9] s108;
wire [PPLEN - 1:0] s109;
wire [PPLEN:1] s110;
assign s0 = {(mul_op1_sign & mul_op1[INLEN - 1]),mul_op1};
assign s1 = {(mul_op2_sign & mul_op2[INLEN - 1]),mul_op2};
assign s2 = mul_op2_sign & s1[INLEN];
assign s3 = {{(PPLEN - INLEN - 1){s0[INLEN]}},s0};
assign s4 = (s3[PPLEN - 1:0] & {(PPLEN - 0){s1[0]}});
assign s5 = (s3[PPLEN - 2:0] & {(PPLEN - 1){s1[1]}});
assign s6 = (s3[PPLEN - 3:0] & {(PPLEN - 2){s1[2]}});
assign s7 = (s3[PPLEN - 4:0] & {(PPLEN - 3){s1[3]}});
assign s8 = (s3[PPLEN - 5:0] & {(PPLEN - 4){s1[4]}});
assign s9 = (s3[PPLEN - 6:0] & {(PPLEN - 5){s1[5]}});
assign s10 = (s3[PPLEN - 7:0] & {(PPLEN - 6){s1[6]}});
assign s11 = (s3[PPLEN - 8:0] & {(PPLEN - 7){s1[7]}});
assign s12 = (s3[PPLEN - 9:0] & {(PPLEN - 8){s1[8]}});
assign s13 = (s3[PPLEN - 10:0] & {(PPLEN - 9){s1[9]}});
assign s14 = (s3[PPLEN - 11:0] & {(PPLEN - 10){s1[10]}});
assign s15 = (s3[PPLEN - 12:0] & {(PPLEN - 11){s1[11]}});
assign s16 = (s3[PPLEN - 13:0] & {(PPLEN - 12){s1[12]}});
assign s17 = (s3[PPLEN - 14:0] & {(PPLEN - 13){s1[13]}});
assign s18 = (s3[PPLEN - 15:0] & {(PPLEN - 14){s1[14]}});
assign s19 = (s3[PPLEN - 16:0] & {(PPLEN - 15){s1[15]}});
assign s20 = (s3[PPLEN - 17:0] & {(PPLEN - 16){s1[16]}});
assign s21 = (s3[PPLEN - 18:0] & {(PPLEN - 17){s1[17]}});
assign s22 = (s3[PPLEN - 19:0] & {(PPLEN - 18){s1[18]}});
assign s23 = (s3[PPLEN - 20:0] & {(PPLEN - 19){s1[19]}});
assign s24 = (s3[PPLEN - 21:0] & {(PPLEN - 20){s1[20]}});
assign s25 = (s3[PPLEN - 22:0] & {(PPLEN - 21){s1[21]}});
assign s26 = (s3[PPLEN - 23:0] & {(PPLEN - 22){s1[22]}});
assign s27 = (s3[PPLEN - 24:0] & {(PPLEN - 23){s1[23]}});
assign s28 = (s3[PPLEN - 25:0] & {(PPLEN - 24){s1[24]}});
assign s29 = (s3[PPLEN - 26:0] & {(PPLEN - 25){s1[25]}});
assign s30 = (s3[PPLEN - 27:0] & {(PPLEN - 26){s1[26]}});
assign s31 = (s3[PPLEN - 28:0] & {(PPLEN - 27){s1[27]}});
assign s32 = (s3[PPLEN - 29:0] & {(PPLEN - 28){s1[28]}});
assign s33 = (s3[PPLEN - 30:0] & {(PPLEN - 29){s1[29]}});
assign s34 = (s3[PPLEN - 31:0] & {(PPLEN - 30){s1[30]}});
assign s35 = (s3[PPLEN - 32:0] & {(PPLEN - 31){s1[31]}});
assign s36 = {(PPLEN - 32){s2}} ^ (s3[PPLEN - 33:0] & {(PPLEN - 32){s1[32]}});
assign s37 = {{(PPLEN - 33){1'b0}},s2};
assign {s39[1],s38[0]} = {1'b0,s4[0]};
assign {s39[2],s38[1]} = {1'b0,s5[1]} + {1'b0,s4[1]};
assign {s39[3],s38[2]} = {1'b0,s6[2]} + {1'b0,s5[2]} + {1'b0,s4[2]};
assign {s39[4],s38[3]} = {1'b0,s6[3]} + {1'b0,s5[3]} + {1'b0,s4[3]};
assign {s39[5],s38[4]} = {1'b0,s6[4]} + {1'b0,s5[4]} + {1'b0,s4[4]};
assign {s39[6],s38[5]} = {1'b0,s6[5]} + {1'b0,s5[5]} + {1'b0,s4[5]};
assign {s39[7],s38[6]} = {1'b0,s6[6]} + {1'b0,s5[6]} + {1'b0,s4[6]};
assign {s39[8],s38[7]} = {1'b0,s6[7]} + {1'b0,s5[7]} + {1'b0,s4[7]};
assign {s39[9],s38[8]} = {1'b0,s6[8]} + {1'b0,s5[8]} + {1'b0,s4[8]};
assign {s39[10],s38[9]} = {1'b0,s6[9]} + {1'b0,s5[9]} + {1'b0,s4[9]};
assign {s39[11],s38[10]} = {1'b0,s6[10]} + {1'b0,s5[10]} + {1'b0,s4[10]};
assign {s39[12],s38[11]} = {1'b0,s6[11]} + {1'b0,s5[11]} + {1'b0,s4[11]};
assign {s39[13],s38[12]} = {1'b0,s6[12]} + {1'b0,s5[12]} + {1'b0,s4[12]};
assign {s39[14],s38[13]} = {1'b0,s6[13]} + {1'b0,s5[13]} + {1'b0,s4[13]};
assign {s39[15],s38[14]} = {1'b0,s6[14]} + {1'b0,s5[14]} + {1'b0,s4[14]};
assign {s39[16],s38[15]} = {1'b0,s6[15]} + {1'b0,s5[15]} + {1'b0,s4[15]};
assign {s39[17],s38[16]} = {1'b0,s6[16]} + {1'b0,s5[16]} + {1'b0,s4[16]};
assign {s39[18],s38[17]} = {1'b0,s6[17]} + {1'b0,s5[17]} + {1'b0,s4[17]};
assign {s39[19],s38[18]} = {1'b0,s6[18]} + {1'b0,s5[18]} + {1'b0,s4[18]};
assign {s39[20],s38[19]} = {1'b0,s6[19]} + {1'b0,s5[19]} + {1'b0,s4[19]};
assign {s39[21],s38[20]} = {1'b0,s6[20]} + {1'b0,s5[20]} + {1'b0,s4[20]};
assign {s39[22],s38[21]} = {1'b0,s6[21]} + {1'b0,s5[21]} + {1'b0,s4[21]};
assign {s39[23],s38[22]} = {1'b0,s6[22]} + {1'b0,s5[22]} + {1'b0,s4[22]};
assign {s39[24],s38[23]} = {1'b0,s6[23]} + {1'b0,s5[23]} + {1'b0,s4[23]};
assign {s39[25],s38[24]} = {1'b0,s6[24]} + {1'b0,s5[24]} + {1'b0,s4[24]};
assign {s39[26],s38[25]} = {1'b0,s6[25]} + {1'b0,s5[25]} + {1'b0,s4[25]};
assign {s39[27],s38[26]} = {1'b0,s6[26]} + {1'b0,s5[26]} + {1'b0,s4[26]};
assign {s39[28],s38[27]} = {1'b0,s6[27]} + {1'b0,s5[27]} + {1'b0,s4[27]};
assign {s39[29],s38[28]} = {1'b0,s6[28]} + {1'b0,s5[28]} + {1'b0,s4[28]};
assign {s39[30],s38[29]} = {1'b0,s6[29]} + {1'b0,s5[29]} + {1'b0,s4[29]};
assign {s39[31],s38[30]} = {1'b0,s6[30]} + {1'b0,s5[30]} + {1'b0,s4[30]};
assign {s39[32],s38[31]} = {1'b0,s6[31]} + {1'b0,s5[31]} + {1'b0,s4[31]};
assign {s39[33],s38[32]} = {1'b0,s6[32]} + {1'b0,s5[32]} + {1'b0,s4[32]};
assign {s39[34],s38[33]} = {1'b0,s6[33]} + {1'b0,s5[33]} + {1'b0,s4[33]};
assign {s39[35],s38[34]} = {1'b0,s6[34]} + {1'b0,s5[34]} + {1'b0,s4[34]};
assign {s39[36],s38[35]} = {1'b0,s6[35]} + {1'b0,s5[35]} + {1'b0,s4[35]};
assign {s39[37],s38[36]} = {1'b0,s6[36]} + {1'b0,s5[36]} + {1'b0,s4[36]};
assign {s39[38],s38[37]} = {1'b0,s6[37]} + {1'b0,s5[37]} + {1'b0,s4[37]};
assign {s39[39],s38[38]} = {1'b0,s6[38]} + {1'b0,s5[38]} + {1'b0,s4[38]};
assign {s39[40],s38[39]} = {1'b0,s6[39]} + {1'b0,s5[39]} + {1'b0,s4[39]};
assign {s39[41],s38[40]} = {1'b0,s6[40]} + {1'b0,s5[40]} + {1'b0,s4[40]};
assign {s39[42],s38[41]} = {1'b0,s6[41]} + {1'b0,s5[41]} + {1'b0,s4[41]};
assign {s39[43],s38[42]} = {1'b0,s6[42]} + {1'b0,s5[42]} + {1'b0,s4[42]};
assign {s39[44],s38[43]} = {1'b0,s6[43]} + {1'b0,s5[43]} + {1'b0,s4[43]};
assign {s39[45],s38[44]} = {1'b0,s6[44]} + {1'b0,s5[44]} + {1'b0,s4[44]};
assign {s39[46],s38[45]} = {1'b0,s6[45]} + {1'b0,s5[45]} + {1'b0,s4[45]};
assign {s39[47],s38[46]} = {1'b0,s6[46]} + {1'b0,s5[46]} + {1'b0,s4[46]};
assign {s39[48],s38[47]} = {1'b0,s6[47]} + {1'b0,s5[47]} + {1'b0,s4[47]};
assign {s39[49],s38[48]} = {1'b0,s6[48]} + {1'b0,s5[48]} + {1'b0,s4[48]};
assign {s39[50],s38[49]} = {1'b0,s6[49]} + {1'b0,s5[49]} + {1'b0,s4[49]};
assign {s39[51],s38[50]} = {1'b0,s6[50]} + {1'b0,s5[50]} + {1'b0,s4[50]};
assign {s39[52],s38[51]} = {1'b0,s6[51]} + {1'b0,s5[51]} + {1'b0,s4[51]};
assign {s39[53],s38[52]} = {1'b0,s6[52]} + {1'b0,s5[52]} + {1'b0,s4[52]};
assign {s39[54],s38[53]} = {1'b0,s6[53]} + {1'b0,s5[53]} + {1'b0,s4[53]};
assign {s39[55],s38[54]} = {1'b0,s6[54]} + {1'b0,s5[54]} + {1'b0,s4[54]};
assign {s39[56],s38[55]} = {1'b0,s6[55]} + {1'b0,s5[55]} + {1'b0,s4[55]};
assign {s39[57],s38[56]} = {1'b0,s6[56]} + {1'b0,s5[56]} + {1'b0,s4[56]};
assign {s39[58],s38[57]} = {1'b0,s6[57]} + {1'b0,s5[57]} + {1'b0,s4[57]};
assign {s39[59],s38[58]} = {1'b0,s6[58]} + {1'b0,s5[58]} + {1'b0,s4[58]};
assign {s39[60],s38[59]} = {1'b0,s6[59]} + {1'b0,s5[59]} + {1'b0,s4[59]};
assign {s39[61],s38[60]} = {1'b0,s6[60]} + {1'b0,s5[60]} + {1'b0,s4[60]};
assign {s39[62],s38[61]} = {1'b0,s6[61]} + {1'b0,s5[61]} + {1'b0,s4[61]};
assign {s39[63],s38[62]} = {1'b0,s6[62]} + {1'b0,s5[62]} + {1'b0,s4[62]};
assign {s39[64],s38[63]} = {1'b0,s6[63]} + {1'b0,s5[63]} + {1'b0,s4[63]};
assign {s39[65],s38[64]} = {1'b0,s6[64]} + {1'b0,s5[64]} + {1'b0,s4[64]};
assign {s39[66],s38[65]} = {1'b0,s6[65]} + {1'b0,s5[65]} + {1'b0,s4[65]};
assign {s39[67],s38[66]} = {1'b0,s6[66]} + {1'b0,s5[66]} + {1'b0,s4[66]};
assign {s41[4],s40[3]} = {1'b0,s7[3]};
assign {s41[5],s40[4]} = {1'b0,s8[4]} + {1'b0,s7[4]};
assign {s41[6],s40[5]} = {1'b0,s9[5]} + {1'b0,s8[5]} + {1'b0,s7[5]};
assign {s41[7],s40[6]} = {1'b0,s9[6]} + {1'b0,s8[6]} + {1'b0,s7[6]};
assign {s41[8],s40[7]} = {1'b0,s9[7]} + {1'b0,s8[7]} + {1'b0,s7[7]};
assign {s41[9],s40[8]} = {1'b0,s9[8]} + {1'b0,s8[8]} + {1'b0,s7[8]};
assign {s41[10],s40[9]} = {1'b0,s9[9]} + {1'b0,s8[9]} + {1'b0,s7[9]};
assign {s41[11],s40[10]} = {1'b0,s9[10]} + {1'b0,s8[10]} + {1'b0,s7[10]};
assign {s41[12],s40[11]} = {1'b0,s9[11]} + {1'b0,s8[11]} + {1'b0,s7[11]};
assign {s41[13],s40[12]} = {1'b0,s9[12]} + {1'b0,s8[12]} + {1'b0,s7[12]};
assign {s41[14],s40[13]} = {1'b0,s9[13]} + {1'b0,s8[13]} + {1'b0,s7[13]};
assign {s41[15],s40[14]} = {1'b0,s9[14]} + {1'b0,s8[14]} + {1'b0,s7[14]};
assign {s41[16],s40[15]} = {1'b0,s9[15]} + {1'b0,s8[15]} + {1'b0,s7[15]};
assign {s41[17],s40[16]} = {1'b0,s9[16]} + {1'b0,s8[16]} + {1'b0,s7[16]};
assign {s41[18],s40[17]} = {1'b0,s9[17]} + {1'b0,s8[17]} + {1'b0,s7[17]};
assign {s41[19],s40[18]} = {1'b0,s9[18]} + {1'b0,s8[18]} + {1'b0,s7[18]};
assign {s41[20],s40[19]} = {1'b0,s9[19]} + {1'b0,s8[19]} + {1'b0,s7[19]};
assign {s41[21],s40[20]} = {1'b0,s9[20]} + {1'b0,s8[20]} + {1'b0,s7[20]};
assign {s41[22],s40[21]} = {1'b0,s9[21]} + {1'b0,s8[21]} + {1'b0,s7[21]};
assign {s41[23],s40[22]} = {1'b0,s9[22]} + {1'b0,s8[22]} + {1'b0,s7[22]};
assign {s41[24],s40[23]} = {1'b0,s9[23]} + {1'b0,s8[23]} + {1'b0,s7[23]};
assign {s41[25],s40[24]} = {1'b0,s9[24]} + {1'b0,s8[24]} + {1'b0,s7[24]};
assign {s41[26],s40[25]} = {1'b0,s9[25]} + {1'b0,s8[25]} + {1'b0,s7[25]};
assign {s41[27],s40[26]} = {1'b0,s9[26]} + {1'b0,s8[26]} + {1'b0,s7[26]};
assign {s41[28],s40[27]} = {1'b0,s9[27]} + {1'b0,s8[27]} + {1'b0,s7[27]};
assign {s41[29],s40[28]} = {1'b0,s9[28]} + {1'b0,s8[28]} + {1'b0,s7[28]};
assign {s41[30],s40[29]} = {1'b0,s9[29]} + {1'b0,s8[29]} + {1'b0,s7[29]};
assign {s41[31],s40[30]} = {1'b0,s9[30]} + {1'b0,s8[30]} + {1'b0,s7[30]};
assign {s41[32],s40[31]} = {1'b0,s9[31]} + {1'b0,s8[31]} + {1'b0,s7[31]};
assign {s41[33],s40[32]} = {1'b0,s9[32]} + {1'b0,s8[32]} + {1'b0,s7[32]};
assign {s41[34],s40[33]} = {1'b0,s9[33]} + {1'b0,s8[33]} + {1'b0,s7[33]};
assign {s41[35],s40[34]} = {1'b0,s9[34]} + {1'b0,s8[34]} + {1'b0,s7[34]};
assign {s41[36],s40[35]} = {1'b0,s9[35]} + {1'b0,s8[35]} + {1'b0,s7[35]};
assign {s41[37],s40[36]} = {1'b0,s9[36]} + {1'b0,s8[36]} + {1'b0,s7[36]};
assign {s41[38],s40[37]} = {1'b0,s9[37]} + {1'b0,s8[37]} + {1'b0,s7[37]};
assign {s41[39],s40[38]} = {1'b0,s9[38]} + {1'b0,s8[38]} + {1'b0,s7[38]};
assign {s41[40],s40[39]} = {1'b0,s9[39]} + {1'b0,s8[39]} + {1'b0,s7[39]};
assign {s41[41],s40[40]} = {1'b0,s9[40]} + {1'b0,s8[40]} + {1'b0,s7[40]};
assign {s41[42],s40[41]} = {1'b0,s9[41]} + {1'b0,s8[41]} + {1'b0,s7[41]};
assign {s41[43],s40[42]} = {1'b0,s9[42]} + {1'b0,s8[42]} + {1'b0,s7[42]};
assign {s41[44],s40[43]} = {1'b0,s9[43]} + {1'b0,s8[43]} + {1'b0,s7[43]};
assign {s41[45],s40[44]} = {1'b0,s9[44]} + {1'b0,s8[44]} + {1'b0,s7[44]};
assign {s41[46],s40[45]} = {1'b0,s9[45]} + {1'b0,s8[45]} + {1'b0,s7[45]};
assign {s41[47],s40[46]} = {1'b0,s9[46]} + {1'b0,s8[46]} + {1'b0,s7[46]};
assign {s41[48],s40[47]} = {1'b0,s9[47]} + {1'b0,s8[47]} + {1'b0,s7[47]};
assign {s41[49],s40[48]} = {1'b0,s9[48]} + {1'b0,s8[48]} + {1'b0,s7[48]};
assign {s41[50],s40[49]} = {1'b0,s9[49]} + {1'b0,s8[49]} + {1'b0,s7[49]};
assign {s41[51],s40[50]} = {1'b0,s9[50]} + {1'b0,s8[50]} + {1'b0,s7[50]};
assign {s41[52],s40[51]} = {1'b0,s9[51]} + {1'b0,s8[51]} + {1'b0,s7[51]};
assign {s41[53],s40[52]} = {1'b0,s9[52]} + {1'b0,s8[52]} + {1'b0,s7[52]};
assign {s41[54],s40[53]} = {1'b0,s9[53]} + {1'b0,s8[53]} + {1'b0,s7[53]};
assign {s41[55],s40[54]} = {1'b0,s9[54]} + {1'b0,s8[54]} + {1'b0,s7[54]};
assign {s41[56],s40[55]} = {1'b0,s9[55]} + {1'b0,s8[55]} + {1'b0,s7[55]};
assign {s41[57],s40[56]} = {1'b0,s9[56]} + {1'b0,s8[56]} + {1'b0,s7[56]};
assign {s41[58],s40[57]} = {1'b0,s9[57]} + {1'b0,s8[57]} + {1'b0,s7[57]};
assign {s41[59],s40[58]} = {1'b0,s9[58]} + {1'b0,s8[58]} + {1'b0,s7[58]};
assign {s41[60],s40[59]} = {1'b0,s9[59]} + {1'b0,s8[59]} + {1'b0,s7[59]};
assign {s41[61],s40[60]} = {1'b0,s9[60]} + {1'b0,s8[60]} + {1'b0,s7[60]};
assign {s41[62],s40[61]} = {1'b0,s9[61]} + {1'b0,s8[61]} + {1'b0,s7[61]};
assign {s41[63],s40[62]} = {1'b0,s9[62]} + {1'b0,s8[62]} + {1'b0,s7[62]};
assign {s41[64],s40[63]} = {1'b0,s9[63]} + {1'b0,s8[63]} + {1'b0,s7[63]};
assign {s41[65],s40[64]} = {1'b0,s9[64]} + {1'b0,s8[64]} + {1'b0,s7[64]};
assign {s41[66],s40[65]} = {1'b0,s9[65]} + {1'b0,s8[65]} + {1'b0,s7[65]};
assign {s41[67],s40[66]} = {1'b0,s9[66]} + {1'b0,s8[66]} + {1'b0,s7[66]};
assign {s43[7],s42[6]} = {1'b0,s10[6]};
assign {s43[8],s42[7]} = {1'b0,s11[7]} + {1'b0,s10[7]};
assign {s43[9],s42[8]} = {1'b0,s12[8]} + {1'b0,s11[8]} + {1'b0,s10[8]};
assign {s43[10],s42[9]} = {1'b0,s12[9]} + {1'b0,s11[9]} + {1'b0,s10[9]};
assign {s43[11],s42[10]} = {1'b0,s12[10]} + {1'b0,s11[10]} + {1'b0,s10[10]};
assign {s43[12],s42[11]} = {1'b0,s12[11]} + {1'b0,s11[11]} + {1'b0,s10[11]};
assign {s43[13],s42[12]} = {1'b0,s12[12]} + {1'b0,s11[12]} + {1'b0,s10[12]};
assign {s43[14],s42[13]} = {1'b0,s12[13]} + {1'b0,s11[13]} + {1'b0,s10[13]};
assign {s43[15],s42[14]} = {1'b0,s12[14]} + {1'b0,s11[14]} + {1'b0,s10[14]};
assign {s43[16],s42[15]} = {1'b0,s12[15]} + {1'b0,s11[15]} + {1'b0,s10[15]};
assign {s43[17],s42[16]} = {1'b0,s12[16]} + {1'b0,s11[16]} + {1'b0,s10[16]};
assign {s43[18],s42[17]} = {1'b0,s12[17]} + {1'b0,s11[17]} + {1'b0,s10[17]};
assign {s43[19],s42[18]} = {1'b0,s12[18]} + {1'b0,s11[18]} + {1'b0,s10[18]};
assign {s43[20],s42[19]} = {1'b0,s12[19]} + {1'b0,s11[19]} + {1'b0,s10[19]};
assign {s43[21],s42[20]} = {1'b0,s12[20]} + {1'b0,s11[20]} + {1'b0,s10[20]};
assign {s43[22],s42[21]} = {1'b0,s12[21]} + {1'b0,s11[21]} + {1'b0,s10[21]};
assign {s43[23],s42[22]} = {1'b0,s12[22]} + {1'b0,s11[22]} + {1'b0,s10[22]};
assign {s43[24],s42[23]} = {1'b0,s12[23]} + {1'b0,s11[23]} + {1'b0,s10[23]};
assign {s43[25],s42[24]} = {1'b0,s12[24]} + {1'b0,s11[24]} + {1'b0,s10[24]};
assign {s43[26],s42[25]} = {1'b0,s12[25]} + {1'b0,s11[25]} + {1'b0,s10[25]};
assign {s43[27],s42[26]} = {1'b0,s12[26]} + {1'b0,s11[26]} + {1'b0,s10[26]};
assign {s43[28],s42[27]} = {1'b0,s12[27]} + {1'b0,s11[27]} + {1'b0,s10[27]};
assign {s43[29],s42[28]} = {1'b0,s12[28]} + {1'b0,s11[28]} + {1'b0,s10[28]};
assign {s43[30],s42[29]} = {1'b0,s12[29]} + {1'b0,s11[29]} + {1'b0,s10[29]};
assign {s43[31],s42[30]} = {1'b0,s12[30]} + {1'b0,s11[30]} + {1'b0,s10[30]};
assign {s43[32],s42[31]} = {1'b0,s12[31]} + {1'b0,s11[31]} + {1'b0,s10[31]};
assign {s43[33],s42[32]} = {1'b0,s12[32]} + {1'b0,s11[32]} + {1'b0,s10[32]};
assign {s43[34],s42[33]} = {1'b0,s12[33]} + {1'b0,s11[33]} + {1'b0,s10[33]};
assign {s43[35],s42[34]} = {1'b0,s12[34]} + {1'b0,s11[34]} + {1'b0,s10[34]};
assign {s43[36],s42[35]} = {1'b0,s12[35]} + {1'b0,s11[35]} + {1'b0,s10[35]};
assign {s43[37],s42[36]} = {1'b0,s12[36]} + {1'b0,s11[36]} + {1'b0,s10[36]};
assign {s43[38],s42[37]} = {1'b0,s12[37]} + {1'b0,s11[37]} + {1'b0,s10[37]};
assign {s43[39],s42[38]} = {1'b0,s12[38]} + {1'b0,s11[38]} + {1'b0,s10[38]};
assign {s43[40],s42[39]} = {1'b0,s12[39]} + {1'b0,s11[39]} + {1'b0,s10[39]};
assign {s43[41],s42[40]} = {1'b0,s12[40]} + {1'b0,s11[40]} + {1'b0,s10[40]};
assign {s43[42],s42[41]} = {1'b0,s12[41]} + {1'b0,s11[41]} + {1'b0,s10[41]};
assign {s43[43],s42[42]} = {1'b0,s12[42]} + {1'b0,s11[42]} + {1'b0,s10[42]};
assign {s43[44],s42[43]} = {1'b0,s12[43]} + {1'b0,s11[43]} + {1'b0,s10[43]};
assign {s43[45],s42[44]} = {1'b0,s12[44]} + {1'b0,s11[44]} + {1'b0,s10[44]};
assign {s43[46],s42[45]} = {1'b0,s12[45]} + {1'b0,s11[45]} + {1'b0,s10[45]};
assign {s43[47],s42[46]} = {1'b0,s12[46]} + {1'b0,s11[46]} + {1'b0,s10[46]};
assign {s43[48],s42[47]} = {1'b0,s12[47]} + {1'b0,s11[47]} + {1'b0,s10[47]};
assign {s43[49],s42[48]} = {1'b0,s12[48]} + {1'b0,s11[48]} + {1'b0,s10[48]};
assign {s43[50],s42[49]} = {1'b0,s12[49]} + {1'b0,s11[49]} + {1'b0,s10[49]};
assign {s43[51],s42[50]} = {1'b0,s12[50]} + {1'b0,s11[50]} + {1'b0,s10[50]};
assign {s43[52],s42[51]} = {1'b0,s12[51]} + {1'b0,s11[51]} + {1'b0,s10[51]};
assign {s43[53],s42[52]} = {1'b0,s12[52]} + {1'b0,s11[52]} + {1'b0,s10[52]};
assign {s43[54],s42[53]} = {1'b0,s12[53]} + {1'b0,s11[53]} + {1'b0,s10[53]};
assign {s43[55],s42[54]} = {1'b0,s12[54]} + {1'b0,s11[54]} + {1'b0,s10[54]};
assign {s43[56],s42[55]} = {1'b0,s12[55]} + {1'b0,s11[55]} + {1'b0,s10[55]};
assign {s43[57],s42[56]} = {1'b0,s12[56]} + {1'b0,s11[56]} + {1'b0,s10[56]};
assign {s43[58],s42[57]} = {1'b0,s12[57]} + {1'b0,s11[57]} + {1'b0,s10[57]};
assign {s43[59],s42[58]} = {1'b0,s12[58]} + {1'b0,s11[58]} + {1'b0,s10[58]};
assign {s43[60],s42[59]} = {1'b0,s12[59]} + {1'b0,s11[59]} + {1'b0,s10[59]};
assign {s43[61],s42[60]} = {1'b0,s12[60]} + {1'b0,s11[60]} + {1'b0,s10[60]};
assign {s43[62],s42[61]} = {1'b0,s12[61]} + {1'b0,s11[61]} + {1'b0,s10[61]};
assign {s43[63],s42[62]} = {1'b0,s12[62]} + {1'b0,s11[62]} + {1'b0,s10[62]};
assign {s43[64],s42[63]} = {1'b0,s12[63]} + {1'b0,s11[63]} + {1'b0,s10[63]};
assign {s43[65],s42[64]} = {1'b0,s12[64]} + {1'b0,s11[64]} + {1'b0,s10[64]};
assign {s43[66],s42[65]} = {1'b0,s12[65]} + {1'b0,s11[65]} + {1'b0,s10[65]};
assign {s43[67],s42[66]} = {1'b0,s12[66]} + {1'b0,s11[66]} + {1'b0,s10[66]};
assign {s45[10],s44[9]} = {1'b0,s13[9]};
assign {s45[11],s44[10]} = {1'b0,s14[10]} + {1'b0,s13[10]};
assign {s45[12],s44[11]} = {1'b0,s15[11]} + {1'b0,s14[11]} + {1'b0,s13[11]};
assign {s45[13],s44[12]} = {1'b0,s15[12]} + {1'b0,s14[12]} + {1'b0,s13[12]};
assign {s45[14],s44[13]} = {1'b0,s15[13]} + {1'b0,s14[13]} + {1'b0,s13[13]};
assign {s45[15],s44[14]} = {1'b0,s15[14]} + {1'b0,s14[14]} + {1'b0,s13[14]};
assign {s45[16],s44[15]} = {1'b0,s15[15]} + {1'b0,s14[15]} + {1'b0,s13[15]};
assign {s45[17],s44[16]} = {1'b0,s15[16]} + {1'b0,s14[16]} + {1'b0,s13[16]};
assign {s45[18],s44[17]} = {1'b0,s15[17]} + {1'b0,s14[17]} + {1'b0,s13[17]};
assign {s45[19],s44[18]} = {1'b0,s15[18]} + {1'b0,s14[18]} + {1'b0,s13[18]};
assign {s45[20],s44[19]} = {1'b0,s15[19]} + {1'b0,s14[19]} + {1'b0,s13[19]};
assign {s45[21],s44[20]} = {1'b0,s15[20]} + {1'b0,s14[20]} + {1'b0,s13[20]};
assign {s45[22],s44[21]} = {1'b0,s15[21]} + {1'b0,s14[21]} + {1'b0,s13[21]};
assign {s45[23],s44[22]} = {1'b0,s15[22]} + {1'b0,s14[22]} + {1'b0,s13[22]};
assign {s45[24],s44[23]} = {1'b0,s15[23]} + {1'b0,s14[23]} + {1'b0,s13[23]};
assign {s45[25],s44[24]} = {1'b0,s15[24]} + {1'b0,s14[24]} + {1'b0,s13[24]};
assign {s45[26],s44[25]} = {1'b0,s15[25]} + {1'b0,s14[25]} + {1'b0,s13[25]};
assign {s45[27],s44[26]} = {1'b0,s15[26]} + {1'b0,s14[26]} + {1'b0,s13[26]};
assign {s45[28],s44[27]} = {1'b0,s15[27]} + {1'b0,s14[27]} + {1'b0,s13[27]};
assign {s45[29],s44[28]} = {1'b0,s15[28]} + {1'b0,s14[28]} + {1'b0,s13[28]};
assign {s45[30],s44[29]} = {1'b0,s15[29]} + {1'b0,s14[29]} + {1'b0,s13[29]};
assign {s45[31],s44[30]} = {1'b0,s15[30]} + {1'b0,s14[30]} + {1'b0,s13[30]};
assign {s45[32],s44[31]} = {1'b0,s15[31]} + {1'b0,s14[31]} + {1'b0,s13[31]};
assign {s45[33],s44[32]} = {1'b0,s15[32]} + {1'b0,s14[32]} + {1'b0,s13[32]};
assign {s45[34],s44[33]} = {1'b0,s15[33]} + {1'b0,s14[33]} + {1'b0,s13[33]};
assign {s45[35],s44[34]} = {1'b0,s15[34]} + {1'b0,s14[34]} + {1'b0,s13[34]};
assign {s45[36],s44[35]} = {1'b0,s15[35]} + {1'b0,s14[35]} + {1'b0,s13[35]};
assign {s45[37],s44[36]} = {1'b0,s15[36]} + {1'b0,s14[36]} + {1'b0,s13[36]};
assign {s45[38],s44[37]} = {1'b0,s15[37]} + {1'b0,s14[37]} + {1'b0,s13[37]};
assign {s45[39],s44[38]} = {1'b0,s15[38]} + {1'b0,s14[38]} + {1'b0,s13[38]};
assign {s45[40],s44[39]} = {1'b0,s15[39]} + {1'b0,s14[39]} + {1'b0,s13[39]};
assign {s45[41],s44[40]} = {1'b0,s15[40]} + {1'b0,s14[40]} + {1'b0,s13[40]};
assign {s45[42],s44[41]} = {1'b0,s15[41]} + {1'b0,s14[41]} + {1'b0,s13[41]};
assign {s45[43],s44[42]} = {1'b0,s15[42]} + {1'b0,s14[42]} + {1'b0,s13[42]};
assign {s45[44],s44[43]} = {1'b0,s15[43]} + {1'b0,s14[43]} + {1'b0,s13[43]};
assign {s45[45],s44[44]} = {1'b0,s15[44]} + {1'b0,s14[44]} + {1'b0,s13[44]};
assign {s45[46],s44[45]} = {1'b0,s15[45]} + {1'b0,s14[45]} + {1'b0,s13[45]};
assign {s45[47],s44[46]} = {1'b0,s15[46]} + {1'b0,s14[46]} + {1'b0,s13[46]};
assign {s45[48],s44[47]} = {1'b0,s15[47]} + {1'b0,s14[47]} + {1'b0,s13[47]};
assign {s45[49],s44[48]} = {1'b0,s15[48]} + {1'b0,s14[48]} + {1'b0,s13[48]};
assign {s45[50],s44[49]} = {1'b0,s15[49]} + {1'b0,s14[49]} + {1'b0,s13[49]};
assign {s45[51],s44[50]} = {1'b0,s15[50]} + {1'b0,s14[50]} + {1'b0,s13[50]};
assign {s45[52],s44[51]} = {1'b0,s15[51]} + {1'b0,s14[51]} + {1'b0,s13[51]};
assign {s45[53],s44[52]} = {1'b0,s15[52]} + {1'b0,s14[52]} + {1'b0,s13[52]};
assign {s45[54],s44[53]} = {1'b0,s15[53]} + {1'b0,s14[53]} + {1'b0,s13[53]};
assign {s45[55],s44[54]} = {1'b0,s15[54]} + {1'b0,s14[54]} + {1'b0,s13[54]};
assign {s45[56],s44[55]} = {1'b0,s15[55]} + {1'b0,s14[55]} + {1'b0,s13[55]};
assign {s45[57],s44[56]} = {1'b0,s15[56]} + {1'b0,s14[56]} + {1'b0,s13[56]};
assign {s45[58],s44[57]} = {1'b0,s15[57]} + {1'b0,s14[57]} + {1'b0,s13[57]};
assign {s45[59],s44[58]} = {1'b0,s15[58]} + {1'b0,s14[58]} + {1'b0,s13[58]};
assign {s45[60],s44[59]} = {1'b0,s15[59]} + {1'b0,s14[59]} + {1'b0,s13[59]};
assign {s45[61],s44[60]} = {1'b0,s15[60]} + {1'b0,s14[60]} + {1'b0,s13[60]};
assign {s45[62],s44[61]} = {1'b0,s15[61]} + {1'b0,s14[61]} + {1'b0,s13[61]};
assign {s45[63],s44[62]} = {1'b0,s15[62]} + {1'b0,s14[62]} + {1'b0,s13[62]};
assign {s45[64],s44[63]} = {1'b0,s15[63]} + {1'b0,s14[63]} + {1'b0,s13[63]};
assign {s45[65],s44[64]} = {1'b0,s15[64]} + {1'b0,s14[64]} + {1'b0,s13[64]};
assign {s45[66],s44[65]} = {1'b0,s15[65]} + {1'b0,s14[65]} + {1'b0,s13[65]};
assign {s45[67],s44[66]} = {1'b0,s15[66]} + {1'b0,s14[66]} + {1'b0,s13[66]};
assign {s47[13],s46[12]} = {1'b0,s16[12]};
assign {s47[14],s46[13]} = {1'b0,s17[13]} + {1'b0,s16[13]};
assign {s47[15],s46[14]} = {1'b0,s18[14]} + {1'b0,s17[14]} + {1'b0,s16[14]};
assign {s47[16],s46[15]} = {1'b0,s18[15]} + {1'b0,s17[15]} + {1'b0,s16[15]};
assign {s47[17],s46[16]} = {1'b0,s18[16]} + {1'b0,s17[16]} + {1'b0,s16[16]};
assign {s47[18],s46[17]} = {1'b0,s18[17]} + {1'b0,s17[17]} + {1'b0,s16[17]};
assign {s47[19],s46[18]} = {1'b0,s18[18]} + {1'b0,s17[18]} + {1'b0,s16[18]};
assign {s47[20],s46[19]} = {1'b0,s18[19]} + {1'b0,s17[19]} + {1'b0,s16[19]};
assign {s47[21],s46[20]} = {1'b0,s18[20]} + {1'b0,s17[20]} + {1'b0,s16[20]};
assign {s47[22],s46[21]} = {1'b0,s18[21]} + {1'b0,s17[21]} + {1'b0,s16[21]};
assign {s47[23],s46[22]} = {1'b0,s18[22]} + {1'b0,s17[22]} + {1'b0,s16[22]};
assign {s47[24],s46[23]} = {1'b0,s18[23]} + {1'b0,s17[23]} + {1'b0,s16[23]};
assign {s47[25],s46[24]} = {1'b0,s18[24]} + {1'b0,s17[24]} + {1'b0,s16[24]};
assign {s47[26],s46[25]} = {1'b0,s18[25]} + {1'b0,s17[25]} + {1'b0,s16[25]};
assign {s47[27],s46[26]} = {1'b0,s18[26]} + {1'b0,s17[26]} + {1'b0,s16[26]};
assign {s47[28],s46[27]} = {1'b0,s18[27]} + {1'b0,s17[27]} + {1'b0,s16[27]};
assign {s47[29],s46[28]} = {1'b0,s18[28]} + {1'b0,s17[28]} + {1'b0,s16[28]};
assign {s47[30],s46[29]} = {1'b0,s18[29]} + {1'b0,s17[29]} + {1'b0,s16[29]};
assign {s47[31],s46[30]} = {1'b0,s18[30]} + {1'b0,s17[30]} + {1'b0,s16[30]};
assign {s47[32],s46[31]} = {1'b0,s18[31]} + {1'b0,s17[31]} + {1'b0,s16[31]};
assign {s47[33],s46[32]} = {1'b0,s18[32]} + {1'b0,s17[32]} + {1'b0,s16[32]};
assign {s47[34],s46[33]} = {1'b0,s18[33]} + {1'b0,s17[33]} + {1'b0,s16[33]};
assign {s47[35],s46[34]} = {1'b0,s18[34]} + {1'b0,s17[34]} + {1'b0,s16[34]};
assign {s47[36],s46[35]} = {1'b0,s18[35]} + {1'b0,s17[35]} + {1'b0,s16[35]};
assign {s47[37],s46[36]} = {1'b0,s18[36]} + {1'b0,s17[36]} + {1'b0,s16[36]};
assign {s47[38],s46[37]} = {1'b0,s18[37]} + {1'b0,s17[37]} + {1'b0,s16[37]};
assign {s47[39],s46[38]} = {1'b0,s18[38]} + {1'b0,s17[38]} + {1'b0,s16[38]};
assign {s47[40],s46[39]} = {1'b0,s18[39]} + {1'b0,s17[39]} + {1'b0,s16[39]};
assign {s47[41],s46[40]} = {1'b0,s18[40]} + {1'b0,s17[40]} + {1'b0,s16[40]};
assign {s47[42],s46[41]} = {1'b0,s18[41]} + {1'b0,s17[41]} + {1'b0,s16[41]};
assign {s47[43],s46[42]} = {1'b0,s18[42]} + {1'b0,s17[42]} + {1'b0,s16[42]};
assign {s47[44],s46[43]} = {1'b0,s18[43]} + {1'b0,s17[43]} + {1'b0,s16[43]};
assign {s47[45],s46[44]} = {1'b0,s18[44]} + {1'b0,s17[44]} + {1'b0,s16[44]};
assign {s47[46],s46[45]} = {1'b0,s18[45]} + {1'b0,s17[45]} + {1'b0,s16[45]};
assign {s47[47],s46[46]} = {1'b0,s18[46]} + {1'b0,s17[46]} + {1'b0,s16[46]};
assign {s47[48],s46[47]} = {1'b0,s18[47]} + {1'b0,s17[47]} + {1'b0,s16[47]};
assign {s47[49],s46[48]} = {1'b0,s18[48]} + {1'b0,s17[48]} + {1'b0,s16[48]};
assign {s47[50],s46[49]} = {1'b0,s18[49]} + {1'b0,s17[49]} + {1'b0,s16[49]};
assign {s47[51],s46[50]} = {1'b0,s18[50]} + {1'b0,s17[50]} + {1'b0,s16[50]};
assign {s47[52],s46[51]} = {1'b0,s18[51]} + {1'b0,s17[51]} + {1'b0,s16[51]};
assign {s47[53],s46[52]} = {1'b0,s18[52]} + {1'b0,s17[52]} + {1'b0,s16[52]};
assign {s47[54],s46[53]} = {1'b0,s18[53]} + {1'b0,s17[53]} + {1'b0,s16[53]};
assign {s47[55],s46[54]} = {1'b0,s18[54]} + {1'b0,s17[54]} + {1'b0,s16[54]};
assign {s47[56],s46[55]} = {1'b0,s18[55]} + {1'b0,s17[55]} + {1'b0,s16[55]};
assign {s47[57],s46[56]} = {1'b0,s18[56]} + {1'b0,s17[56]} + {1'b0,s16[56]};
assign {s47[58],s46[57]} = {1'b0,s18[57]} + {1'b0,s17[57]} + {1'b0,s16[57]};
assign {s47[59],s46[58]} = {1'b0,s18[58]} + {1'b0,s17[58]} + {1'b0,s16[58]};
assign {s47[60],s46[59]} = {1'b0,s18[59]} + {1'b0,s17[59]} + {1'b0,s16[59]};
assign {s47[61],s46[60]} = {1'b0,s18[60]} + {1'b0,s17[60]} + {1'b0,s16[60]};
assign {s47[62],s46[61]} = {1'b0,s18[61]} + {1'b0,s17[61]} + {1'b0,s16[61]};
assign {s47[63],s46[62]} = {1'b0,s18[62]} + {1'b0,s17[62]} + {1'b0,s16[62]};
assign {s47[64],s46[63]} = {1'b0,s18[63]} + {1'b0,s17[63]} + {1'b0,s16[63]};
assign {s47[65],s46[64]} = {1'b0,s18[64]} + {1'b0,s17[64]} + {1'b0,s16[64]};
assign {s47[66],s46[65]} = {1'b0,s18[65]} + {1'b0,s17[65]} + {1'b0,s16[65]};
assign {s47[67],s46[66]} = {1'b0,s18[66]} + {1'b0,s17[66]} + {1'b0,s16[66]};
assign {s49[16],s48[15]} = {1'b0,s19[15]};
assign {s49[17],s48[16]} = {1'b0,s20[16]} + {1'b0,s19[16]};
assign {s49[18],s48[17]} = {1'b0,s21[17]} + {1'b0,s20[17]} + {1'b0,s19[17]};
assign {s49[19],s48[18]} = {1'b0,s21[18]} + {1'b0,s20[18]} + {1'b0,s19[18]};
assign {s49[20],s48[19]} = {1'b0,s21[19]} + {1'b0,s20[19]} + {1'b0,s19[19]};
assign {s49[21],s48[20]} = {1'b0,s21[20]} + {1'b0,s20[20]} + {1'b0,s19[20]};
assign {s49[22],s48[21]} = {1'b0,s21[21]} + {1'b0,s20[21]} + {1'b0,s19[21]};
assign {s49[23],s48[22]} = {1'b0,s21[22]} + {1'b0,s20[22]} + {1'b0,s19[22]};
assign {s49[24],s48[23]} = {1'b0,s21[23]} + {1'b0,s20[23]} + {1'b0,s19[23]};
assign {s49[25],s48[24]} = {1'b0,s21[24]} + {1'b0,s20[24]} + {1'b0,s19[24]};
assign {s49[26],s48[25]} = {1'b0,s21[25]} + {1'b0,s20[25]} + {1'b0,s19[25]};
assign {s49[27],s48[26]} = {1'b0,s21[26]} + {1'b0,s20[26]} + {1'b0,s19[26]};
assign {s49[28],s48[27]} = {1'b0,s21[27]} + {1'b0,s20[27]} + {1'b0,s19[27]};
assign {s49[29],s48[28]} = {1'b0,s21[28]} + {1'b0,s20[28]} + {1'b0,s19[28]};
assign {s49[30],s48[29]} = {1'b0,s21[29]} + {1'b0,s20[29]} + {1'b0,s19[29]};
assign {s49[31],s48[30]} = {1'b0,s21[30]} + {1'b0,s20[30]} + {1'b0,s19[30]};
assign {s49[32],s48[31]} = {1'b0,s21[31]} + {1'b0,s20[31]} + {1'b0,s19[31]};
assign {s49[33],s48[32]} = {1'b0,s21[32]} + {1'b0,s20[32]} + {1'b0,s19[32]};
assign {s49[34],s48[33]} = {1'b0,s21[33]} + {1'b0,s20[33]} + {1'b0,s19[33]};
assign {s49[35],s48[34]} = {1'b0,s21[34]} + {1'b0,s20[34]} + {1'b0,s19[34]};
assign {s49[36],s48[35]} = {1'b0,s21[35]} + {1'b0,s20[35]} + {1'b0,s19[35]};
assign {s49[37],s48[36]} = {1'b0,s21[36]} + {1'b0,s20[36]} + {1'b0,s19[36]};
assign {s49[38],s48[37]} = {1'b0,s21[37]} + {1'b0,s20[37]} + {1'b0,s19[37]};
assign {s49[39],s48[38]} = {1'b0,s21[38]} + {1'b0,s20[38]} + {1'b0,s19[38]};
assign {s49[40],s48[39]} = {1'b0,s21[39]} + {1'b0,s20[39]} + {1'b0,s19[39]};
assign {s49[41],s48[40]} = {1'b0,s21[40]} + {1'b0,s20[40]} + {1'b0,s19[40]};
assign {s49[42],s48[41]} = {1'b0,s21[41]} + {1'b0,s20[41]} + {1'b0,s19[41]};
assign {s49[43],s48[42]} = {1'b0,s21[42]} + {1'b0,s20[42]} + {1'b0,s19[42]};
assign {s49[44],s48[43]} = {1'b0,s21[43]} + {1'b0,s20[43]} + {1'b0,s19[43]};
assign {s49[45],s48[44]} = {1'b0,s21[44]} + {1'b0,s20[44]} + {1'b0,s19[44]};
assign {s49[46],s48[45]} = {1'b0,s21[45]} + {1'b0,s20[45]} + {1'b0,s19[45]};
assign {s49[47],s48[46]} = {1'b0,s21[46]} + {1'b0,s20[46]} + {1'b0,s19[46]};
assign {s49[48],s48[47]} = {1'b0,s21[47]} + {1'b0,s20[47]} + {1'b0,s19[47]};
assign {s49[49],s48[48]} = {1'b0,s21[48]} + {1'b0,s20[48]} + {1'b0,s19[48]};
assign {s49[50],s48[49]} = {1'b0,s21[49]} + {1'b0,s20[49]} + {1'b0,s19[49]};
assign {s49[51],s48[50]} = {1'b0,s21[50]} + {1'b0,s20[50]} + {1'b0,s19[50]};
assign {s49[52],s48[51]} = {1'b0,s21[51]} + {1'b0,s20[51]} + {1'b0,s19[51]};
assign {s49[53],s48[52]} = {1'b0,s21[52]} + {1'b0,s20[52]} + {1'b0,s19[52]};
assign {s49[54],s48[53]} = {1'b0,s21[53]} + {1'b0,s20[53]} + {1'b0,s19[53]};
assign {s49[55],s48[54]} = {1'b0,s21[54]} + {1'b0,s20[54]} + {1'b0,s19[54]};
assign {s49[56],s48[55]} = {1'b0,s21[55]} + {1'b0,s20[55]} + {1'b0,s19[55]};
assign {s49[57],s48[56]} = {1'b0,s21[56]} + {1'b0,s20[56]} + {1'b0,s19[56]};
assign {s49[58],s48[57]} = {1'b0,s21[57]} + {1'b0,s20[57]} + {1'b0,s19[57]};
assign {s49[59],s48[58]} = {1'b0,s21[58]} + {1'b0,s20[58]} + {1'b0,s19[58]};
assign {s49[60],s48[59]} = {1'b0,s21[59]} + {1'b0,s20[59]} + {1'b0,s19[59]};
assign {s49[61],s48[60]} = {1'b0,s21[60]} + {1'b0,s20[60]} + {1'b0,s19[60]};
assign {s49[62],s48[61]} = {1'b0,s21[61]} + {1'b0,s20[61]} + {1'b0,s19[61]};
assign {s49[63],s48[62]} = {1'b0,s21[62]} + {1'b0,s20[62]} + {1'b0,s19[62]};
assign {s49[64],s48[63]} = {1'b0,s21[63]} + {1'b0,s20[63]} + {1'b0,s19[63]};
assign {s49[65],s48[64]} = {1'b0,s21[64]} + {1'b0,s20[64]} + {1'b0,s19[64]};
assign {s49[66],s48[65]} = {1'b0,s21[65]} + {1'b0,s20[65]} + {1'b0,s19[65]};
assign {s49[67],s48[66]} = {1'b0,s21[66]} + {1'b0,s20[66]} + {1'b0,s19[66]};
assign {s51[19],s50[18]} = {1'b0,s22[18]};
assign {s51[20],s50[19]} = {1'b0,s23[19]} + {1'b0,s22[19]};
assign {s51[21],s50[20]} = {1'b0,s24[20]} + {1'b0,s23[20]} + {1'b0,s22[20]};
assign {s51[22],s50[21]} = {1'b0,s24[21]} + {1'b0,s23[21]} + {1'b0,s22[21]};
assign {s51[23],s50[22]} = {1'b0,s24[22]} + {1'b0,s23[22]} + {1'b0,s22[22]};
assign {s51[24],s50[23]} = {1'b0,s24[23]} + {1'b0,s23[23]} + {1'b0,s22[23]};
assign {s51[25],s50[24]} = {1'b0,s24[24]} + {1'b0,s23[24]} + {1'b0,s22[24]};
assign {s51[26],s50[25]} = {1'b0,s24[25]} + {1'b0,s23[25]} + {1'b0,s22[25]};
assign {s51[27],s50[26]} = {1'b0,s24[26]} + {1'b0,s23[26]} + {1'b0,s22[26]};
assign {s51[28],s50[27]} = {1'b0,s24[27]} + {1'b0,s23[27]} + {1'b0,s22[27]};
assign {s51[29],s50[28]} = {1'b0,s24[28]} + {1'b0,s23[28]} + {1'b0,s22[28]};
assign {s51[30],s50[29]} = {1'b0,s24[29]} + {1'b0,s23[29]} + {1'b0,s22[29]};
assign {s51[31],s50[30]} = {1'b0,s24[30]} + {1'b0,s23[30]} + {1'b0,s22[30]};
assign {s51[32],s50[31]} = {1'b0,s24[31]} + {1'b0,s23[31]} + {1'b0,s22[31]};
assign {s51[33],s50[32]} = {1'b0,s24[32]} + {1'b0,s23[32]} + {1'b0,s22[32]};
assign {s51[34],s50[33]} = {1'b0,s24[33]} + {1'b0,s23[33]} + {1'b0,s22[33]};
assign {s51[35],s50[34]} = {1'b0,s24[34]} + {1'b0,s23[34]} + {1'b0,s22[34]};
assign {s51[36],s50[35]} = {1'b0,s24[35]} + {1'b0,s23[35]} + {1'b0,s22[35]};
assign {s51[37],s50[36]} = {1'b0,s24[36]} + {1'b0,s23[36]} + {1'b0,s22[36]};
assign {s51[38],s50[37]} = {1'b0,s24[37]} + {1'b0,s23[37]} + {1'b0,s22[37]};
assign {s51[39],s50[38]} = {1'b0,s24[38]} + {1'b0,s23[38]} + {1'b0,s22[38]};
assign {s51[40],s50[39]} = {1'b0,s24[39]} + {1'b0,s23[39]} + {1'b0,s22[39]};
assign {s51[41],s50[40]} = {1'b0,s24[40]} + {1'b0,s23[40]} + {1'b0,s22[40]};
assign {s51[42],s50[41]} = {1'b0,s24[41]} + {1'b0,s23[41]} + {1'b0,s22[41]};
assign {s51[43],s50[42]} = {1'b0,s24[42]} + {1'b0,s23[42]} + {1'b0,s22[42]};
assign {s51[44],s50[43]} = {1'b0,s24[43]} + {1'b0,s23[43]} + {1'b0,s22[43]};
assign {s51[45],s50[44]} = {1'b0,s24[44]} + {1'b0,s23[44]} + {1'b0,s22[44]};
assign {s51[46],s50[45]} = {1'b0,s24[45]} + {1'b0,s23[45]} + {1'b0,s22[45]};
assign {s51[47],s50[46]} = {1'b0,s24[46]} + {1'b0,s23[46]} + {1'b0,s22[46]};
assign {s51[48],s50[47]} = {1'b0,s24[47]} + {1'b0,s23[47]} + {1'b0,s22[47]};
assign {s51[49],s50[48]} = {1'b0,s24[48]} + {1'b0,s23[48]} + {1'b0,s22[48]};
assign {s51[50],s50[49]} = {1'b0,s24[49]} + {1'b0,s23[49]} + {1'b0,s22[49]};
assign {s51[51],s50[50]} = {1'b0,s24[50]} + {1'b0,s23[50]} + {1'b0,s22[50]};
assign {s51[52],s50[51]} = {1'b0,s24[51]} + {1'b0,s23[51]} + {1'b0,s22[51]};
assign {s51[53],s50[52]} = {1'b0,s24[52]} + {1'b0,s23[52]} + {1'b0,s22[52]};
assign {s51[54],s50[53]} = {1'b0,s24[53]} + {1'b0,s23[53]} + {1'b0,s22[53]};
assign {s51[55],s50[54]} = {1'b0,s24[54]} + {1'b0,s23[54]} + {1'b0,s22[54]};
assign {s51[56],s50[55]} = {1'b0,s24[55]} + {1'b0,s23[55]} + {1'b0,s22[55]};
assign {s51[57],s50[56]} = {1'b0,s24[56]} + {1'b0,s23[56]} + {1'b0,s22[56]};
assign {s51[58],s50[57]} = {1'b0,s24[57]} + {1'b0,s23[57]} + {1'b0,s22[57]};
assign {s51[59],s50[58]} = {1'b0,s24[58]} + {1'b0,s23[58]} + {1'b0,s22[58]};
assign {s51[60],s50[59]} = {1'b0,s24[59]} + {1'b0,s23[59]} + {1'b0,s22[59]};
assign {s51[61],s50[60]} = {1'b0,s24[60]} + {1'b0,s23[60]} + {1'b0,s22[60]};
assign {s51[62],s50[61]} = {1'b0,s24[61]} + {1'b0,s23[61]} + {1'b0,s22[61]};
assign {s51[63],s50[62]} = {1'b0,s24[62]} + {1'b0,s23[62]} + {1'b0,s22[62]};
assign {s51[64],s50[63]} = {1'b0,s24[63]} + {1'b0,s23[63]} + {1'b0,s22[63]};
assign {s51[65],s50[64]} = {1'b0,s24[64]} + {1'b0,s23[64]} + {1'b0,s22[64]};
assign {s51[66],s50[65]} = {1'b0,s24[65]} + {1'b0,s23[65]} + {1'b0,s22[65]};
assign {s51[67],s50[66]} = {1'b0,s24[66]} + {1'b0,s23[66]} + {1'b0,s22[66]};
assign {s53[22],s52[21]} = {1'b0,s25[21]};
assign {s53[23],s52[22]} = {1'b0,s26[22]} + {1'b0,s25[22]};
assign {s53[24],s52[23]} = {1'b0,s27[23]} + {1'b0,s26[23]} + {1'b0,s25[23]};
assign {s53[25],s52[24]} = {1'b0,s27[24]} + {1'b0,s26[24]} + {1'b0,s25[24]};
assign {s53[26],s52[25]} = {1'b0,s27[25]} + {1'b0,s26[25]} + {1'b0,s25[25]};
assign {s53[27],s52[26]} = {1'b0,s27[26]} + {1'b0,s26[26]} + {1'b0,s25[26]};
assign {s53[28],s52[27]} = {1'b0,s27[27]} + {1'b0,s26[27]} + {1'b0,s25[27]};
assign {s53[29],s52[28]} = {1'b0,s27[28]} + {1'b0,s26[28]} + {1'b0,s25[28]};
assign {s53[30],s52[29]} = {1'b0,s27[29]} + {1'b0,s26[29]} + {1'b0,s25[29]};
assign {s53[31],s52[30]} = {1'b0,s27[30]} + {1'b0,s26[30]} + {1'b0,s25[30]};
assign {s53[32],s52[31]} = {1'b0,s27[31]} + {1'b0,s26[31]} + {1'b0,s25[31]};
assign {s53[33],s52[32]} = {1'b0,s27[32]} + {1'b0,s26[32]} + {1'b0,s25[32]};
assign {s53[34],s52[33]} = {1'b0,s27[33]} + {1'b0,s26[33]} + {1'b0,s25[33]};
assign {s53[35],s52[34]} = {1'b0,s27[34]} + {1'b0,s26[34]} + {1'b0,s25[34]};
assign {s53[36],s52[35]} = {1'b0,s27[35]} + {1'b0,s26[35]} + {1'b0,s25[35]};
assign {s53[37],s52[36]} = {1'b0,s27[36]} + {1'b0,s26[36]} + {1'b0,s25[36]};
assign {s53[38],s52[37]} = {1'b0,s27[37]} + {1'b0,s26[37]} + {1'b0,s25[37]};
assign {s53[39],s52[38]} = {1'b0,s27[38]} + {1'b0,s26[38]} + {1'b0,s25[38]};
assign {s53[40],s52[39]} = {1'b0,s27[39]} + {1'b0,s26[39]} + {1'b0,s25[39]};
assign {s53[41],s52[40]} = {1'b0,s27[40]} + {1'b0,s26[40]} + {1'b0,s25[40]};
assign {s53[42],s52[41]} = {1'b0,s27[41]} + {1'b0,s26[41]} + {1'b0,s25[41]};
assign {s53[43],s52[42]} = {1'b0,s27[42]} + {1'b0,s26[42]} + {1'b0,s25[42]};
assign {s53[44],s52[43]} = {1'b0,s27[43]} + {1'b0,s26[43]} + {1'b0,s25[43]};
assign {s53[45],s52[44]} = {1'b0,s27[44]} + {1'b0,s26[44]} + {1'b0,s25[44]};
assign {s53[46],s52[45]} = {1'b0,s27[45]} + {1'b0,s26[45]} + {1'b0,s25[45]};
assign {s53[47],s52[46]} = {1'b0,s27[46]} + {1'b0,s26[46]} + {1'b0,s25[46]};
assign {s53[48],s52[47]} = {1'b0,s27[47]} + {1'b0,s26[47]} + {1'b0,s25[47]};
assign {s53[49],s52[48]} = {1'b0,s27[48]} + {1'b0,s26[48]} + {1'b0,s25[48]};
assign {s53[50],s52[49]} = {1'b0,s27[49]} + {1'b0,s26[49]} + {1'b0,s25[49]};
assign {s53[51],s52[50]} = {1'b0,s27[50]} + {1'b0,s26[50]} + {1'b0,s25[50]};
assign {s53[52],s52[51]} = {1'b0,s27[51]} + {1'b0,s26[51]} + {1'b0,s25[51]};
assign {s53[53],s52[52]} = {1'b0,s27[52]} + {1'b0,s26[52]} + {1'b0,s25[52]};
assign {s53[54],s52[53]} = {1'b0,s27[53]} + {1'b0,s26[53]} + {1'b0,s25[53]};
assign {s53[55],s52[54]} = {1'b0,s27[54]} + {1'b0,s26[54]} + {1'b0,s25[54]};
assign {s53[56],s52[55]} = {1'b0,s27[55]} + {1'b0,s26[55]} + {1'b0,s25[55]};
assign {s53[57],s52[56]} = {1'b0,s27[56]} + {1'b0,s26[56]} + {1'b0,s25[56]};
assign {s53[58],s52[57]} = {1'b0,s27[57]} + {1'b0,s26[57]} + {1'b0,s25[57]};
assign {s53[59],s52[58]} = {1'b0,s27[58]} + {1'b0,s26[58]} + {1'b0,s25[58]};
assign {s53[60],s52[59]} = {1'b0,s27[59]} + {1'b0,s26[59]} + {1'b0,s25[59]};
assign {s53[61],s52[60]} = {1'b0,s27[60]} + {1'b0,s26[60]} + {1'b0,s25[60]};
assign {s53[62],s52[61]} = {1'b0,s27[61]} + {1'b0,s26[61]} + {1'b0,s25[61]};
assign {s53[63],s52[62]} = {1'b0,s27[62]} + {1'b0,s26[62]} + {1'b0,s25[62]};
assign {s53[64],s52[63]} = {1'b0,s27[63]} + {1'b0,s26[63]} + {1'b0,s25[63]};
assign {s53[65],s52[64]} = {1'b0,s27[64]} + {1'b0,s26[64]} + {1'b0,s25[64]};
assign {s53[66],s52[65]} = {1'b0,s27[65]} + {1'b0,s26[65]} + {1'b0,s25[65]};
assign {s53[67],s52[66]} = {1'b0,s27[66]} + {1'b0,s26[66]} + {1'b0,s25[66]};
assign {s55[25],s54[24]} = {1'b0,s28[24]};
assign {s55[26],s54[25]} = {1'b0,s29[25]} + {1'b0,s28[25]};
assign {s55[27],s54[26]} = {1'b0,s30[26]} + {1'b0,s29[26]} + {1'b0,s28[26]};
assign {s55[28],s54[27]} = {1'b0,s30[27]} + {1'b0,s29[27]} + {1'b0,s28[27]};
assign {s55[29],s54[28]} = {1'b0,s30[28]} + {1'b0,s29[28]} + {1'b0,s28[28]};
assign {s55[30],s54[29]} = {1'b0,s30[29]} + {1'b0,s29[29]} + {1'b0,s28[29]};
assign {s55[31],s54[30]} = {1'b0,s30[30]} + {1'b0,s29[30]} + {1'b0,s28[30]};
assign {s55[32],s54[31]} = {1'b0,s30[31]} + {1'b0,s29[31]} + {1'b0,s28[31]};
assign {s55[33],s54[32]} = {1'b0,s30[32]} + {1'b0,s29[32]} + {1'b0,s28[32]};
assign {s55[34],s54[33]} = {1'b0,s30[33]} + {1'b0,s29[33]} + {1'b0,s28[33]};
assign {s55[35],s54[34]} = {1'b0,s30[34]} + {1'b0,s29[34]} + {1'b0,s28[34]};
assign {s55[36],s54[35]} = {1'b0,s30[35]} + {1'b0,s29[35]} + {1'b0,s28[35]};
assign {s55[37],s54[36]} = {1'b0,s30[36]} + {1'b0,s29[36]} + {1'b0,s28[36]};
assign {s55[38],s54[37]} = {1'b0,s30[37]} + {1'b0,s29[37]} + {1'b0,s28[37]};
assign {s55[39],s54[38]} = {1'b0,s30[38]} + {1'b0,s29[38]} + {1'b0,s28[38]};
assign {s55[40],s54[39]} = {1'b0,s30[39]} + {1'b0,s29[39]} + {1'b0,s28[39]};
assign {s55[41],s54[40]} = {1'b0,s30[40]} + {1'b0,s29[40]} + {1'b0,s28[40]};
assign {s55[42],s54[41]} = {1'b0,s30[41]} + {1'b0,s29[41]} + {1'b0,s28[41]};
assign {s55[43],s54[42]} = {1'b0,s30[42]} + {1'b0,s29[42]} + {1'b0,s28[42]};
assign {s55[44],s54[43]} = {1'b0,s30[43]} + {1'b0,s29[43]} + {1'b0,s28[43]};
assign {s55[45],s54[44]} = {1'b0,s30[44]} + {1'b0,s29[44]} + {1'b0,s28[44]};
assign {s55[46],s54[45]} = {1'b0,s30[45]} + {1'b0,s29[45]} + {1'b0,s28[45]};
assign {s55[47],s54[46]} = {1'b0,s30[46]} + {1'b0,s29[46]} + {1'b0,s28[46]};
assign {s55[48],s54[47]} = {1'b0,s30[47]} + {1'b0,s29[47]} + {1'b0,s28[47]};
assign {s55[49],s54[48]} = {1'b0,s30[48]} + {1'b0,s29[48]} + {1'b0,s28[48]};
assign {s55[50],s54[49]} = {1'b0,s30[49]} + {1'b0,s29[49]} + {1'b0,s28[49]};
assign {s55[51],s54[50]} = {1'b0,s30[50]} + {1'b0,s29[50]} + {1'b0,s28[50]};
assign {s55[52],s54[51]} = {1'b0,s30[51]} + {1'b0,s29[51]} + {1'b0,s28[51]};
assign {s55[53],s54[52]} = {1'b0,s30[52]} + {1'b0,s29[52]} + {1'b0,s28[52]};
assign {s55[54],s54[53]} = {1'b0,s30[53]} + {1'b0,s29[53]} + {1'b0,s28[53]};
assign {s55[55],s54[54]} = {1'b0,s30[54]} + {1'b0,s29[54]} + {1'b0,s28[54]};
assign {s55[56],s54[55]} = {1'b0,s30[55]} + {1'b0,s29[55]} + {1'b0,s28[55]};
assign {s55[57],s54[56]} = {1'b0,s30[56]} + {1'b0,s29[56]} + {1'b0,s28[56]};
assign {s55[58],s54[57]} = {1'b0,s30[57]} + {1'b0,s29[57]} + {1'b0,s28[57]};
assign {s55[59],s54[58]} = {1'b0,s30[58]} + {1'b0,s29[58]} + {1'b0,s28[58]};
assign {s55[60],s54[59]} = {1'b0,s30[59]} + {1'b0,s29[59]} + {1'b0,s28[59]};
assign {s55[61],s54[60]} = {1'b0,s30[60]} + {1'b0,s29[60]} + {1'b0,s28[60]};
assign {s55[62],s54[61]} = {1'b0,s30[61]} + {1'b0,s29[61]} + {1'b0,s28[61]};
assign {s55[63],s54[62]} = {1'b0,s30[62]} + {1'b0,s29[62]} + {1'b0,s28[62]};
assign {s55[64],s54[63]} = {1'b0,s30[63]} + {1'b0,s29[63]} + {1'b0,s28[63]};
assign {s55[65],s54[64]} = {1'b0,s30[64]} + {1'b0,s29[64]} + {1'b0,s28[64]};
assign {s55[66],s54[65]} = {1'b0,s30[65]} + {1'b0,s29[65]} + {1'b0,s28[65]};
assign {s55[67],s54[66]} = {1'b0,s30[66]} + {1'b0,s29[66]} + {1'b0,s28[66]};
assign {s57[28],s56[27]} = {1'b0,s31[27]};
assign {s57[29],s56[28]} = {1'b0,s32[28]} + {1'b0,s31[28]};
assign {s57[30],s56[29]} = {1'b0,s33[29]} + {1'b0,s32[29]} + {1'b0,s31[29]};
assign {s57[31],s56[30]} = {1'b0,s33[30]} + {1'b0,s32[30]} + {1'b0,s31[30]};
assign {s57[32],s56[31]} = {1'b0,s33[31]} + {1'b0,s32[31]} + {1'b0,s31[31]};
assign {s57[33],s56[32]} = {1'b0,s33[32]} + {1'b0,s32[32]} + {1'b0,s31[32]};
assign {s57[34],s56[33]} = {1'b0,s33[33]} + {1'b0,s32[33]} + {1'b0,s31[33]};
assign {s57[35],s56[34]} = {1'b0,s33[34]} + {1'b0,s32[34]} + {1'b0,s31[34]};
assign {s57[36],s56[35]} = {1'b0,s33[35]} + {1'b0,s32[35]} + {1'b0,s31[35]};
assign {s57[37],s56[36]} = {1'b0,s33[36]} + {1'b0,s32[36]} + {1'b0,s31[36]};
assign {s57[38],s56[37]} = {1'b0,s33[37]} + {1'b0,s32[37]} + {1'b0,s31[37]};
assign {s57[39],s56[38]} = {1'b0,s33[38]} + {1'b0,s32[38]} + {1'b0,s31[38]};
assign {s57[40],s56[39]} = {1'b0,s33[39]} + {1'b0,s32[39]} + {1'b0,s31[39]};
assign {s57[41],s56[40]} = {1'b0,s33[40]} + {1'b0,s32[40]} + {1'b0,s31[40]};
assign {s57[42],s56[41]} = {1'b0,s33[41]} + {1'b0,s32[41]} + {1'b0,s31[41]};
assign {s57[43],s56[42]} = {1'b0,s33[42]} + {1'b0,s32[42]} + {1'b0,s31[42]};
assign {s57[44],s56[43]} = {1'b0,s33[43]} + {1'b0,s32[43]} + {1'b0,s31[43]};
assign {s57[45],s56[44]} = {1'b0,s33[44]} + {1'b0,s32[44]} + {1'b0,s31[44]};
assign {s57[46],s56[45]} = {1'b0,s33[45]} + {1'b0,s32[45]} + {1'b0,s31[45]};
assign {s57[47],s56[46]} = {1'b0,s33[46]} + {1'b0,s32[46]} + {1'b0,s31[46]};
assign {s57[48],s56[47]} = {1'b0,s33[47]} + {1'b0,s32[47]} + {1'b0,s31[47]};
assign {s57[49],s56[48]} = {1'b0,s33[48]} + {1'b0,s32[48]} + {1'b0,s31[48]};
assign {s57[50],s56[49]} = {1'b0,s33[49]} + {1'b0,s32[49]} + {1'b0,s31[49]};
assign {s57[51],s56[50]} = {1'b0,s33[50]} + {1'b0,s32[50]} + {1'b0,s31[50]};
assign {s57[52],s56[51]} = {1'b0,s33[51]} + {1'b0,s32[51]} + {1'b0,s31[51]};
assign {s57[53],s56[52]} = {1'b0,s33[52]} + {1'b0,s32[52]} + {1'b0,s31[52]};
assign {s57[54],s56[53]} = {1'b0,s33[53]} + {1'b0,s32[53]} + {1'b0,s31[53]};
assign {s57[55],s56[54]} = {1'b0,s33[54]} + {1'b0,s32[54]} + {1'b0,s31[54]};
assign {s57[56],s56[55]} = {1'b0,s33[55]} + {1'b0,s32[55]} + {1'b0,s31[55]};
assign {s57[57],s56[56]} = {1'b0,s33[56]} + {1'b0,s32[56]} + {1'b0,s31[56]};
assign {s57[58],s56[57]} = {1'b0,s33[57]} + {1'b0,s32[57]} + {1'b0,s31[57]};
assign {s57[59],s56[58]} = {1'b0,s33[58]} + {1'b0,s32[58]} + {1'b0,s31[58]};
assign {s57[60],s56[59]} = {1'b0,s33[59]} + {1'b0,s32[59]} + {1'b0,s31[59]};
assign {s57[61],s56[60]} = {1'b0,s33[60]} + {1'b0,s32[60]} + {1'b0,s31[60]};
assign {s57[62],s56[61]} = {1'b0,s33[61]} + {1'b0,s32[61]} + {1'b0,s31[61]};
assign {s57[63],s56[62]} = {1'b0,s33[62]} + {1'b0,s32[62]} + {1'b0,s31[62]};
assign {s57[64],s56[63]} = {1'b0,s33[63]} + {1'b0,s32[63]} + {1'b0,s31[63]};
assign {s57[65],s56[64]} = {1'b0,s33[64]} + {1'b0,s32[64]} + {1'b0,s31[64]};
assign {s57[66],s56[65]} = {1'b0,s33[65]} + {1'b0,s32[65]} + {1'b0,s31[65]};
assign {s57[67],s56[66]} = {1'b0,s33[66]} + {1'b0,s32[66]} + {1'b0,s31[66]};
assign {s59[31],s58[30]} = {1'b0,s34[30]};
assign {s59[32],s58[31]} = {1'b0,s35[31]} + {1'b0,s34[31]};
assign {s59[33],s58[32]} = {1'b0,s36[32]} + {1'b0,s35[32]} + {1'b0,s34[32]};
assign {s59[34],s58[33]} = {1'b0,s36[33]} + {1'b0,s35[33]} + {1'b0,s34[33]};
assign {s59[35],s58[34]} = {1'b0,s36[34]} + {1'b0,s35[34]} + {1'b0,s34[34]};
assign {s59[36],s58[35]} = {1'b0,s36[35]} + {1'b0,s35[35]} + {1'b0,s34[35]};
assign {s59[37],s58[36]} = {1'b0,s36[36]} + {1'b0,s35[36]} + {1'b0,s34[36]};
assign {s59[38],s58[37]} = {1'b0,s36[37]} + {1'b0,s35[37]} + {1'b0,s34[37]};
assign {s59[39],s58[38]} = {1'b0,s36[38]} + {1'b0,s35[38]} + {1'b0,s34[38]};
assign {s59[40],s58[39]} = {1'b0,s36[39]} + {1'b0,s35[39]} + {1'b0,s34[39]};
assign {s59[41],s58[40]} = {1'b0,s36[40]} + {1'b0,s35[40]} + {1'b0,s34[40]};
assign {s59[42],s58[41]} = {1'b0,s36[41]} + {1'b0,s35[41]} + {1'b0,s34[41]};
assign {s59[43],s58[42]} = {1'b0,s36[42]} + {1'b0,s35[42]} + {1'b0,s34[42]};
assign {s59[44],s58[43]} = {1'b0,s36[43]} + {1'b0,s35[43]} + {1'b0,s34[43]};
assign {s59[45],s58[44]} = {1'b0,s36[44]} + {1'b0,s35[44]} + {1'b0,s34[44]};
assign {s59[46],s58[45]} = {1'b0,s36[45]} + {1'b0,s35[45]} + {1'b0,s34[45]};
assign {s59[47],s58[46]} = {1'b0,s36[46]} + {1'b0,s35[46]} + {1'b0,s34[46]};
assign {s59[48],s58[47]} = {1'b0,s36[47]} + {1'b0,s35[47]} + {1'b0,s34[47]};
assign {s59[49],s58[48]} = {1'b0,s36[48]} + {1'b0,s35[48]} + {1'b0,s34[48]};
assign {s59[50],s58[49]} = {1'b0,s36[49]} + {1'b0,s35[49]} + {1'b0,s34[49]};
assign {s59[51],s58[50]} = {1'b0,s36[50]} + {1'b0,s35[50]} + {1'b0,s34[50]};
assign {s59[52],s58[51]} = {1'b0,s36[51]} + {1'b0,s35[51]} + {1'b0,s34[51]};
assign {s59[53],s58[52]} = {1'b0,s36[52]} + {1'b0,s35[52]} + {1'b0,s34[52]};
assign {s59[54],s58[53]} = {1'b0,s36[53]} + {1'b0,s35[53]} + {1'b0,s34[53]};
assign {s59[55],s58[54]} = {1'b0,s36[54]} + {1'b0,s35[54]} + {1'b0,s34[54]};
assign {s59[56],s58[55]} = {1'b0,s36[55]} + {1'b0,s35[55]} + {1'b0,s34[55]};
assign {s59[57],s58[56]} = {1'b0,s36[56]} + {1'b0,s35[56]} + {1'b0,s34[56]};
assign {s59[58],s58[57]} = {1'b0,s36[57]} + {1'b0,s35[57]} + {1'b0,s34[57]};
assign {s59[59],s58[58]} = {1'b0,s36[58]} + {1'b0,s35[58]} + {1'b0,s34[58]};
assign {s59[60],s58[59]} = {1'b0,s36[59]} + {1'b0,s35[59]} + {1'b0,s34[59]};
assign {s59[61],s58[60]} = {1'b0,s36[60]} + {1'b0,s35[60]} + {1'b0,s34[60]};
assign {s59[62],s58[61]} = {1'b0,s36[61]} + {1'b0,s35[61]} + {1'b0,s34[61]};
assign {s59[63],s58[62]} = {1'b0,s36[62]} + {1'b0,s35[62]} + {1'b0,s34[62]};
assign {s59[64],s58[63]} = {1'b0,s36[63]} + {1'b0,s35[63]} + {1'b0,s34[63]};
assign {s59[65],s58[64]} = {1'b0,s36[64]} + {1'b0,s35[64]} + {1'b0,s34[64]};
assign {s59[66],s58[65]} = {1'b0,s36[65]} + {1'b0,s35[65]} + {1'b0,s34[65]};
assign {s59[67],s58[66]} = {1'b0,s36[66]} + {1'b0,s35[66]} + {1'b0,s34[66]};
assign s60 = s37[(PPLEN - 1):32];
assign {s62[1],s61[0]} = {1'b0,s38[0]};
assign {s62[2],s61[1]} = {1'b0,s39[1]} + {1'b0,s38[1]};
assign {s62[3],s61[2]} = {1'b0,s39[2]} + {1'b0,s38[2]};
assign {s62[4],s61[3]} = {1'b0,s40[3]} + {1'b0,s39[3]} + {1'b0,s38[3]};
assign {s62[5],s61[4]} = {1'b0,s40[4]} + {1'b0,s39[4]} + {1'b0,s38[4]};
assign {s62[6],s61[5]} = {1'b0,s40[5]} + {1'b0,s39[5]} + {1'b0,s38[5]};
assign {s62[7],s61[6]} = {1'b0,s40[6]} + {1'b0,s39[6]} + {1'b0,s38[6]};
assign {s62[8],s61[7]} = {1'b0,s40[7]} + {1'b0,s39[7]} + {1'b0,s38[7]};
assign {s62[9],s61[8]} = {1'b0,s40[8]} + {1'b0,s39[8]} + {1'b0,s38[8]};
assign {s62[10],s61[9]} = {1'b0,s40[9]} + {1'b0,s39[9]} + {1'b0,s38[9]};
assign {s62[11],s61[10]} = {1'b0,s40[10]} + {1'b0,s39[10]} + {1'b0,s38[10]};
assign {s62[12],s61[11]} = {1'b0,s40[11]} + {1'b0,s39[11]} + {1'b0,s38[11]};
assign {s62[13],s61[12]} = {1'b0,s40[12]} + {1'b0,s39[12]} + {1'b0,s38[12]};
assign {s62[14],s61[13]} = {1'b0,s40[13]} + {1'b0,s39[13]} + {1'b0,s38[13]};
assign {s62[15],s61[14]} = {1'b0,s40[14]} + {1'b0,s39[14]} + {1'b0,s38[14]};
assign {s62[16],s61[15]} = {1'b0,s40[15]} + {1'b0,s39[15]} + {1'b0,s38[15]};
assign {s62[17],s61[16]} = {1'b0,s40[16]} + {1'b0,s39[16]} + {1'b0,s38[16]};
assign {s62[18],s61[17]} = {1'b0,s40[17]} + {1'b0,s39[17]} + {1'b0,s38[17]};
assign {s62[19],s61[18]} = {1'b0,s40[18]} + {1'b0,s39[18]} + {1'b0,s38[18]};
assign {s62[20],s61[19]} = {1'b0,s40[19]} + {1'b0,s39[19]} + {1'b0,s38[19]};
assign {s62[21],s61[20]} = {1'b0,s40[20]} + {1'b0,s39[20]} + {1'b0,s38[20]};
assign {s62[22],s61[21]} = {1'b0,s40[21]} + {1'b0,s39[21]} + {1'b0,s38[21]};
assign {s62[23],s61[22]} = {1'b0,s40[22]} + {1'b0,s39[22]} + {1'b0,s38[22]};
assign {s62[24],s61[23]} = {1'b0,s40[23]} + {1'b0,s39[23]} + {1'b0,s38[23]};
assign {s62[25],s61[24]} = {1'b0,s40[24]} + {1'b0,s39[24]} + {1'b0,s38[24]};
assign {s62[26],s61[25]} = {1'b0,s40[25]} + {1'b0,s39[25]} + {1'b0,s38[25]};
assign {s62[27],s61[26]} = {1'b0,s40[26]} + {1'b0,s39[26]} + {1'b0,s38[26]};
assign {s62[28],s61[27]} = {1'b0,s40[27]} + {1'b0,s39[27]} + {1'b0,s38[27]};
assign {s62[29],s61[28]} = {1'b0,s40[28]} + {1'b0,s39[28]} + {1'b0,s38[28]};
assign {s62[30],s61[29]} = {1'b0,s40[29]} + {1'b0,s39[29]} + {1'b0,s38[29]};
assign {s62[31],s61[30]} = {1'b0,s40[30]} + {1'b0,s39[30]} + {1'b0,s38[30]};
assign {s62[32],s61[31]} = {1'b0,s40[31]} + {1'b0,s39[31]} + {1'b0,s38[31]};
assign {s62[33],s61[32]} = {1'b0,s40[32]} + {1'b0,s39[32]} + {1'b0,s38[32]};
assign {s62[34],s61[33]} = {1'b0,s40[33]} + {1'b0,s39[33]} + {1'b0,s38[33]};
assign {s62[35],s61[34]} = {1'b0,s40[34]} + {1'b0,s39[34]} + {1'b0,s38[34]};
assign {s62[36],s61[35]} = {1'b0,s40[35]} + {1'b0,s39[35]} + {1'b0,s38[35]};
assign {s62[37],s61[36]} = {1'b0,s40[36]} + {1'b0,s39[36]} + {1'b0,s38[36]};
assign {s62[38],s61[37]} = {1'b0,s40[37]} + {1'b0,s39[37]} + {1'b0,s38[37]};
assign {s62[39],s61[38]} = {1'b0,s40[38]} + {1'b0,s39[38]} + {1'b0,s38[38]};
assign {s62[40],s61[39]} = {1'b0,s40[39]} + {1'b0,s39[39]} + {1'b0,s38[39]};
assign {s62[41],s61[40]} = {1'b0,s40[40]} + {1'b0,s39[40]} + {1'b0,s38[40]};
assign {s62[42],s61[41]} = {1'b0,s40[41]} + {1'b0,s39[41]} + {1'b0,s38[41]};
assign {s62[43],s61[42]} = {1'b0,s40[42]} + {1'b0,s39[42]} + {1'b0,s38[42]};
assign {s62[44],s61[43]} = {1'b0,s40[43]} + {1'b0,s39[43]} + {1'b0,s38[43]};
assign {s62[45],s61[44]} = {1'b0,s40[44]} + {1'b0,s39[44]} + {1'b0,s38[44]};
assign {s62[46],s61[45]} = {1'b0,s40[45]} + {1'b0,s39[45]} + {1'b0,s38[45]};
assign {s62[47],s61[46]} = {1'b0,s40[46]} + {1'b0,s39[46]} + {1'b0,s38[46]};
assign {s62[48],s61[47]} = {1'b0,s40[47]} + {1'b0,s39[47]} + {1'b0,s38[47]};
assign {s62[49],s61[48]} = {1'b0,s40[48]} + {1'b0,s39[48]} + {1'b0,s38[48]};
assign {s62[50],s61[49]} = {1'b0,s40[49]} + {1'b0,s39[49]} + {1'b0,s38[49]};
assign {s62[51],s61[50]} = {1'b0,s40[50]} + {1'b0,s39[50]} + {1'b0,s38[50]};
assign {s62[52],s61[51]} = {1'b0,s40[51]} + {1'b0,s39[51]} + {1'b0,s38[51]};
assign {s62[53],s61[52]} = {1'b0,s40[52]} + {1'b0,s39[52]} + {1'b0,s38[52]};
assign {s62[54],s61[53]} = {1'b0,s40[53]} + {1'b0,s39[53]} + {1'b0,s38[53]};
assign {s62[55],s61[54]} = {1'b0,s40[54]} + {1'b0,s39[54]} + {1'b0,s38[54]};
assign {s62[56],s61[55]} = {1'b0,s40[55]} + {1'b0,s39[55]} + {1'b0,s38[55]};
assign {s62[57],s61[56]} = {1'b0,s40[56]} + {1'b0,s39[56]} + {1'b0,s38[56]};
assign {s62[58],s61[57]} = {1'b0,s40[57]} + {1'b0,s39[57]} + {1'b0,s38[57]};
assign {s62[59],s61[58]} = {1'b0,s40[58]} + {1'b0,s39[58]} + {1'b0,s38[58]};
assign {s62[60],s61[59]} = {1'b0,s40[59]} + {1'b0,s39[59]} + {1'b0,s38[59]};
assign {s62[61],s61[60]} = {1'b0,s40[60]} + {1'b0,s39[60]} + {1'b0,s38[60]};
assign {s62[62],s61[61]} = {1'b0,s40[61]} + {1'b0,s39[61]} + {1'b0,s38[61]};
assign {s62[63],s61[62]} = {1'b0,s40[62]} + {1'b0,s39[62]} + {1'b0,s38[62]};
assign {s62[64],s61[63]} = {1'b0,s40[63]} + {1'b0,s39[63]} + {1'b0,s38[63]};
assign {s62[65],s61[64]} = {1'b0,s40[64]} + {1'b0,s39[64]} + {1'b0,s38[64]};
assign {s62[66],s61[65]} = {1'b0,s40[65]} + {1'b0,s39[65]} + {1'b0,s38[65]};
assign {s62[67],s61[66]} = {1'b0,s40[66]} + {1'b0,s39[66]} + {1'b0,s38[66]};
assign {s64[5],s63[4]} = {1'b0,s41[4]};
assign {s64[6],s63[5]} = {1'b0,s41[5]};
assign {s64[7],s63[6]} = {1'b0,s42[6]} + {1'b0,s41[6]};
assign {s64[8],s63[7]} = {1'b0,s43[7]} + {1'b0,s42[7]} + {1'b0,s41[7]};
assign {s64[9],s63[8]} = {1'b0,s43[8]} + {1'b0,s42[8]} + {1'b0,s41[8]};
assign {s64[10],s63[9]} = {1'b0,s43[9]} + {1'b0,s42[9]} + {1'b0,s41[9]};
assign {s64[11],s63[10]} = {1'b0,s43[10]} + {1'b0,s42[10]} + {1'b0,s41[10]};
assign {s64[12],s63[11]} = {1'b0,s43[11]} + {1'b0,s42[11]} + {1'b0,s41[11]};
assign {s64[13],s63[12]} = {1'b0,s43[12]} + {1'b0,s42[12]} + {1'b0,s41[12]};
assign {s64[14],s63[13]} = {1'b0,s43[13]} + {1'b0,s42[13]} + {1'b0,s41[13]};
assign {s64[15],s63[14]} = {1'b0,s43[14]} + {1'b0,s42[14]} + {1'b0,s41[14]};
assign {s64[16],s63[15]} = {1'b0,s43[15]} + {1'b0,s42[15]} + {1'b0,s41[15]};
assign {s64[17],s63[16]} = {1'b0,s43[16]} + {1'b0,s42[16]} + {1'b0,s41[16]};
assign {s64[18],s63[17]} = {1'b0,s43[17]} + {1'b0,s42[17]} + {1'b0,s41[17]};
assign {s64[19],s63[18]} = {1'b0,s43[18]} + {1'b0,s42[18]} + {1'b0,s41[18]};
assign {s64[20],s63[19]} = {1'b0,s43[19]} + {1'b0,s42[19]} + {1'b0,s41[19]};
assign {s64[21],s63[20]} = {1'b0,s43[20]} + {1'b0,s42[20]} + {1'b0,s41[20]};
assign {s64[22],s63[21]} = {1'b0,s43[21]} + {1'b0,s42[21]} + {1'b0,s41[21]};
assign {s64[23],s63[22]} = {1'b0,s43[22]} + {1'b0,s42[22]} + {1'b0,s41[22]};
assign {s64[24],s63[23]} = {1'b0,s43[23]} + {1'b0,s42[23]} + {1'b0,s41[23]};
assign {s64[25],s63[24]} = {1'b0,s43[24]} + {1'b0,s42[24]} + {1'b0,s41[24]};
assign {s64[26],s63[25]} = {1'b0,s43[25]} + {1'b0,s42[25]} + {1'b0,s41[25]};
assign {s64[27],s63[26]} = {1'b0,s43[26]} + {1'b0,s42[26]} + {1'b0,s41[26]};
assign {s64[28],s63[27]} = {1'b0,s43[27]} + {1'b0,s42[27]} + {1'b0,s41[27]};
assign {s64[29],s63[28]} = {1'b0,s43[28]} + {1'b0,s42[28]} + {1'b0,s41[28]};
assign {s64[30],s63[29]} = {1'b0,s43[29]} + {1'b0,s42[29]} + {1'b0,s41[29]};
assign {s64[31],s63[30]} = {1'b0,s43[30]} + {1'b0,s42[30]} + {1'b0,s41[30]};
assign {s64[32],s63[31]} = {1'b0,s43[31]} + {1'b0,s42[31]} + {1'b0,s41[31]};
assign {s64[33],s63[32]} = {1'b0,s43[32]} + {1'b0,s42[32]} + {1'b0,s41[32]};
assign {s64[34],s63[33]} = {1'b0,s43[33]} + {1'b0,s42[33]} + {1'b0,s41[33]};
assign {s64[35],s63[34]} = {1'b0,s43[34]} + {1'b0,s42[34]} + {1'b0,s41[34]};
assign {s64[36],s63[35]} = {1'b0,s43[35]} + {1'b0,s42[35]} + {1'b0,s41[35]};
assign {s64[37],s63[36]} = {1'b0,s43[36]} + {1'b0,s42[36]} + {1'b0,s41[36]};
assign {s64[38],s63[37]} = {1'b0,s43[37]} + {1'b0,s42[37]} + {1'b0,s41[37]};
assign {s64[39],s63[38]} = {1'b0,s43[38]} + {1'b0,s42[38]} + {1'b0,s41[38]};
assign {s64[40],s63[39]} = {1'b0,s43[39]} + {1'b0,s42[39]} + {1'b0,s41[39]};
assign {s64[41],s63[40]} = {1'b0,s43[40]} + {1'b0,s42[40]} + {1'b0,s41[40]};
assign {s64[42],s63[41]} = {1'b0,s43[41]} + {1'b0,s42[41]} + {1'b0,s41[41]};
assign {s64[43],s63[42]} = {1'b0,s43[42]} + {1'b0,s42[42]} + {1'b0,s41[42]};
assign {s64[44],s63[43]} = {1'b0,s43[43]} + {1'b0,s42[43]} + {1'b0,s41[43]};
assign {s64[45],s63[44]} = {1'b0,s43[44]} + {1'b0,s42[44]} + {1'b0,s41[44]};
assign {s64[46],s63[45]} = {1'b0,s43[45]} + {1'b0,s42[45]} + {1'b0,s41[45]};
assign {s64[47],s63[46]} = {1'b0,s43[46]} + {1'b0,s42[46]} + {1'b0,s41[46]};
assign {s64[48],s63[47]} = {1'b0,s43[47]} + {1'b0,s42[47]} + {1'b0,s41[47]};
assign {s64[49],s63[48]} = {1'b0,s43[48]} + {1'b0,s42[48]} + {1'b0,s41[48]};
assign {s64[50],s63[49]} = {1'b0,s43[49]} + {1'b0,s42[49]} + {1'b0,s41[49]};
assign {s64[51],s63[50]} = {1'b0,s43[50]} + {1'b0,s42[50]} + {1'b0,s41[50]};
assign {s64[52],s63[51]} = {1'b0,s43[51]} + {1'b0,s42[51]} + {1'b0,s41[51]};
assign {s64[53],s63[52]} = {1'b0,s43[52]} + {1'b0,s42[52]} + {1'b0,s41[52]};
assign {s64[54],s63[53]} = {1'b0,s43[53]} + {1'b0,s42[53]} + {1'b0,s41[53]};
assign {s64[55],s63[54]} = {1'b0,s43[54]} + {1'b0,s42[54]} + {1'b0,s41[54]};
assign {s64[56],s63[55]} = {1'b0,s43[55]} + {1'b0,s42[55]} + {1'b0,s41[55]};
assign {s64[57],s63[56]} = {1'b0,s43[56]} + {1'b0,s42[56]} + {1'b0,s41[56]};
assign {s64[58],s63[57]} = {1'b0,s43[57]} + {1'b0,s42[57]} + {1'b0,s41[57]};
assign {s64[59],s63[58]} = {1'b0,s43[58]} + {1'b0,s42[58]} + {1'b0,s41[58]};
assign {s64[60],s63[59]} = {1'b0,s43[59]} + {1'b0,s42[59]} + {1'b0,s41[59]};
assign {s64[61],s63[60]} = {1'b0,s43[60]} + {1'b0,s42[60]} + {1'b0,s41[60]};
assign {s64[62],s63[61]} = {1'b0,s43[61]} + {1'b0,s42[61]} + {1'b0,s41[61]};
assign {s64[63],s63[62]} = {1'b0,s43[62]} + {1'b0,s42[62]} + {1'b0,s41[62]};
assign {s64[64],s63[63]} = {1'b0,s43[63]} + {1'b0,s42[63]} + {1'b0,s41[63]};
assign {s64[65],s63[64]} = {1'b0,s43[64]} + {1'b0,s42[64]} + {1'b0,s41[64]};
assign {s64[66],s63[65]} = {1'b0,s43[65]} + {1'b0,s42[65]} + {1'b0,s41[65]};
assign {s64[67],s63[66]} = {1'b0,s43[66]} + {1'b0,s42[66]} + {1'b0,s41[66]};
assign {s66[10],s65[9]} = {1'b0,s44[9]};
assign {s66[11],s65[10]} = {1'b0,s45[10]} + {1'b0,s44[10]};
assign {s66[12],s65[11]} = {1'b0,s45[11]} + {1'b0,s44[11]};
assign {s66[13],s65[12]} = {1'b0,s46[12]} + {1'b0,s45[12]} + {1'b0,s44[12]};
assign {s66[14],s65[13]} = {1'b0,s46[13]} + {1'b0,s45[13]} + {1'b0,s44[13]};
assign {s66[15],s65[14]} = {1'b0,s46[14]} + {1'b0,s45[14]} + {1'b0,s44[14]};
assign {s66[16],s65[15]} = {1'b0,s46[15]} + {1'b0,s45[15]} + {1'b0,s44[15]};
assign {s66[17],s65[16]} = {1'b0,s46[16]} + {1'b0,s45[16]} + {1'b0,s44[16]};
assign {s66[18],s65[17]} = {1'b0,s46[17]} + {1'b0,s45[17]} + {1'b0,s44[17]};
assign {s66[19],s65[18]} = {1'b0,s46[18]} + {1'b0,s45[18]} + {1'b0,s44[18]};
assign {s66[20],s65[19]} = {1'b0,s46[19]} + {1'b0,s45[19]} + {1'b0,s44[19]};
assign {s66[21],s65[20]} = {1'b0,s46[20]} + {1'b0,s45[20]} + {1'b0,s44[20]};
assign {s66[22],s65[21]} = {1'b0,s46[21]} + {1'b0,s45[21]} + {1'b0,s44[21]};
assign {s66[23],s65[22]} = {1'b0,s46[22]} + {1'b0,s45[22]} + {1'b0,s44[22]};
assign {s66[24],s65[23]} = {1'b0,s46[23]} + {1'b0,s45[23]} + {1'b0,s44[23]};
assign {s66[25],s65[24]} = {1'b0,s46[24]} + {1'b0,s45[24]} + {1'b0,s44[24]};
assign {s66[26],s65[25]} = {1'b0,s46[25]} + {1'b0,s45[25]} + {1'b0,s44[25]};
assign {s66[27],s65[26]} = {1'b0,s46[26]} + {1'b0,s45[26]} + {1'b0,s44[26]};
assign {s66[28],s65[27]} = {1'b0,s46[27]} + {1'b0,s45[27]} + {1'b0,s44[27]};
assign {s66[29],s65[28]} = {1'b0,s46[28]} + {1'b0,s45[28]} + {1'b0,s44[28]};
assign {s66[30],s65[29]} = {1'b0,s46[29]} + {1'b0,s45[29]} + {1'b0,s44[29]};
assign {s66[31],s65[30]} = {1'b0,s46[30]} + {1'b0,s45[30]} + {1'b0,s44[30]};
assign {s66[32],s65[31]} = {1'b0,s46[31]} + {1'b0,s45[31]} + {1'b0,s44[31]};
assign {s66[33],s65[32]} = {1'b0,s46[32]} + {1'b0,s45[32]} + {1'b0,s44[32]};
assign {s66[34],s65[33]} = {1'b0,s46[33]} + {1'b0,s45[33]} + {1'b0,s44[33]};
assign {s66[35],s65[34]} = {1'b0,s46[34]} + {1'b0,s45[34]} + {1'b0,s44[34]};
assign {s66[36],s65[35]} = {1'b0,s46[35]} + {1'b0,s45[35]} + {1'b0,s44[35]};
assign {s66[37],s65[36]} = {1'b0,s46[36]} + {1'b0,s45[36]} + {1'b0,s44[36]};
assign {s66[38],s65[37]} = {1'b0,s46[37]} + {1'b0,s45[37]} + {1'b0,s44[37]};
assign {s66[39],s65[38]} = {1'b0,s46[38]} + {1'b0,s45[38]} + {1'b0,s44[38]};
assign {s66[40],s65[39]} = {1'b0,s46[39]} + {1'b0,s45[39]} + {1'b0,s44[39]};
assign {s66[41],s65[40]} = {1'b0,s46[40]} + {1'b0,s45[40]} + {1'b0,s44[40]};
assign {s66[42],s65[41]} = {1'b0,s46[41]} + {1'b0,s45[41]} + {1'b0,s44[41]};
assign {s66[43],s65[42]} = {1'b0,s46[42]} + {1'b0,s45[42]} + {1'b0,s44[42]};
assign {s66[44],s65[43]} = {1'b0,s46[43]} + {1'b0,s45[43]} + {1'b0,s44[43]};
assign {s66[45],s65[44]} = {1'b0,s46[44]} + {1'b0,s45[44]} + {1'b0,s44[44]};
assign {s66[46],s65[45]} = {1'b0,s46[45]} + {1'b0,s45[45]} + {1'b0,s44[45]};
assign {s66[47],s65[46]} = {1'b0,s46[46]} + {1'b0,s45[46]} + {1'b0,s44[46]};
assign {s66[48],s65[47]} = {1'b0,s46[47]} + {1'b0,s45[47]} + {1'b0,s44[47]};
assign {s66[49],s65[48]} = {1'b0,s46[48]} + {1'b0,s45[48]} + {1'b0,s44[48]};
assign {s66[50],s65[49]} = {1'b0,s46[49]} + {1'b0,s45[49]} + {1'b0,s44[49]};
assign {s66[51],s65[50]} = {1'b0,s46[50]} + {1'b0,s45[50]} + {1'b0,s44[50]};
assign {s66[52],s65[51]} = {1'b0,s46[51]} + {1'b0,s45[51]} + {1'b0,s44[51]};
assign {s66[53],s65[52]} = {1'b0,s46[52]} + {1'b0,s45[52]} + {1'b0,s44[52]};
assign {s66[54],s65[53]} = {1'b0,s46[53]} + {1'b0,s45[53]} + {1'b0,s44[53]};
assign {s66[55],s65[54]} = {1'b0,s46[54]} + {1'b0,s45[54]} + {1'b0,s44[54]};
assign {s66[56],s65[55]} = {1'b0,s46[55]} + {1'b0,s45[55]} + {1'b0,s44[55]};
assign {s66[57],s65[56]} = {1'b0,s46[56]} + {1'b0,s45[56]} + {1'b0,s44[56]};
assign {s66[58],s65[57]} = {1'b0,s46[57]} + {1'b0,s45[57]} + {1'b0,s44[57]};
assign {s66[59],s65[58]} = {1'b0,s46[58]} + {1'b0,s45[58]} + {1'b0,s44[58]};
assign {s66[60],s65[59]} = {1'b0,s46[59]} + {1'b0,s45[59]} + {1'b0,s44[59]};
assign {s66[61],s65[60]} = {1'b0,s46[60]} + {1'b0,s45[60]} + {1'b0,s44[60]};
assign {s66[62],s65[61]} = {1'b0,s46[61]} + {1'b0,s45[61]} + {1'b0,s44[61]};
assign {s66[63],s65[62]} = {1'b0,s46[62]} + {1'b0,s45[62]} + {1'b0,s44[62]};
assign {s66[64],s65[63]} = {1'b0,s46[63]} + {1'b0,s45[63]} + {1'b0,s44[63]};
assign {s66[65],s65[64]} = {1'b0,s46[64]} + {1'b0,s45[64]} + {1'b0,s44[64]};
assign {s66[66],s65[65]} = {1'b0,s46[65]} + {1'b0,s45[65]} + {1'b0,s44[65]};
assign {s66[67],s65[66]} = {1'b0,s46[66]} + {1'b0,s45[66]} + {1'b0,s44[66]};
assign {s68[14],s67[13]} = {1'b0,s47[13]};
assign {s68[15],s67[14]} = {1'b0,s47[14]};
assign {s68[16],s67[15]} = {1'b0,s48[15]} + {1'b0,s47[15]};
assign {s68[17],s67[16]} = {1'b0,s49[16]} + {1'b0,s48[16]} + {1'b0,s47[16]};
assign {s68[18],s67[17]} = {1'b0,s49[17]} + {1'b0,s48[17]} + {1'b0,s47[17]};
assign {s68[19],s67[18]} = {1'b0,s49[18]} + {1'b0,s48[18]} + {1'b0,s47[18]};
assign {s68[20],s67[19]} = {1'b0,s49[19]} + {1'b0,s48[19]} + {1'b0,s47[19]};
assign {s68[21],s67[20]} = {1'b0,s49[20]} + {1'b0,s48[20]} + {1'b0,s47[20]};
assign {s68[22],s67[21]} = {1'b0,s49[21]} + {1'b0,s48[21]} + {1'b0,s47[21]};
assign {s68[23],s67[22]} = {1'b0,s49[22]} + {1'b0,s48[22]} + {1'b0,s47[22]};
assign {s68[24],s67[23]} = {1'b0,s49[23]} + {1'b0,s48[23]} + {1'b0,s47[23]};
assign {s68[25],s67[24]} = {1'b0,s49[24]} + {1'b0,s48[24]} + {1'b0,s47[24]};
assign {s68[26],s67[25]} = {1'b0,s49[25]} + {1'b0,s48[25]} + {1'b0,s47[25]};
assign {s68[27],s67[26]} = {1'b0,s49[26]} + {1'b0,s48[26]} + {1'b0,s47[26]};
assign {s68[28],s67[27]} = {1'b0,s49[27]} + {1'b0,s48[27]} + {1'b0,s47[27]};
assign {s68[29],s67[28]} = {1'b0,s49[28]} + {1'b0,s48[28]} + {1'b0,s47[28]};
assign {s68[30],s67[29]} = {1'b0,s49[29]} + {1'b0,s48[29]} + {1'b0,s47[29]};
assign {s68[31],s67[30]} = {1'b0,s49[30]} + {1'b0,s48[30]} + {1'b0,s47[30]};
assign {s68[32],s67[31]} = {1'b0,s49[31]} + {1'b0,s48[31]} + {1'b0,s47[31]};
assign {s68[33],s67[32]} = {1'b0,s49[32]} + {1'b0,s48[32]} + {1'b0,s47[32]};
assign {s68[34],s67[33]} = {1'b0,s49[33]} + {1'b0,s48[33]} + {1'b0,s47[33]};
assign {s68[35],s67[34]} = {1'b0,s49[34]} + {1'b0,s48[34]} + {1'b0,s47[34]};
assign {s68[36],s67[35]} = {1'b0,s49[35]} + {1'b0,s48[35]} + {1'b0,s47[35]};
assign {s68[37],s67[36]} = {1'b0,s49[36]} + {1'b0,s48[36]} + {1'b0,s47[36]};
assign {s68[38],s67[37]} = {1'b0,s49[37]} + {1'b0,s48[37]} + {1'b0,s47[37]};
assign {s68[39],s67[38]} = {1'b0,s49[38]} + {1'b0,s48[38]} + {1'b0,s47[38]};
assign {s68[40],s67[39]} = {1'b0,s49[39]} + {1'b0,s48[39]} + {1'b0,s47[39]};
assign {s68[41],s67[40]} = {1'b0,s49[40]} + {1'b0,s48[40]} + {1'b0,s47[40]};
assign {s68[42],s67[41]} = {1'b0,s49[41]} + {1'b0,s48[41]} + {1'b0,s47[41]};
assign {s68[43],s67[42]} = {1'b0,s49[42]} + {1'b0,s48[42]} + {1'b0,s47[42]};
assign {s68[44],s67[43]} = {1'b0,s49[43]} + {1'b0,s48[43]} + {1'b0,s47[43]};
assign {s68[45],s67[44]} = {1'b0,s49[44]} + {1'b0,s48[44]} + {1'b0,s47[44]};
assign {s68[46],s67[45]} = {1'b0,s49[45]} + {1'b0,s48[45]} + {1'b0,s47[45]};
assign {s68[47],s67[46]} = {1'b0,s49[46]} + {1'b0,s48[46]} + {1'b0,s47[46]};
assign {s68[48],s67[47]} = {1'b0,s49[47]} + {1'b0,s48[47]} + {1'b0,s47[47]};
assign {s68[49],s67[48]} = {1'b0,s49[48]} + {1'b0,s48[48]} + {1'b0,s47[48]};
assign {s68[50],s67[49]} = {1'b0,s49[49]} + {1'b0,s48[49]} + {1'b0,s47[49]};
assign {s68[51],s67[50]} = {1'b0,s49[50]} + {1'b0,s48[50]} + {1'b0,s47[50]};
assign {s68[52],s67[51]} = {1'b0,s49[51]} + {1'b0,s48[51]} + {1'b0,s47[51]};
assign {s68[53],s67[52]} = {1'b0,s49[52]} + {1'b0,s48[52]} + {1'b0,s47[52]};
assign {s68[54],s67[53]} = {1'b0,s49[53]} + {1'b0,s48[53]} + {1'b0,s47[53]};
assign {s68[55],s67[54]} = {1'b0,s49[54]} + {1'b0,s48[54]} + {1'b0,s47[54]};
assign {s68[56],s67[55]} = {1'b0,s49[55]} + {1'b0,s48[55]} + {1'b0,s47[55]};
assign {s68[57],s67[56]} = {1'b0,s49[56]} + {1'b0,s48[56]} + {1'b0,s47[56]};
assign {s68[58],s67[57]} = {1'b0,s49[57]} + {1'b0,s48[57]} + {1'b0,s47[57]};
assign {s68[59],s67[58]} = {1'b0,s49[58]} + {1'b0,s48[58]} + {1'b0,s47[58]};
assign {s68[60],s67[59]} = {1'b0,s49[59]} + {1'b0,s48[59]} + {1'b0,s47[59]};
assign {s68[61],s67[60]} = {1'b0,s49[60]} + {1'b0,s48[60]} + {1'b0,s47[60]};
assign {s68[62],s67[61]} = {1'b0,s49[61]} + {1'b0,s48[61]} + {1'b0,s47[61]};
assign {s68[63],s67[62]} = {1'b0,s49[62]} + {1'b0,s48[62]} + {1'b0,s47[62]};
assign {s68[64],s67[63]} = {1'b0,s49[63]} + {1'b0,s48[63]} + {1'b0,s47[63]};
assign {s68[65],s67[64]} = {1'b0,s49[64]} + {1'b0,s48[64]} + {1'b0,s47[64]};
assign {s68[66],s67[65]} = {1'b0,s49[65]} + {1'b0,s48[65]} + {1'b0,s47[65]};
assign {s68[67],s67[66]} = {1'b0,s49[66]} + {1'b0,s48[66]} + {1'b0,s47[66]};
assign {s70[19],s69[18]} = {1'b0,s50[18]};
assign {s70[20],s69[19]} = {1'b0,s51[19]} + {1'b0,s50[19]};
assign {s70[21],s69[20]} = {1'b0,s51[20]} + {1'b0,s50[20]};
assign {s70[22],s69[21]} = {1'b0,s52[21]} + {1'b0,s51[21]} + {1'b0,s50[21]};
assign {s70[23],s69[22]} = {1'b0,s52[22]} + {1'b0,s51[22]} + {1'b0,s50[22]};
assign {s70[24],s69[23]} = {1'b0,s52[23]} + {1'b0,s51[23]} + {1'b0,s50[23]};
assign {s70[25],s69[24]} = {1'b0,s52[24]} + {1'b0,s51[24]} + {1'b0,s50[24]};
assign {s70[26],s69[25]} = {1'b0,s52[25]} + {1'b0,s51[25]} + {1'b0,s50[25]};
assign {s70[27],s69[26]} = {1'b0,s52[26]} + {1'b0,s51[26]} + {1'b0,s50[26]};
assign {s70[28],s69[27]} = {1'b0,s52[27]} + {1'b0,s51[27]} + {1'b0,s50[27]};
assign {s70[29],s69[28]} = {1'b0,s52[28]} + {1'b0,s51[28]} + {1'b0,s50[28]};
assign {s70[30],s69[29]} = {1'b0,s52[29]} + {1'b0,s51[29]} + {1'b0,s50[29]};
assign {s70[31],s69[30]} = {1'b0,s52[30]} + {1'b0,s51[30]} + {1'b0,s50[30]};
assign {s70[32],s69[31]} = {1'b0,s52[31]} + {1'b0,s51[31]} + {1'b0,s50[31]};
assign {s70[33],s69[32]} = {1'b0,s52[32]} + {1'b0,s51[32]} + {1'b0,s50[32]};
assign {s70[34],s69[33]} = {1'b0,s52[33]} + {1'b0,s51[33]} + {1'b0,s50[33]};
assign {s70[35],s69[34]} = {1'b0,s52[34]} + {1'b0,s51[34]} + {1'b0,s50[34]};
assign {s70[36],s69[35]} = {1'b0,s52[35]} + {1'b0,s51[35]} + {1'b0,s50[35]};
assign {s70[37],s69[36]} = {1'b0,s52[36]} + {1'b0,s51[36]} + {1'b0,s50[36]};
assign {s70[38],s69[37]} = {1'b0,s52[37]} + {1'b0,s51[37]} + {1'b0,s50[37]};
assign {s70[39],s69[38]} = {1'b0,s52[38]} + {1'b0,s51[38]} + {1'b0,s50[38]};
assign {s70[40],s69[39]} = {1'b0,s52[39]} + {1'b0,s51[39]} + {1'b0,s50[39]};
assign {s70[41],s69[40]} = {1'b0,s52[40]} + {1'b0,s51[40]} + {1'b0,s50[40]};
assign {s70[42],s69[41]} = {1'b0,s52[41]} + {1'b0,s51[41]} + {1'b0,s50[41]};
assign {s70[43],s69[42]} = {1'b0,s52[42]} + {1'b0,s51[42]} + {1'b0,s50[42]};
assign {s70[44],s69[43]} = {1'b0,s52[43]} + {1'b0,s51[43]} + {1'b0,s50[43]};
assign {s70[45],s69[44]} = {1'b0,s52[44]} + {1'b0,s51[44]} + {1'b0,s50[44]};
assign {s70[46],s69[45]} = {1'b0,s52[45]} + {1'b0,s51[45]} + {1'b0,s50[45]};
assign {s70[47],s69[46]} = {1'b0,s52[46]} + {1'b0,s51[46]} + {1'b0,s50[46]};
assign {s70[48],s69[47]} = {1'b0,s52[47]} + {1'b0,s51[47]} + {1'b0,s50[47]};
assign {s70[49],s69[48]} = {1'b0,s52[48]} + {1'b0,s51[48]} + {1'b0,s50[48]};
assign {s70[50],s69[49]} = {1'b0,s52[49]} + {1'b0,s51[49]} + {1'b0,s50[49]};
assign {s70[51],s69[50]} = {1'b0,s52[50]} + {1'b0,s51[50]} + {1'b0,s50[50]};
assign {s70[52],s69[51]} = {1'b0,s52[51]} + {1'b0,s51[51]} + {1'b0,s50[51]};
assign {s70[53],s69[52]} = {1'b0,s52[52]} + {1'b0,s51[52]} + {1'b0,s50[52]};
assign {s70[54],s69[53]} = {1'b0,s52[53]} + {1'b0,s51[53]} + {1'b0,s50[53]};
assign {s70[55],s69[54]} = {1'b0,s52[54]} + {1'b0,s51[54]} + {1'b0,s50[54]};
assign {s70[56],s69[55]} = {1'b0,s52[55]} + {1'b0,s51[55]} + {1'b0,s50[55]};
assign {s70[57],s69[56]} = {1'b0,s52[56]} + {1'b0,s51[56]} + {1'b0,s50[56]};
assign {s70[58],s69[57]} = {1'b0,s52[57]} + {1'b0,s51[57]} + {1'b0,s50[57]};
assign {s70[59],s69[58]} = {1'b0,s52[58]} + {1'b0,s51[58]} + {1'b0,s50[58]};
assign {s70[60],s69[59]} = {1'b0,s52[59]} + {1'b0,s51[59]} + {1'b0,s50[59]};
assign {s70[61],s69[60]} = {1'b0,s52[60]} + {1'b0,s51[60]} + {1'b0,s50[60]};
assign {s70[62],s69[61]} = {1'b0,s52[61]} + {1'b0,s51[61]} + {1'b0,s50[61]};
assign {s70[63],s69[62]} = {1'b0,s52[62]} + {1'b0,s51[62]} + {1'b0,s50[62]};
assign {s70[64],s69[63]} = {1'b0,s52[63]} + {1'b0,s51[63]} + {1'b0,s50[63]};
assign {s70[65],s69[64]} = {1'b0,s52[64]} + {1'b0,s51[64]} + {1'b0,s50[64]};
assign {s70[66],s69[65]} = {1'b0,s52[65]} + {1'b0,s51[65]} + {1'b0,s50[65]};
assign {s70[67],s69[66]} = {1'b0,s52[66]} + {1'b0,s51[66]} + {1'b0,s50[66]};
assign {s72[23],s71[22]} = {1'b0,s53[22]};
assign {s72[24],s71[23]} = {1'b0,s53[23]};
assign {s72[25],s71[24]} = {1'b0,s54[24]} + {1'b0,s53[24]};
assign {s72[26],s71[25]} = {1'b0,s55[25]} + {1'b0,s54[25]} + {1'b0,s53[25]};
assign {s72[27],s71[26]} = {1'b0,s55[26]} + {1'b0,s54[26]} + {1'b0,s53[26]};
assign {s72[28],s71[27]} = {1'b0,s55[27]} + {1'b0,s54[27]} + {1'b0,s53[27]};
assign {s72[29],s71[28]} = {1'b0,s55[28]} + {1'b0,s54[28]} + {1'b0,s53[28]};
assign {s72[30],s71[29]} = {1'b0,s55[29]} + {1'b0,s54[29]} + {1'b0,s53[29]};
assign {s72[31],s71[30]} = {1'b0,s55[30]} + {1'b0,s54[30]} + {1'b0,s53[30]};
assign {s72[32],s71[31]} = {1'b0,s55[31]} + {1'b0,s54[31]} + {1'b0,s53[31]};
assign {s72[33],s71[32]} = {1'b0,s55[32]} + {1'b0,s54[32]} + {1'b0,s53[32]};
assign {s72[34],s71[33]} = {1'b0,s55[33]} + {1'b0,s54[33]} + {1'b0,s53[33]};
assign {s72[35],s71[34]} = {1'b0,s55[34]} + {1'b0,s54[34]} + {1'b0,s53[34]};
assign {s72[36],s71[35]} = {1'b0,s55[35]} + {1'b0,s54[35]} + {1'b0,s53[35]};
assign {s72[37],s71[36]} = {1'b0,s55[36]} + {1'b0,s54[36]} + {1'b0,s53[36]};
assign {s72[38],s71[37]} = {1'b0,s55[37]} + {1'b0,s54[37]} + {1'b0,s53[37]};
assign {s72[39],s71[38]} = {1'b0,s55[38]} + {1'b0,s54[38]} + {1'b0,s53[38]};
assign {s72[40],s71[39]} = {1'b0,s55[39]} + {1'b0,s54[39]} + {1'b0,s53[39]};
assign {s72[41],s71[40]} = {1'b0,s55[40]} + {1'b0,s54[40]} + {1'b0,s53[40]};
assign {s72[42],s71[41]} = {1'b0,s55[41]} + {1'b0,s54[41]} + {1'b0,s53[41]};
assign {s72[43],s71[42]} = {1'b0,s55[42]} + {1'b0,s54[42]} + {1'b0,s53[42]};
assign {s72[44],s71[43]} = {1'b0,s55[43]} + {1'b0,s54[43]} + {1'b0,s53[43]};
assign {s72[45],s71[44]} = {1'b0,s55[44]} + {1'b0,s54[44]} + {1'b0,s53[44]};
assign {s72[46],s71[45]} = {1'b0,s55[45]} + {1'b0,s54[45]} + {1'b0,s53[45]};
assign {s72[47],s71[46]} = {1'b0,s55[46]} + {1'b0,s54[46]} + {1'b0,s53[46]};
assign {s72[48],s71[47]} = {1'b0,s55[47]} + {1'b0,s54[47]} + {1'b0,s53[47]};
assign {s72[49],s71[48]} = {1'b0,s55[48]} + {1'b0,s54[48]} + {1'b0,s53[48]};
assign {s72[50],s71[49]} = {1'b0,s55[49]} + {1'b0,s54[49]} + {1'b0,s53[49]};
assign {s72[51],s71[50]} = {1'b0,s55[50]} + {1'b0,s54[50]} + {1'b0,s53[50]};
assign {s72[52],s71[51]} = {1'b0,s55[51]} + {1'b0,s54[51]} + {1'b0,s53[51]};
assign {s72[53],s71[52]} = {1'b0,s55[52]} + {1'b0,s54[52]} + {1'b0,s53[52]};
assign {s72[54],s71[53]} = {1'b0,s55[53]} + {1'b0,s54[53]} + {1'b0,s53[53]};
assign {s72[55],s71[54]} = {1'b0,s55[54]} + {1'b0,s54[54]} + {1'b0,s53[54]};
assign {s72[56],s71[55]} = {1'b0,s55[55]} + {1'b0,s54[55]} + {1'b0,s53[55]};
assign {s72[57],s71[56]} = {1'b0,s55[56]} + {1'b0,s54[56]} + {1'b0,s53[56]};
assign {s72[58],s71[57]} = {1'b0,s55[57]} + {1'b0,s54[57]} + {1'b0,s53[57]};
assign {s72[59],s71[58]} = {1'b0,s55[58]} + {1'b0,s54[58]} + {1'b0,s53[58]};
assign {s72[60],s71[59]} = {1'b0,s55[59]} + {1'b0,s54[59]} + {1'b0,s53[59]};
assign {s72[61],s71[60]} = {1'b0,s55[60]} + {1'b0,s54[60]} + {1'b0,s53[60]};
assign {s72[62],s71[61]} = {1'b0,s55[61]} + {1'b0,s54[61]} + {1'b0,s53[61]};
assign {s72[63],s71[62]} = {1'b0,s55[62]} + {1'b0,s54[62]} + {1'b0,s53[62]};
assign {s72[64],s71[63]} = {1'b0,s55[63]} + {1'b0,s54[63]} + {1'b0,s53[63]};
assign {s72[65],s71[64]} = {1'b0,s55[64]} + {1'b0,s54[64]} + {1'b0,s53[64]};
assign {s72[66],s71[65]} = {1'b0,s55[65]} + {1'b0,s54[65]} + {1'b0,s53[65]};
assign {s72[67],s71[66]} = {1'b0,s55[66]} + {1'b0,s54[66]} + {1'b0,s53[66]};
assign {s74[28],s73[27]} = {1'b0,s56[27]};
assign {s74[29],s73[28]} = {1'b0,s57[28]} + {1'b0,s56[28]};
assign {s74[30],s73[29]} = {1'b0,s57[29]} + {1'b0,s56[29]};
assign {s74[31],s73[30]} = {1'b0,s58[30]} + {1'b0,s57[30]} + {1'b0,s56[30]};
assign {s74[32],s73[31]} = {1'b0,s58[31]} + {1'b0,s57[31]} + {1'b0,s56[31]};
assign {s74[33],s73[32]} = {1'b0,s58[32]} + {1'b0,s57[32]} + {1'b0,s56[32]};
assign {s74[34],s73[33]} = {1'b0,s58[33]} + {1'b0,s57[33]} + {1'b0,s56[33]};
assign {s74[35],s73[34]} = {1'b0,s58[34]} + {1'b0,s57[34]} + {1'b0,s56[34]};
assign {s74[36],s73[35]} = {1'b0,s58[35]} + {1'b0,s57[35]} + {1'b0,s56[35]};
assign {s74[37],s73[36]} = {1'b0,s58[36]} + {1'b0,s57[36]} + {1'b0,s56[36]};
assign {s74[38],s73[37]} = {1'b0,s58[37]} + {1'b0,s57[37]} + {1'b0,s56[37]};
assign {s74[39],s73[38]} = {1'b0,s58[38]} + {1'b0,s57[38]} + {1'b0,s56[38]};
assign {s74[40],s73[39]} = {1'b0,s58[39]} + {1'b0,s57[39]} + {1'b0,s56[39]};
assign {s74[41],s73[40]} = {1'b0,s58[40]} + {1'b0,s57[40]} + {1'b0,s56[40]};
assign {s74[42],s73[41]} = {1'b0,s58[41]} + {1'b0,s57[41]} + {1'b0,s56[41]};
assign {s74[43],s73[42]} = {1'b0,s58[42]} + {1'b0,s57[42]} + {1'b0,s56[42]};
assign {s74[44],s73[43]} = {1'b0,s58[43]} + {1'b0,s57[43]} + {1'b0,s56[43]};
assign {s74[45],s73[44]} = {1'b0,s58[44]} + {1'b0,s57[44]} + {1'b0,s56[44]};
assign {s74[46],s73[45]} = {1'b0,s58[45]} + {1'b0,s57[45]} + {1'b0,s56[45]};
assign {s74[47],s73[46]} = {1'b0,s58[46]} + {1'b0,s57[46]} + {1'b0,s56[46]};
assign {s74[48],s73[47]} = {1'b0,s58[47]} + {1'b0,s57[47]} + {1'b0,s56[47]};
assign {s74[49],s73[48]} = {1'b0,s58[48]} + {1'b0,s57[48]} + {1'b0,s56[48]};
assign {s74[50],s73[49]} = {1'b0,s58[49]} + {1'b0,s57[49]} + {1'b0,s56[49]};
assign {s74[51],s73[50]} = {1'b0,s58[50]} + {1'b0,s57[50]} + {1'b0,s56[50]};
assign {s74[52],s73[51]} = {1'b0,s58[51]} + {1'b0,s57[51]} + {1'b0,s56[51]};
assign {s74[53],s73[52]} = {1'b0,s58[52]} + {1'b0,s57[52]} + {1'b0,s56[52]};
assign {s74[54],s73[53]} = {1'b0,s58[53]} + {1'b0,s57[53]} + {1'b0,s56[53]};
assign {s74[55],s73[54]} = {1'b0,s58[54]} + {1'b0,s57[54]} + {1'b0,s56[54]};
assign {s74[56],s73[55]} = {1'b0,s58[55]} + {1'b0,s57[55]} + {1'b0,s56[55]};
assign {s74[57],s73[56]} = {1'b0,s58[56]} + {1'b0,s57[56]} + {1'b0,s56[56]};
assign {s74[58],s73[57]} = {1'b0,s58[57]} + {1'b0,s57[57]} + {1'b0,s56[57]};
assign {s74[59],s73[58]} = {1'b0,s58[58]} + {1'b0,s57[58]} + {1'b0,s56[58]};
assign {s74[60],s73[59]} = {1'b0,s58[59]} + {1'b0,s57[59]} + {1'b0,s56[59]};
assign {s74[61],s73[60]} = {1'b0,s58[60]} + {1'b0,s57[60]} + {1'b0,s56[60]};
assign {s74[62],s73[61]} = {1'b0,s58[61]} + {1'b0,s57[61]} + {1'b0,s56[61]};
assign {s74[63],s73[62]} = {1'b0,s58[62]} + {1'b0,s57[62]} + {1'b0,s56[62]};
assign {s74[64],s73[63]} = {1'b0,s58[63]} + {1'b0,s57[63]} + {1'b0,s56[63]};
assign {s74[65],s73[64]} = {1'b0,s58[64]} + {1'b0,s57[64]} + {1'b0,s56[64]};
assign {s74[66],s73[65]} = {1'b0,s58[65]} + {1'b0,s57[65]} + {1'b0,s56[65]};
assign {s74[67],s73[66]} = {1'b0,s58[66]} + {1'b0,s57[66]} + {1'b0,s56[66]};
assign s75 = s59[(PPLEN - 1):31];
assign s76 = s60[(PPLEN - 1):32];
assign {s78[1],s77[0]} = {1'b0,s61[0]};
assign {s78[2],s77[1]} = {1'b0,s62[1]} + {1'b0,s61[1]};
assign {s78[3],s77[2]} = {1'b0,s62[2]} + {1'b0,s61[2]};
assign {s78[4],s77[3]} = {1'b0,s62[3]} + {1'b0,s61[3]};
assign {s78[5],s77[4]} = {1'b0,s63[4]} + {1'b0,s62[4]} + {1'b0,s61[4]};
assign {s78[6],s77[5]} = {1'b0,s63[5]} + {1'b0,s62[5]} + {1'b0,s61[5]};
assign {s78[7],s77[6]} = {1'b0,s63[6]} + {1'b0,s62[6]} + {1'b0,s61[6]};
assign {s78[8],s77[7]} = {1'b0,s63[7]} + {1'b0,s62[7]} + {1'b0,s61[7]};
assign {s78[9],s77[8]} = {1'b0,s63[8]} + {1'b0,s62[8]} + {1'b0,s61[8]};
assign {s78[10],s77[9]} = {1'b0,s63[9]} + {1'b0,s62[9]} + {1'b0,s61[9]};
assign {s78[11],s77[10]} = {1'b0,s63[10]} + {1'b0,s62[10]} + {1'b0,s61[10]};
assign {s78[12],s77[11]} = {1'b0,s63[11]} + {1'b0,s62[11]} + {1'b0,s61[11]};
assign {s78[13],s77[12]} = {1'b0,s63[12]} + {1'b0,s62[12]} + {1'b0,s61[12]};
assign {s78[14],s77[13]} = {1'b0,s63[13]} + {1'b0,s62[13]} + {1'b0,s61[13]};
assign {s78[15],s77[14]} = {1'b0,s63[14]} + {1'b0,s62[14]} + {1'b0,s61[14]};
assign {s78[16],s77[15]} = {1'b0,s63[15]} + {1'b0,s62[15]} + {1'b0,s61[15]};
assign {s78[17],s77[16]} = {1'b0,s63[16]} + {1'b0,s62[16]} + {1'b0,s61[16]};
assign {s78[18],s77[17]} = {1'b0,s63[17]} + {1'b0,s62[17]} + {1'b0,s61[17]};
assign {s78[19],s77[18]} = {1'b0,s63[18]} + {1'b0,s62[18]} + {1'b0,s61[18]};
assign {s78[20],s77[19]} = {1'b0,s63[19]} + {1'b0,s62[19]} + {1'b0,s61[19]};
assign {s78[21],s77[20]} = {1'b0,s63[20]} + {1'b0,s62[20]} + {1'b0,s61[20]};
assign {s78[22],s77[21]} = {1'b0,s63[21]} + {1'b0,s62[21]} + {1'b0,s61[21]};
assign {s78[23],s77[22]} = {1'b0,s63[22]} + {1'b0,s62[22]} + {1'b0,s61[22]};
assign {s78[24],s77[23]} = {1'b0,s63[23]} + {1'b0,s62[23]} + {1'b0,s61[23]};
assign {s78[25],s77[24]} = {1'b0,s63[24]} + {1'b0,s62[24]} + {1'b0,s61[24]};
assign {s78[26],s77[25]} = {1'b0,s63[25]} + {1'b0,s62[25]} + {1'b0,s61[25]};
assign {s78[27],s77[26]} = {1'b0,s63[26]} + {1'b0,s62[26]} + {1'b0,s61[26]};
assign {s78[28],s77[27]} = {1'b0,s63[27]} + {1'b0,s62[27]} + {1'b0,s61[27]};
assign {s78[29],s77[28]} = {1'b0,s63[28]} + {1'b0,s62[28]} + {1'b0,s61[28]};
assign {s78[30],s77[29]} = {1'b0,s63[29]} + {1'b0,s62[29]} + {1'b0,s61[29]};
assign {s78[31],s77[30]} = {1'b0,s63[30]} + {1'b0,s62[30]} + {1'b0,s61[30]};
assign {s78[32],s77[31]} = {1'b0,s63[31]} + {1'b0,s62[31]} + {1'b0,s61[31]};
assign {s78[33],s77[32]} = {1'b0,s63[32]} + {1'b0,s62[32]} + {1'b0,s61[32]};
assign {s78[34],s77[33]} = {1'b0,s63[33]} + {1'b0,s62[33]} + {1'b0,s61[33]};
assign {s78[35],s77[34]} = {1'b0,s63[34]} + {1'b0,s62[34]} + {1'b0,s61[34]};
assign {s78[36],s77[35]} = {1'b0,s63[35]} + {1'b0,s62[35]} + {1'b0,s61[35]};
assign {s78[37],s77[36]} = {1'b0,s63[36]} + {1'b0,s62[36]} + {1'b0,s61[36]};
assign {s78[38],s77[37]} = {1'b0,s63[37]} + {1'b0,s62[37]} + {1'b0,s61[37]};
assign {s78[39],s77[38]} = {1'b0,s63[38]} + {1'b0,s62[38]} + {1'b0,s61[38]};
assign {s78[40],s77[39]} = {1'b0,s63[39]} + {1'b0,s62[39]} + {1'b0,s61[39]};
assign {s78[41],s77[40]} = {1'b0,s63[40]} + {1'b0,s62[40]} + {1'b0,s61[40]};
assign {s78[42],s77[41]} = {1'b0,s63[41]} + {1'b0,s62[41]} + {1'b0,s61[41]};
assign {s78[43],s77[42]} = {1'b0,s63[42]} + {1'b0,s62[42]} + {1'b0,s61[42]};
assign {s78[44],s77[43]} = {1'b0,s63[43]} + {1'b0,s62[43]} + {1'b0,s61[43]};
assign {s78[45],s77[44]} = {1'b0,s63[44]} + {1'b0,s62[44]} + {1'b0,s61[44]};
assign {s78[46],s77[45]} = {1'b0,s63[45]} + {1'b0,s62[45]} + {1'b0,s61[45]};
assign {s78[47],s77[46]} = {1'b0,s63[46]} + {1'b0,s62[46]} + {1'b0,s61[46]};
assign {s78[48],s77[47]} = {1'b0,s63[47]} + {1'b0,s62[47]} + {1'b0,s61[47]};
assign {s78[49],s77[48]} = {1'b0,s63[48]} + {1'b0,s62[48]} + {1'b0,s61[48]};
assign {s78[50],s77[49]} = {1'b0,s63[49]} + {1'b0,s62[49]} + {1'b0,s61[49]};
assign {s78[51],s77[50]} = {1'b0,s63[50]} + {1'b0,s62[50]} + {1'b0,s61[50]};
assign {s78[52],s77[51]} = {1'b0,s63[51]} + {1'b0,s62[51]} + {1'b0,s61[51]};
assign {s78[53],s77[52]} = {1'b0,s63[52]} + {1'b0,s62[52]} + {1'b0,s61[52]};
assign {s78[54],s77[53]} = {1'b0,s63[53]} + {1'b0,s62[53]} + {1'b0,s61[53]};
assign {s78[55],s77[54]} = {1'b0,s63[54]} + {1'b0,s62[54]} + {1'b0,s61[54]};
assign {s78[56],s77[55]} = {1'b0,s63[55]} + {1'b0,s62[55]} + {1'b0,s61[55]};
assign {s78[57],s77[56]} = {1'b0,s63[56]} + {1'b0,s62[56]} + {1'b0,s61[56]};
assign {s78[58],s77[57]} = {1'b0,s63[57]} + {1'b0,s62[57]} + {1'b0,s61[57]};
assign {s78[59],s77[58]} = {1'b0,s63[58]} + {1'b0,s62[58]} + {1'b0,s61[58]};
assign {s78[60],s77[59]} = {1'b0,s63[59]} + {1'b0,s62[59]} + {1'b0,s61[59]};
assign {s78[61],s77[60]} = {1'b0,s63[60]} + {1'b0,s62[60]} + {1'b0,s61[60]};
assign {s78[62],s77[61]} = {1'b0,s63[61]} + {1'b0,s62[61]} + {1'b0,s61[61]};
assign {s78[63],s77[62]} = {1'b0,s63[62]} + {1'b0,s62[62]} + {1'b0,s61[62]};
assign {s78[64],s77[63]} = {1'b0,s63[63]} + {1'b0,s62[63]} + {1'b0,s61[63]};
assign {s78[65],s77[64]} = {1'b0,s63[64]} + {1'b0,s62[64]} + {1'b0,s61[64]};
assign {s78[66],s77[65]} = {1'b0,s63[65]} + {1'b0,s62[65]} + {1'b0,s61[65]};
assign {s78[67],s77[66]} = {1'b0,s63[66]} + {1'b0,s62[66]} + {1'b0,s61[66]};
assign {s80[6],s79[5]} = {1'b0,s64[5]};
assign {s80[7],s79[6]} = {1'b0,s64[6]};
assign {s80[8],s79[7]} = {1'b0,s64[7]};
assign {s80[9],s79[8]} = {1'b0,s64[8]};
assign {s80[10],s79[9]} = {1'b0,s65[9]} + {1'b0,s64[9]};
assign {s80[11],s79[10]} = {1'b0,s66[10]} + {1'b0,s65[10]} + {1'b0,s64[10]};
assign {s80[12],s79[11]} = {1'b0,s66[11]} + {1'b0,s65[11]} + {1'b0,s64[11]};
assign {s80[13],s79[12]} = {1'b0,s66[12]} + {1'b0,s65[12]} + {1'b0,s64[12]};
assign {s80[14],s79[13]} = {1'b0,s66[13]} + {1'b0,s65[13]} + {1'b0,s64[13]};
assign {s80[15],s79[14]} = {1'b0,s66[14]} + {1'b0,s65[14]} + {1'b0,s64[14]};
assign {s80[16],s79[15]} = {1'b0,s66[15]} + {1'b0,s65[15]} + {1'b0,s64[15]};
assign {s80[17],s79[16]} = {1'b0,s66[16]} + {1'b0,s65[16]} + {1'b0,s64[16]};
assign {s80[18],s79[17]} = {1'b0,s66[17]} + {1'b0,s65[17]} + {1'b0,s64[17]};
assign {s80[19],s79[18]} = {1'b0,s66[18]} + {1'b0,s65[18]} + {1'b0,s64[18]};
assign {s80[20],s79[19]} = {1'b0,s66[19]} + {1'b0,s65[19]} + {1'b0,s64[19]};
assign {s80[21],s79[20]} = {1'b0,s66[20]} + {1'b0,s65[20]} + {1'b0,s64[20]};
assign {s80[22],s79[21]} = {1'b0,s66[21]} + {1'b0,s65[21]} + {1'b0,s64[21]};
assign {s80[23],s79[22]} = {1'b0,s66[22]} + {1'b0,s65[22]} + {1'b0,s64[22]};
assign {s80[24],s79[23]} = {1'b0,s66[23]} + {1'b0,s65[23]} + {1'b0,s64[23]};
assign {s80[25],s79[24]} = {1'b0,s66[24]} + {1'b0,s65[24]} + {1'b0,s64[24]};
assign {s80[26],s79[25]} = {1'b0,s66[25]} + {1'b0,s65[25]} + {1'b0,s64[25]};
assign {s80[27],s79[26]} = {1'b0,s66[26]} + {1'b0,s65[26]} + {1'b0,s64[26]};
assign {s80[28],s79[27]} = {1'b0,s66[27]} + {1'b0,s65[27]} + {1'b0,s64[27]};
assign {s80[29],s79[28]} = {1'b0,s66[28]} + {1'b0,s65[28]} + {1'b0,s64[28]};
assign {s80[30],s79[29]} = {1'b0,s66[29]} + {1'b0,s65[29]} + {1'b0,s64[29]};
assign {s80[31],s79[30]} = {1'b0,s66[30]} + {1'b0,s65[30]} + {1'b0,s64[30]};
assign {s80[32],s79[31]} = {1'b0,s66[31]} + {1'b0,s65[31]} + {1'b0,s64[31]};
assign {s80[33],s79[32]} = {1'b0,s66[32]} + {1'b0,s65[32]} + {1'b0,s64[32]};
assign {s80[34],s79[33]} = {1'b0,s66[33]} + {1'b0,s65[33]} + {1'b0,s64[33]};
assign {s80[35],s79[34]} = {1'b0,s66[34]} + {1'b0,s65[34]} + {1'b0,s64[34]};
assign {s80[36],s79[35]} = {1'b0,s66[35]} + {1'b0,s65[35]} + {1'b0,s64[35]};
assign {s80[37],s79[36]} = {1'b0,s66[36]} + {1'b0,s65[36]} + {1'b0,s64[36]};
assign {s80[38],s79[37]} = {1'b0,s66[37]} + {1'b0,s65[37]} + {1'b0,s64[37]};
assign {s80[39],s79[38]} = {1'b0,s66[38]} + {1'b0,s65[38]} + {1'b0,s64[38]};
assign {s80[40],s79[39]} = {1'b0,s66[39]} + {1'b0,s65[39]} + {1'b0,s64[39]};
assign {s80[41],s79[40]} = {1'b0,s66[40]} + {1'b0,s65[40]} + {1'b0,s64[40]};
assign {s80[42],s79[41]} = {1'b0,s66[41]} + {1'b0,s65[41]} + {1'b0,s64[41]};
assign {s80[43],s79[42]} = {1'b0,s66[42]} + {1'b0,s65[42]} + {1'b0,s64[42]};
assign {s80[44],s79[43]} = {1'b0,s66[43]} + {1'b0,s65[43]} + {1'b0,s64[43]};
assign {s80[45],s79[44]} = {1'b0,s66[44]} + {1'b0,s65[44]} + {1'b0,s64[44]};
assign {s80[46],s79[45]} = {1'b0,s66[45]} + {1'b0,s65[45]} + {1'b0,s64[45]};
assign {s80[47],s79[46]} = {1'b0,s66[46]} + {1'b0,s65[46]} + {1'b0,s64[46]};
assign {s80[48],s79[47]} = {1'b0,s66[47]} + {1'b0,s65[47]} + {1'b0,s64[47]};
assign {s80[49],s79[48]} = {1'b0,s66[48]} + {1'b0,s65[48]} + {1'b0,s64[48]};
assign {s80[50],s79[49]} = {1'b0,s66[49]} + {1'b0,s65[49]} + {1'b0,s64[49]};
assign {s80[51],s79[50]} = {1'b0,s66[50]} + {1'b0,s65[50]} + {1'b0,s64[50]};
assign {s80[52],s79[51]} = {1'b0,s66[51]} + {1'b0,s65[51]} + {1'b0,s64[51]};
assign {s80[53],s79[52]} = {1'b0,s66[52]} + {1'b0,s65[52]} + {1'b0,s64[52]};
assign {s80[54],s79[53]} = {1'b0,s66[53]} + {1'b0,s65[53]} + {1'b0,s64[53]};
assign {s80[55],s79[54]} = {1'b0,s66[54]} + {1'b0,s65[54]} + {1'b0,s64[54]};
assign {s80[56],s79[55]} = {1'b0,s66[55]} + {1'b0,s65[55]} + {1'b0,s64[55]};
assign {s80[57],s79[56]} = {1'b0,s66[56]} + {1'b0,s65[56]} + {1'b0,s64[56]};
assign {s80[58],s79[57]} = {1'b0,s66[57]} + {1'b0,s65[57]} + {1'b0,s64[57]};
assign {s80[59],s79[58]} = {1'b0,s66[58]} + {1'b0,s65[58]} + {1'b0,s64[58]};
assign {s80[60],s79[59]} = {1'b0,s66[59]} + {1'b0,s65[59]} + {1'b0,s64[59]};
assign {s80[61],s79[60]} = {1'b0,s66[60]} + {1'b0,s65[60]} + {1'b0,s64[60]};
assign {s80[62],s79[61]} = {1'b0,s66[61]} + {1'b0,s65[61]} + {1'b0,s64[61]};
assign {s80[63],s79[62]} = {1'b0,s66[62]} + {1'b0,s65[62]} + {1'b0,s64[62]};
assign {s80[64],s79[63]} = {1'b0,s66[63]} + {1'b0,s65[63]} + {1'b0,s64[63]};
assign {s80[65],s79[64]} = {1'b0,s66[64]} + {1'b0,s65[64]} + {1'b0,s64[64]};
assign {s80[66],s79[65]} = {1'b0,s66[65]} + {1'b0,s65[65]} + {1'b0,s64[65]};
assign {s80[67],s79[66]} = {1'b0,s66[66]} + {1'b0,s65[66]} + {1'b0,s64[66]};
assign {s82[14],s81[13]} = {1'b0,s67[13]};
assign {s82[15],s81[14]} = {1'b0,s68[14]} + {1'b0,s67[14]};
assign {s82[16],s81[15]} = {1'b0,s68[15]} + {1'b0,s67[15]};
assign {s82[17],s81[16]} = {1'b0,s68[16]} + {1'b0,s67[16]};
assign {s82[18],s81[17]} = {1'b0,s68[17]} + {1'b0,s67[17]};
assign {s82[19],s81[18]} = {1'b0,s69[18]} + {1'b0,s68[18]} + {1'b0,s67[18]};
assign {s82[20],s81[19]} = {1'b0,s69[19]} + {1'b0,s68[19]} + {1'b0,s67[19]};
assign {s82[21],s81[20]} = {1'b0,s69[20]} + {1'b0,s68[20]} + {1'b0,s67[20]};
assign {s82[22],s81[21]} = {1'b0,s69[21]} + {1'b0,s68[21]} + {1'b0,s67[21]};
assign {s82[23],s81[22]} = {1'b0,s69[22]} + {1'b0,s68[22]} + {1'b0,s67[22]};
assign {s82[24],s81[23]} = {1'b0,s69[23]} + {1'b0,s68[23]} + {1'b0,s67[23]};
assign {s82[25],s81[24]} = {1'b0,s69[24]} + {1'b0,s68[24]} + {1'b0,s67[24]};
assign {s82[26],s81[25]} = {1'b0,s69[25]} + {1'b0,s68[25]} + {1'b0,s67[25]};
assign {s82[27],s81[26]} = {1'b0,s69[26]} + {1'b0,s68[26]} + {1'b0,s67[26]};
assign {s82[28],s81[27]} = {1'b0,s69[27]} + {1'b0,s68[27]} + {1'b0,s67[27]};
assign {s82[29],s81[28]} = {1'b0,s69[28]} + {1'b0,s68[28]} + {1'b0,s67[28]};
assign {s82[30],s81[29]} = {1'b0,s69[29]} + {1'b0,s68[29]} + {1'b0,s67[29]};
assign {s82[31],s81[30]} = {1'b0,s69[30]} + {1'b0,s68[30]} + {1'b0,s67[30]};
assign {s82[32],s81[31]} = {1'b0,s69[31]} + {1'b0,s68[31]} + {1'b0,s67[31]};
assign {s82[33],s81[32]} = {1'b0,s69[32]} + {1'b0,s68[32]} + {1'b0,s67[32]};
assign {s82[34],s81[33]} = {1'b0,s69[33]} + {1'b0,s68[33]} + {1'b0,s67[33]};
assign {s82[35],s81[34]} = {1'b0,s69[34]} + {1'b0,s68[34]} + {1'b0,s67[34]};
assign {s82[36],s81[35]} = {1'b0,s69[35]} + {1'b0,s68[35]} + {1'b0,s67[35]};
assign {s82[37],s81[36]} = {1'b0,s69[36]} + {1'b0,s68[36]} + {1'b0,s67[36]};
assign {s82[38],s81[37]} = {1'b0,s69[37]} + {1'b0,s68[37]} + {1'b0,s67[37]};
assign {s82[39],s81[38]} = {1'b0,s69[38]} + {1'b0,s68[38]} + {1'b0,s67[38]};
assign {s82[40],s81[39]} = {1'b0,s69[39]} + {1'b0,s68[39]} + {1'b0,s67[39]};
assign {s82[41],s81[40]} = {1'b0,s69[40]} + {1'b0,s68[40]} + {1'b0,s67[40]};
assign {s82[42],s81[41]} = {1'b0,s69[41]} + {1'b0,s68[41]} + {1'b0,s67[41]};
assign {s82[43],s81[42]} = {1'b0,s69[42]} + {1'b0,s68[42]} + {1'b0,s67[42]};
assign {s82[44],s81[43]} = {1'b0,s69[43]} + {1'b0,s68[43]} + {1'b0,s67[43]};
assign {s82[45],s81[44]} = {1'b0,s69[44]} + {1'b0,s68[44]} + {1'b0,s67[44]};
assign {s82[46],s81[45]} = {1'b0,s69[45]} + {1'b0,s68[45]} + {1'b0,s67[45]};
assign {s82[47],s81[46]} = {1'b0,s69[46]} + {1'b0,s68[46]} + {1'b0,s67[46]};
assign {s82[48],s81[47]} = {1'b0,s69[47]} + {1'b0,s68[47]} + {1'b0,s67[47]};
assign {s82[49],s81[48]} = {1'b0,s69[48]} + {1'b0,s68[48]} + {1'b0,s67[48]};
assign {s82[50],s81[49]} = {1'b0,s69[49]} + {1'b0,s68[49]} + {1'b0,s67[49]};
assign {s82[51],s81[50]} = {1'b0,s69[50]} + {1'b0,s68[50]} + {1'b0,s67[50]};
assign {s82[52],s81[51]} = {1'b0,s69[51]} + {1'b0,s68[51]} + {1'b0,s67[51]};
assign {s82[53],s81[52]} = {1'b0,s69[52]} + {1'b0,s68[52]} + {1'b0,s67[52]};
assign {s82[54],s81[53]} = {1'b0,s69[53]} + {1'b0,s68[53]} + {1'b0,s67[53]};
assign {s82[55],s81[54]} = {1'b0,s69[54]} + {1'b0,s68[54]} + {1'b0,s67[54]};
assign {s82[56],s81[55]} = {1'b0,s69[55]} + {1'b0,s68[55]} + {1'b0,s67[55]};
assign {s82[57],s81[56]} = {1'b0,s69[56]} + {1'b0,s68[56]} + {1'b0,s67[56]};
assign {s82[58],s81[57]} = {1'b0,s69[57]} + {1'b0,s68[57]} + {1'b0,s67[57]};
assign {s82[59],s81[58]} = {1'b0,s69[58]} + {1'b0,s68[58]} + {1'b0,s67[58]};
assign {s82[60],s81[59]} = {1'b0,s69[59]} + {1'b0,s68[59]} + {1'b0,s67[59]};
assign {s82[61],s81[60]} = {1'b0,s69[60]} + {1'b0,s68[60]} + {1'b0,s67[60]};
assign {s82[62],s81[61]} = {1'b0,s69[61]} + {1'b0,s68[61]} + {1'b0,s67[61]};
assign {s82[63],s81[62]} = {1'b0,s69[62]} + {1'b0,s68[62]} + {1'b0,s67[62]};
assign {s82[64],s81[63]} = {1'b0,s69[63]} + {1'b0,s68[63]} + {1'b0,s67[63]};
assign {s82[65],s81[64]} = {1'b0,s69[64]} + {1'b0,s68[64]} + {1'b0,s67[64]};
assign {s82[66],s81[65]} = {1'b0,s69[65]} + {1'b0,s68[65]} + {1'b0,s67[65]};
assign {s82[67],s81[66]} = {1'b0,s69[66]} + {1'b0,s68[66]} + {1'b0,s67[66]};
assign {s84[20],s83[19]} = {1'b0,s70[19]};
assign {s84[21],s83[20]} = {1'b0,s70[20]};
assign {s84[22],s83[21]} = {1'b0,s70[21]};
assign {s84[23],s83[22]} = {1'b0,s71[22]} + {1'b0,s70[22]};
assign {s84[24],s83[23]} = {1'b0,s72[23]} + {1'b0,s71[23]} + {1'b0,s70[23]};
assign {s84[25],s83[24]} = {1'b0,s72[24]} + {1'b0,s71[24]} + {1'b0,s70[24]};
assign {s84[26],s83[25]} = {1'b0,s72[25]} + {1'b0,s71[25]} + {1'b0,s70[25]};
assign {s84[27],s83[26]} = {1'b0,s72[26]} + {1'b0,s71[26]} + {1'b0,s70[26]};
assign {s84[28],s83[27]} = {1'b0,s72[27]} + {1'b0,s71[27]} + {1'b0,s70[27]};
assign {s84[29],s83[28]} = {1'b0,s72[28]} + {1'b0,s71[28]} + {1'b0,s70[28]};
assign {s84[30],s83[29]} = {1'b0,s72[29]} + {1'b0,s71[29]} + {1'b0,s70[29]};
assign {s84[31],s83[30]} = {1'b0,s72[30]} + {1'b0,s71[30]} + {1'b0,s70[30]};
assign {s84[32],s83[31]} = {1'b0,s72[31]} + {1'b0,s71[31]} + {1'b0,s70[31]};
assign {s84[33],s83[32]} = {1'b0,s72[32]} + {1'b0,s71[32]} + {1'b0,s70[32]};
assign {s84[34],s83[33]} = {1'b0,s72[33]} + {1'b0,s71[33]} + {1'b0,s70[33]};
assign {s84[35],s83[34]} = {1'b0,s72[34]} + {1'b0,s71[34]} + {1'b0,s70[34]};
assign {s84[36],s83[35]} = {1'b0,s72[35]} + {1'b0,s71[35]} + {1'b0,s70[35]};
assign {s84[37],s83[36]} = {1'b0,s72[36]} + {1'b0,s71[36]} + {1'b0,s70[36]};
assign {s84[38],s83[37]} = {1'b0,s72[37]} + {1'b0,s71[37]} + {1'b0,s70[37]};
assign {s84[39],s83[38]} = {1'b0,s72[38]} + {1'b0,s71[38]} + {1'b0,s70[38]};
assign {s84[40],s83[39]} = {1'b0,s72[39]} + {1'b0,s71[39]} + {1'b0,s70[39]};
assign {s84[41],s83[40]} = {1'b0,s72[40]} + {1'b0,s71[40]} + {1'b0,s70[40]};
assign {s84[42],s83[41]} = {1'b0,s72[41]} + {1'b0,s71[41]} + {1'b0,s70[41]};
assign {s84[43],s83[42]} = {1'b0,s72[42]} + {1'b0,s71[42]} + {1'b0,s70[42]};
assign {s84[44],s83[43]} = {1'b0,s72[43]} + {1'b0,s71[43]} + {1'b0,s70[43]};
assign {s84[45],s83[44]} = {1'b0,s72[44]} + {1'b0,s71[44]} + {1'b0,s70[44]};
assign {s84[46],s83[45]} = {1'b0,s72[45]} + {1'b0,s71[45]} + {1'b0,s70[45]};
assign {s84[47],s83[46]} = {1'b0,s72[46]} + {1'b0,s71[46]} + {1'b0,s70[46]};
assign {s84[48],s83[47]} = {1'b0,s72[47]} + {1'b0,s71[47]} + {1'b0,s70[47]};
assign {s84[49],s83[48]} = {1'b0,s72[48]} + {1'b0,s71[48]} + {1'b0,s70[48]};
assign {s84[50],s83[49]} = {1'b0,s72[49]} + {1'b0,s71[49]} + {1'b0,s70[49]};
assign {s84[51],s83[50]} = {1'b0,s72[50]} + {1'b0,s71[50]} + {1'b0,s70[50]};
assign {s84[52],s83[51]} = {1'b0,s72[51]} + {1'b0,s71[51]} + {1'b0,s70[51]};
assign {s84[53],s83[52]} = {1'b0,s72[52]} + {1'b0,s71[52]} + {1'b0,s70[52]};
assign {s84[54],s83[53]} = {1'b0,s72[53]} + {1'b0,s71[53]} + {1'b0,s70[53]};
assign {s84[55],s83[54]} = {1'b0,s72[54]} + {1'b0,s71[54]} + {1'b0,s70[54]};
assign {s84[56],s83[55]} = {1'b0,s72[55]} + {1'b0,s71[55]} + {1'b0,s70[55]};
assign {s84[57],s83[56]} = {1'b0,s72[56]} + {1'b0,s71[56]} + {1'b0,s70[56]};
assign {s84[58],s83[57]} = {1'b0,s72[57]} + {1'b0,s71[57]} + {1'b0,s70[57]};
assign {s84[59],s83[58]} = {1'b0,s72[58]} + {1'b0,s71[58]} + {1'b0,s70[58]};
assign {s84[60],s83[59]} = {1'b0,s72[59]} + {1'b0,s71[59]} + {1'b0,s70[59]};
assign {s84[61],s83[60]} = {1'b0,s72[60]} + {1'b0,s71[60]} + {1'b0,s70[60]};
assign {s84[62],s83[61]} = {1'b0,s72[61]} + {1'b0,s71[61]} + {1'b0,s70[61]};
assign {s84[63],s83[62]} = {1'b0,s72[62]} + {1'b0,s71[62]} + {1'b0,s70[62]};
assign {s84[64],s83[63]} = {1'b0,s72[63]} + {1'b0,s71[63]} + {1'b0,s70[63]};
assign {s84[65],s83[64]} = {1'b0,s72[64]} + {1'b0,s71[64]} + {1'b0,s70[64]};
assign {s84[66],s83[65]} = {1'b0,s72[65]} + {1'b0,s71[65]} + {1'b0,s70[65]};
assign {s84[67],s83[66]} = {1'b0,s72[66]} + {1'b0,s71[66]} + {1'b0,s70[66]};
assign {s86[28],s85[27]} = {1'b0,s73[27]};
assign {s86[29],s85[28]} = {1'b0,s74[28]} + {1'b0,s73[28]};
assign {s86[30],s85[29]} = {1'b0,s74[29]} + {1'b0,s73[29]};
assign {s86[31],s85[30]} = {1'b0,s74[30]} + {1'b0,s73[30]};
assign {s86[32],s85[31]} = {1'b0,s75[31]} + {1'b0,s74[31]} + {1'b0,s73[31]};
assign {s86[33],s85[32]} = {1'b0,s75[32]} + {1'b0,s74[32]} + {1'b0,s73[32]};
assign {s86[34],s85[33]} = {1'b0,s75[33]} + {1'b0,s74[33]} + {1'b0,s73[33]};
assign {s86[35],s85[34]} = {1'b0,s75[34]} + {1'b0,s74[34]} + {1'b0,s73[34]};
assign {s86[36],s85[35]} = {1'b0,s75[35]} + {1'b0,s74[35]} + {1'b0,s73[35]};
assign {s86[37],s85[36]} = {1'b0,s75[36]} + {1'b0,s74[36]} + {1'b0,s73[36]};
assign {s86[38],s85[37]} = {1'b0,s75[37]} + {1'b0,s74[37]} + {1'b0,s73[37]};
assign {s86[39],s85[38]} = {1'b0,s75[38]} + {1'b0,s74[38]} + {1'b0,s73[38]};
assign {s86[40],s85[39]} = {1'b0,s75[39]} + {1'b0,s74[39]} + {1'b0,s73[39]};
assign {s86[41],s85[40]} = {1'b0,s75[40]} + {1'b0,s74[40]} + {1'b0,s73[40]};
assign {s86[42],s85[41]} = {1'b0,s75[41]} + {1'b0,s74[41]} + {1'b0,s73[41]};
assign {s86[43],s85[42]} = {1'b0,s75[42]} + {1'b0,s74[42]} + {1'b0,s73[42]};
assign {s86[44],s85[43]} = {1'b0,s75[43]} + {1'b0,s74[43]} + {1'b0,s73[43]};
assign {s86[45],s85[44]} = {1'b0,s75[44]} + {1'b0,s74[44]} + {1'b0,s73[44]};
assign {s86[46],s85[45]} = {1'b0,s75[45]} + {1'b0,s74[45]} + {1'b0,s73[45]};
assign {s86[47],s85[46]} = {1'b0,s75[46]} + {1'b0,s74[46]} + {1'b0,s73[46]};
assign {s86[48],s85[47]} = {1'b0,s75[47]} + {1'b0,s74[47]} + {1'b0,s73[47]};
assign {s86[49],s85[48]} = {1'b0,s75[48]} + {1'b0,s74[48]} + {1'b0,s73[48]};
assign {s86[50],s85[49]} = {1'b0,s75[49]} + {1'b0,s74[49]} + {1'b0,s73[49]};
assign {s86[51],s85[50]} = {1'b0,s75[50]} + {1'b0,s74[50]} + {1'b0,s73[50]};
assign {s86[52],s85[51]} = {1'b0,s75[51]} + {1'b0,s74[51]} + {1'b0,s73[51]};
assign {s86[53],s85[52]} = {1'b0,s75[52]} + {1'b0,s74[52]} + {1'b0,s73[52]};
assign {s86[54],s85[53]} = {1'b0,s75[53]} + {1'b0,s74[53]} + {1'b0,s73[53]};
assign {s86[55],s85[54]} = {1'b0,s75[54]} + {1'b0,s74[54]} + {1'b0,s73[54]};
assign {s86[56],s85[55]} = {1'b0,s75[55]} + {1'b0,s74[55]} + {1'b0,s73[55]};
assign {s86[57],s85[56]} = {1'b0,s75[56]} + {1'b0,s74[56]} + {1'b0,s73[56]};
assign {s86[58],s85[57]} = {1'b0,s75[57]} + {1'b0,s74[57]} + {1'b0,s73[57]};
assign {s86[59],s85[58]} = {1'b0,s75[58]} + {1'b0,s74[58]} + {1'b0,s73[58]};
assign {s86[60],s85[59]} = {1'b0,s75[59]} + {1'b0,s74[59]} + {1'b0,s73[59]};
assign {s86[61],s85[60]} = {1'b0,s75[60]} + {1'b0,s74[60]} + {1'b0,s73[60]};
assign {s86[62],s85[61]} = {1'b0,s75[61]} + {1'b0,s74[61]} + {1'b0,s73[61]};
assign {s86[63],s85[62]} = {1'b0,s75[62]} + {1'b0,s74[62]} + {1'b0,s73[62]};
assign {s86[64],s85[63]} = {1'b0,s75[63]} + {1'b0,s74[63]} + {1'b0,s73[63]};
assign {s86[65],s85[64]} = {1'b0,s75[64]} + {1'b0,s74[64]} + {1'b0,s73[64]};
assign {s86[66],s85[65]} = {1'b0,s75[65]} + {1'b0,s74[65]} + {1'b0,s73[65]};
assign {s86[67],s85[66]} = {1'b0,s75[66]} + {1'b0,s74[66]} + {1'b0,s73[66]};
assign s87 = s76[(PPLEN - 1):32];
assign {s89[1],s88[0]} = {1'b0,s77[0]};
assign {s89[2],s88[1]} = {1'b0,s78[1]} + {1'b0,s77[1]};
assign {s89[3],s88[2]} = {1'b0,s78[2]} + {1'b0,s77[2]};
assign {s89[4],s88[3]} = {1'b0,s78[3]} + {1'b0,s77[3]};
assign {s89[5],s88[4]} = {1'b0,s78[4]} + {1'b0,s77[4]};
assign {s89[6],s88[5]} = {1'b0,s79[5]} + {1'b0,s78[5]} + {1'b0,s77[5]};
assign {s89[7],s88[6]} = {1'b0,s79[6]} + {1'b0,s78[6]} + {1'b0,s77[6]};
assign {s89[8],s88[7]} = {1'b0,s79[7]} + {1'b0,s78[7]} + {1'b0,s77[7]};
assign {s89[9],s88[8]} = {1'b0,s79[8]} + {1'b0,s78[8]} + {1'b0,s77[8]};
assign {s89[10],s88[9]} = {1'b0,s79[9]} + {1'b0,s78[9]} + {1'b0,s77[9]};
assign {s89[11],s88[10]} = {1'b0,s79[10]} + {1'b0,s78[10]} + {1'b0,s77[10]};
assign {s89[12],s88[11]} = {1'b0,s79[11]} + {1'b0,s78[11]} + {1'b0,s77[11]};
assign {s89[13],s88[12]} = {1'b0,s79[12]} + {1'b0,s78[12]} + {1'b0,s77[12]};
assign {s89[14],s88[13]} = {1'b0,s79[13]} + {1'b0,s78[13]} + {1'b0,s77[13]};
assign {s89[15],s88[14]} = {1'b0,s79[14]} + {1'b0,s78[14]} + {1'b0,s77[14]};
assign {s89[16],s88[15]} = {1'b0,s79[15]} + {1'b0,s78[15]} + {1'b0,s77[15]};
assign {s89[17],s88[16]} = {1'b0,s79[16]} + {1'b0,s78[16]} + {1'b0,s77[16]};
assign {s89[18],s88[17]} = {1'b0,s79[17]} + {1'b0,s78[17]} + {1'b0,s77[17]};
assign {s89[19],s88[18]} = {1'b0,s79[18]} + {1'b0,s78[18]} + {1'b0,s77[18]};
assign {s89[20],s88[19]} = {1'b0,s79[19]} + {1'b0,s78[19]} + {1'b0,s77[19]};
assign {s89[21],s88[20]} = {1'b0,s79[20]} + {1'b0,s78[20]} + {1'b0,s77[20]};
assign {s89[22],s88[21]} = {1'b0,s79[21]} + {1'b0,s78[21]} + {1'b0,s77[21]};
assign {s89[23],s88[22]} = {1'b0,s79[22]} + {1'b0,s78[22]} + {1'b0,s77[22]};
assign {s89[24],s88[23]} = {1'b0,s79[23]} + {1'b0,s78[23]} + {1'b0,s77[23]};
assign {s89[25],s88[24]} = {1'b0,s79[24]} + {1'b0,s78[24]} + {1'b0,s77[24]};
assign {s89[26],s88[25]} = {1'b0,s79[25]} + {1'b0,s78[25]} + {1'b0,s77[25]};
assign {s89[27],s88[26]} = {1'b0,s79[26]} + {1'b0,s78[26]} + {1'b0,s77[26]};
assign {s89[28],s88[27]} = {1'b0,s79[27]} + {1'b0,s78[27]} + {1'b0,s77[27]};
assign {s89[29],s88[28]} = {1'b0,s79[28]} + {1'b0,s78[28]} + {1'b0,s77[28]};
assign {s89[30],s88[29]} = {1'b0,s79[29]} + {1'b0,s78[29]} + {1'b0,s77[29]};
assign {s89[31],s88[30]} = {1'b0,s79[30]} + {1'b0,s78[30]} + {1'b0,s77[30]};
assign {s89[32],s88[31]} = {1'b0,s79[31]} + {1'b0,s78[31]} + {1'b0,s77[31]};
assign {s89[33],s88[32]} = {1'b0,s79[32]} + {1'b0,s78[32]} + {1'b0,s77[32]};
assign {s89[34],s88[33]} = {1'b0,s79[33]} + {1'b0,s78[33]} + {1'b0,s77[33]};
assign {s89[35],s88[34]} = {1'b0,s79[34]} + {1'b0,s78[34]} + {1'b0,s77[34]};
assign {s89[36],s88[35]} = {1'b0,s79[35]} + {1'b0,s78[35]} + {1'b0,s77[35]};
assign {s89[37],s88[36]} = {1'b0,s79[36]} + {1'b0,s78[36]} + {1'b0,s77[36]};
assign {s89[38],s88[37]} = {1'b0,s79[37]} + {1'b0,s78[37]} + {1'b0,s77[37]};
assign {s89[39],s88[38]} = {1'b0,s79[38]} + {1'b0,s78[38]} + {1'b0,s77[38]};
assign {s89[40],s88[39]} = {1'b0,s79[39]} + {1'b0,s78[39]} + {1'b0,s77[39]};
assign {s89[41],s88[40]} = {1'b0,s79[40]} + {1'b0,s78[40]} + {1'b0,s77[40]};
assign {s89[42],s88[41]} = {1'b0,s79[41]} + {1'b0,s78[41]} + {1'b0,s77[41]};
assign {s89[43],s88[42]} = {1'b0,s79[42]} + {1'b0,s78[42]} + {1'b0,s77[42]};
assign {s89[44],s88[43]} = {1'b0,s79[43]} + {1'b0,s78[43]} + {1'b0,s77[43]};
assign {s89[45],s88[44]} = {1'b0,s79[44]} + {1'b0,s78[44]} + {1'b0,s77[44]};
assign {s89[46],s88[45]} = {1'b0,s79[45]} + {1'b0,s78[45]} + {1'b0,s77[45]};
assign {s89[47],s88[46]} = {1'b0,s79[46]} + {1'b0,s78[46]} + {1'b0,s77[46]};
assign {s89[48],s88[47]} = {1'b0,s79[47]} + {1'b0,s78[47]} + {1'b0,s77[47]};
assign {s89[49],s88[48]} = {1'b0,s79[48]} + {1'b0,s78[48]} + {1'b0,s77[48]};
assign {s89[50],s88[49]} = {1'b0,s79[49]} + {1'b0,s78[49]} + {1'b0,s77[49]};
assign {s89[51],s88[50]} = {1'b0,s79[50]} + {1'b0,s78[50]} + {1'b0,s77[50]};
assign {s89[52],s88[51]} = {1'b0,s79[51]} + {1'b0,s78[51]} + {1'b0,s77[51]};
assign {s89[53],s88[52]} = {1'b0,s79[52]} + {1'b0,s78[52]} + {1'b0,s77[52]};
assign {s89[54],s88[53]} = {1'b0,s79[53]} + {1'b0,s78[53]} + {1'b0,s77[53]};
assign {s89[55],s88[54]} = {1'b0,s79[54]} + {1'b0,s78[54]} + {1'b0,s77[54]};
assign {s89[56],s88[55]} = {1'b0,s79[55]} + {1'b0,s78[55]} + {1'b0,s77[55]};
assign {s89[57],s88[56]} = {1'b0,s79[56]} + {1'b0,s78[56]} + {1'b0,s77[56]};
assign {s89[58],s88[57]} = {1'b0,s79[57]} + {1'b0,s78[57]} + {1'b0,s77[57]};
assign {s89[59],s88[58]} = {1'b0,s79[58]} + {1'b0,s78[58]} + {1'b0,s77[58]};
assign {s89[60],s88[59]} = {1'b0,s79[59]} + {1'b0,s78[59]} + {1'b0,s77[59]};
assign {s89[61],s88[60]} = {1'b0,s79[60]} + {1'b0,s78[60]} + {1'b0,s77[60]};
assign {s89[62],s88[61]} = {1'b0,s79[61]} + {1'b0,s78[61]} + {1'b0,s77[61]};
assign {s89[63],s88[62]} = {1'b0,s79[62]} + {1'b0,s78[62]} + {1'b0,s77[62]};
assign {s89[64],s88[63]} = {1'b0,s79[63]} + {1'b0,s78[63]} + {1'b0,s77[63]};
assign {s89[65],s88[64]} = {1'b0,s79[64]} + {1'b0,s78[64]} + {1'b0,s77[64]};
assign {s89[66],s88[65]} = {1'b0,s79[65]} + {1'b0,s78[65]} + {1'b0,s77[65]};
assign {s89[67],s88[66]} = {1'b0,s79[66]} + {1'b0,s78[66]} + {1'b0,s77[66]};
assign {s91[7],s90[6]} = {1'b0,s80[6]};
assign {s91[8],s90[7]} = {1'b0,s80[7]};
assign {s91[9],s90[8]} = {1'b0,s80[8]};
assign {s91[10],s90[9]} = {1'b0,s80[9]};
assign {s91[11],s90[10]} = {1'b0,s80[10]};
assign {s91[12],s90[11]} = {1'b0,s80[11]};
assign {s91[13],s90[12]} = {1'b0,s80[12]};
assign {s91[14],s90[13]} = {1'b0,s81[13]} + {1'b0,s80[13]};
assign {s91[15],s90[14]} = {1'b0,s82[14]} + {1'b0,s81[14]} + {1'b0,s80[14]};
assign {s91[16],s90[15]} = {1'b0,s82[15]} + {1'b0,s81[15]} + {1'b0,s80[15]};
assign {s91[17],s90[16]} = {1'b0,s82[16]} + {1'b0,s81[16]} + {1'b0,s80[16]};
assign {s91[18],s90[17]} = {1'b0,s82[17]} + {1'b0,s81[17]} + {1'b0,s80[17]};
assign {s91[19],s90[18]} = {1'b0,s82[18]} + {1'b0,s81[18]} + {1'b0,s80[18]};
assign {s91[20],s90[19]} = {1'b0,s82[19]} + {1'b0,s81[19]} + {1'b0,s80[19]};
assign {s91[21],s90[20]} = {1'b0,s82[20]} + {1'b0,s81[20]} + {1'b0,s80[20]};
assign {s91[22],s90[21]} = {1'b0,s82[21]} + {1'b0,s81[21]} + {1'b0,s80[21]};
assign {s91[23],s90[22]} = {1'b0,s82[22]} + {1'b0,s81[22]} + {1'b0,s80[22]};
assign {s91[24],s90[23]} = {1'b0,s82[23]} + {1'b0,s81[23]} + {1'b0,s80[23]};
assign {s91[25],s90[24]} = {1'b0,s82[24]} + {1'b0,s81[24]} + {1'b0,s80[24]};
assign {s91[26],s90[25]} = {1'b0,s82[25]} + {1'b0,s81[25]} + {1'b0,s80[25]};
assign {s91[27],s90[26]} = {1'b0,s82[26]} + {1'b0,s81[26]} + {1'b0,s80[26]};
assign {s91[28],s90[27]} = {1'b0,s82[27]} + {1'b0,s81[27]} + {1'b0,s80[27]};
assign {s91[29],s90[28]} = {1'b0,s82[28]} + {1'b0,s81[28]} + {1'b0,s80[28]};
assign {s91[30],s90[29]} = {1'b0,s82[29]} + {1'b0,s81[29]} + {1'b0,s80[29]};
assign {s91[31],s90[30]} = {1'b0,s82[30]} + {1'b0,s81[30]} + {1'b0,s80[30]};
assign {s91[32],s90[31]} = {1'b0,s82[31]} + {1'b0,s81[31]} + {1'b0,s80[31]};
assign {s91[33],s90[32]} = {1'b0,s82[32]} + {1'b0,s81[32]} + {1'b0,s80[32]};
assign {s91[34],s90[33]} = {1'b0,s82[33]} + {1'b0,s81[33]} + {1'b0,s80[33]};
assign {s91[35],s90[34]} = {1'b0,s82[34]} + {1'b0,s81[34]} + {1'b0,s80[34]};
assign {s91[36],s90[35]} = {1'b0,s82[35]} + {1'b0,s81[35]} + {1'b0,s80[35]};
assign {s91[37],s90[36]} = {1'b0,s82[36]} + {1'b0,s81[36]} + {1'b0,s80[36]};
assign {s91[38],s90[37]} = {1'b0,s82[37]} + {1'b0,s81[37]} + {1'b0,s80[37]};
assign {s91[39],s90[38]} = {1'b0,s82[38]} + {1'b0,s81[38]} + {1'b0,s80[38]};
assign {s91[40],s90[39]} = {1'b0,s82[39]} + {1'b0,s81[39]} + {1'b0,s80[39]};
assign {s91[41],s90[40]} = {1'b0,s82[40]} + {1'b0,s81[40]} + {1'b0,s80[40]};
assign {s91[42],s90[41]} = {1'b0,s82[41]} + {1'b0,s81[41]} + {1'b0,s80[41]};
assign {s91[43],s90[42]} = {1'b0,s82[42]} + {1'b0,s81[42]} + {1'b0,s80[42]};
assign {s91[44],s90[43]} = {1'b0,s82[43]} + {1'b0,s81[43]} + {1'b0,s80[43]};
assign {s91[45],s90[44]} = {1'b0,s82[44]} + {1'b0,s81[44]} + {1'b0,s80[44]};
assign {s91[46],s90[45]} = {1'b0,s82[45]} + {1'b0,s81[45]} + {1'b0,s80[45]};
assign {s91[47],s90[46]} = {1'b0,s82[46]} + {1'b0,s81[46]} + {1'b0,s80[46]};
assign {s91[48],s90[47]} = {1'b0,s82[47]} + {1'b0,s81[47]} + {1'b0,s80[47]};
assign {s91[49],s90[48]} = {1'b0,s82[48]} + {1'b0,s81[48]} + {1'b0,s80[48]};
assign {s91[50],s90[49]} = {1'b0,s82[49]} + {1'b0,s81[49]} + {1'b0,s80[49]};
assign {s91[51],s90[50]} = {1'b0,s82[50]} + {1'b0,s81[50]} + {1'b0,s80[50]};
assign {s91[52],s90[51]} = {1'b0,s82[51]} + {1'b0,s81[51]} + {1'b0,s80[51]};
assign {s91[53],s90[52]} = {1'b0,s82[52]} + {1'b0,s81[52]} + {1'b0,s80[52]};
assign {s91[54],s90[53]} = {1'b0,s82[53]} + {1'b0,s81[53]} + {1'b0,s80[53]};
assign {s91[55],s90[54]} = {1'b0,s82[54]} + {1'b0,s81[54]} + {1'b0,s80[54]};
assign {s91[56],s90[55]} = {1'b0,s82[55]} + {1'b0,s81[55]} + {1'b0,s80[55]};
assign {s91[57],s90[56]} = {1'b0,s82[56]} + {1'b0,s81[56]} + {1'b0,s80[56]};
assign {s91[58],s90[57]} = {1'b0,s82[57]} + {1'b0,s81[57]} + {1'b0,s80[57]};
assign {s91[59],s90[58]} = {1'b0,s82[58]} + {1'b0,s81[58]} + {1'b0,s80[58]};
assign {s91[60],s90[59]} = {1'b0,s82[59]} + {1'b0,s81[59]} + {1'b0,s80[59]};
assign {s91[61],s90[60]} = {1'b0,s82[60]} + {1'b0,s81[60]} + {1'b0,s80[60]};
assign {s91[62],s90[61]} = {1'b0,s82[61]} + {1'b0,s81[61]} + {1'b0,s80[61]};
assign {s91[63],s90[62]} = {1'b0,s82[62]} + {1'b0,s81[62]} + {1'b0,s80[62]};
assign {s91[64],s90[63]} = {1'b0,s82[63]} + {1'b0,s81[63]} + {1'b0,s80[63]};
assign {s91[65],s90[64]} = {1'b0,s82[64]} + {1'b0,s81[64]} + {1'b0,s80[64]};
assign {s91[66],s90[65]} = {1'b0,s82[65]} + {1'b0,s81[65]} + {1'b0,s80[65]};
assign {s91[67],s90[66]} = {1'b0,s82[66]} + {1'b0,s81[66]} + {1'b0,s80[66]};
assign {s93[20],s92[19]} = {1'b0,s83[19]};
assign {s93[21],s92[20]} = {1'b0,s84[20]} + {1'b0,s83[20]};
assign {s93[22],s92[21]} = {1'b0,s84[21]} + {1'b0,s83[21]};
assign {s93[23],s92[22]} = {1'b0,s84[22]} + {1'b0,s83[22]};
assign {s93[24],s92[23]} = {1'b0,s84[23]} + {1'b0,s83[23]};
assign {s93[25],s92[24]} = {1'b0,s84[24]} + {1'b0,s83[24]};
assign {s93[26],s92[25]} = {1'b0,s84[25]} + {1'b0,s83[25]};
assign {s93[27],s92[26]} = {1'b0,s84[26]} + {1'b0,s83[26]};
assign {s93[28],s92[27]} = {1'b0,s85[27]} + {1'b0,s84[27]} + {1'b0,s83[27]};
assign {s93[29],s92[28]} = {1'b0,s85[28]} + {1'b0,s84[28]} + {1'b0,s83[28]};
assign {s93[30],s92[29]} = {1'b0,s85[29]} + {1'b0,s84[29]} + {1'b0,s83[29]};
assign {s93[31],s92[30]} = {1'b0,s85[30]} + {1'b0,s84[30]} + {1'b0,s83[30]};
assign {s93[32],s92[31]} = {1'b0,s85[31]} + {1'b0,s84[31]} + {1'b0,s83[31]};
assign {s93[33],s92[32]} = {1'b0,s85[32]} + {1'b0,s84[32]} + {1'b0,s83[32]};
assign {s93[34],s92[33]} = {1'b0,s85[33]} + {1'b0,s84[33]} + {1'b0,s83[33]};
assign {s93[35],s92[34]} = {1'b0,s85[34]} + {1'b0,s84[34]} + {1'b0,s83[34]};
assign {s93[36],s92[35]} = {1'b0,s85[35]} + {1'b0,s84[35]} + {1'b0,s83[35]};
assign {s93[37],s92[36]} = {1'b0,s85[36]} + {1'b0,s84[36]} + {1'b0,s83[36]};
assign {s93[38],s92[37]} = {1'b0,s85[37]} + {1'b0,s84[37]} + {1'b0,s83[37]};
assign {s93[39],s92[38]} = {1'b0,s85[38]} + {1'b0,s84[38]} + {1'b0,s83[38]};
assign {s93[40],s92[39]} = {1'b0,s85[39]} + {1'b0,s84[39]} + {1'b0,s83[39]};
assign {s93[41],s92[40]} = {1'b0,s85[40]} + {1'b0,s84[40]} + {1'b0,s83[40]};
assign {s93[42],s92[41]} = {1'b0,s85[41]} + {1'b0,s84[41]} + {1'b0,s83[41]};
assign {s93[43],s92[42]} = {1'b0,s85[42]} + {1'b0,s84[42]} + {1'b0,s83[42]};
assign {s93[44],s92[43]} = {1'b0,s85[43]} + {1'b0,s84[43]} + {1'b0,s83[43]};
assign {s93[45],s92[44]} = {1'b0,s85[44]} + {1'b0,s84[44]} + {1'b0,s83[44]};
assign {s93[46],s92[45]} = {1'b0,s85[45]} + {1'b0,s84[45]} + {1'b0,s83[45]};
assign {s93[47],s92[46]} = {1'b0,s85[46]} + {1'b0,s84[46]} + {1'b0,s83[46]};
assign {s93[48],s92[47]} = {1'b0,s85[47]} + {1'b0,s84[47]} + {1'b0,s83[47]};
assign {s93[49],s92[48]} = {1'b0,s85[48]} + {1'b0,s84[48]} + {1'b0,s83[48]};
assign {s93[50],s92[49]} = {1'b0,s85[49]} + {1'b0,s84[49]} + {1'b0,s83[49]};
assign {s93[51],s92[50]} = {1'b0,s85[50]} + {1'b0,s84[50]} + {1'b0,s83[50]};
assign {s93[52],s92[51]} = {1'b0,s85[51]} + {1'b0,s84[51]} + {1'b0,s83[51]};
assign {s93[53],s92[52]} = {1'b0,s85[52]} + {1'b0,s84[52]} + {1'b0,s83[52]};
assign {s93[54],s92[53]} = {1'b0,s85[53]} + {1'b0,s84[53]} + {1'b0,s83[53]};
assign {s93[55],s92[54]} = {1'b0,s85[54]} + {1'b0,s84[54]} + {1'b0,s83[54]};
assign {s93[56],s92[55]} = {1'b0,s85[55]} + {1'b0,s84[55]} + {1'b0,s83[55]};
assign {s93[57],s92[56]} = {1'b0,s85[56]} + {1'b0,s84[56]} + {1'b0,s83[56]};
assign {s93[58],s92[57]} = {1'b0,s85[57]} + {1'b0,s84[57]} + {1'b0,s83[57]};
assign {s93[59],s92[58]} = {1'b0,s85[58]} + {1'b0,s84[58]} + {1'b0,s83[58]};
assign {s93[60],s92[59]} = {1'b0,s85[59]} + {1'b0,s84[59]} + {1'b0,s83[59]};
assign {s93[61],s92[60]} = {1'b0,s85[60]} + {1'b0,s84[60]} + {1'b0,s83[60]};
assign {s93[62],s92[61]} = {1'b0,s85[61]} + {1'b0,s84[61]} + {1'b0,s83[61]};
assign {s93[63],s92[62]} = {1'b0,s85[62]} + {1'b0,s84[62]} + {1'b0,s83[62]};
assign {s93[64],s92[63]} = {1'b0,s85[63]} + {1'b0,s84[63]} + {1'b0,s83[63]};
assign {s93[65],s92[64]} = {1'b0,s85[64]} + {1'b0,s84[64]} + {1'b0,s83[64]};
assign {s93[66],s92[65]} = {1'b0,s85[65]} + {1'b0,s84[65]} + {1'b0,s83[65]};
assign {s93[67],s92[66]} = {1'b0,s85[66]} + {1'b0,s84[66]} + {1'b0,s83[66]};
assign s94 = s86[(PPLEN - 1):28];
assign s95 = s87[(PPLEN - 1):32];
assign {s97[1],s96[0]} = {1'b0,s88[0]};
assign {s97[2],s96[1]} = {1'b0,s89[1]} + {1'b0,s88[1]};
assign {s97[3],s96[2]} = {1'b0,s89[2]} + {1'b0,s88[2]};
assign {s97[4],s96[3]} = {1'b0,s89[3]} + {1'b0,s88[3]};
assign {s97[5],s96[4]} = {1'b0,s89[4]} + {1'b0,s88[4]};
assign {s97[6],s96[5]} = {1'b0,s89[5]} + {1'b0,s88[5]};
assign {s97[7],s96[6]} = {1'b0,s90[6]} + {1'b0,s89[6]} + {1'b0,s88[6]};
assign {s97[8],s96[7]} = {1'b0,s90[7]} + {1'b0,s89[7]} + {1'b0,s88[7]};
assign {s97[9],s96[8]} = {1'b0,s90[8]} + {1'b0,s89[8]} + {1'b0,s88[8]};
assign {s97[10],s96[9]} = {1'b0,s90[9]} + {1'b0,s89[9]} + {1'b0,s88[9]};
assign {s97[11],s96[10]} = {1'b0,s90[10]} + {1'b0,s89[10]} + {1'b0,s88[10]};
assign {s97[12],s96[11]} = {1'b0,s90[11]} + {1'b0,s89[11]} + {1'b0,s88[11]};
assign {s97[13],s96[12]} = {1'b0,s90[12]} + {1'b0,s89[12]} + {1'b0,s88[12]};
assign {s97[14],s96[13]} = {1'b0,s90[13]} + {1'b0,s89[13]} + {1'b0,s88[13]};
assign {s97[15],s96[14]} = {1'b0,s90[14]} + {1'b0,s89[14]} + {1'b0,s88[14]};
assign {s97[16],s96[15]} = {1'b0,s90[15]} + {1'b0,s89[15]} + {1'b0,s88[15]};
assign {s97[17],s96[16]} = {1'b0,s90[16]} + {1'b0,s89[16]} + {1'b0,s88[16]};
assign {s97[18],s96[17]} = {1'b0,s90[17]} + {1'b0,s89[17]} + {1'b0,s88[17]};
assign {s97[19],s96[18]} = {1'b0,s90[18]} + {1'b0,s89[18]} + {1'b0,s88[18]};
assign {s97[20],s96[19]} = {1'b0,s90[19]} + {1'b0,s89[19]} + {1'b0,s88[19]};
assign {s97[21],s96[20]} = {1'b0,s90[20]} + {1'b0,s89[20]} + {1'b0,s88[20]};
assign {s97[22],s96[21]} = {1'b0,s90[21]} + {1'b0,s89[21]} + {1'b0,s88[21]};
assign {s97[23],s96[22]} = {1'b0,s90[22]} + {1'b0,s89[22]} + {1'b0,s88[22]};
assign {s97[24],s96[23]} = {1'b0,s90[23]} + {1'b0,s89[23]} + {1'b0,s88[23]};
assign {s97[25],s96[24]} = {1'b0,s90[24]} + {1'b0,s89[24]} + {1'b0,s88[24]};
assign {s97[26],s96[25]} = {1'b0,s90[25]} + {1'b0,s89[25]} + {1'b0,s88[25]};
assign {s97[27],s96[26]} = {1'b0,s90[26]} + {1'b0,s89[26]} + {1'b0,s88[26]};
assign {s97[28],s96[27]} = {1'b0,s90[27]} + {1'b0,s89[27]} + {1'b0,s88[27]};
assign {s97[29],s96[28]} = {1'b0,s90[28]} + {1'b0,s89[28]} + {1'b0,s88[28]};
assign {s97[30],s96[29]} = {1'b0,s90[29]} + {1'b0,s89[29]} + {1'b0,s88[29]};
assign {s97[31],s96[30]} = {1'b0,s90[30]} + {1'b0,s89[30]} + {1'b0,s88[30]};
assign {s97[32],s96[31]} = {1'b0,s90[31]} + {1'b0,s89[31]} + {1'b0,s88[31]};
assign {s97[33],s96[32]} = {1'b0,s90[32]} + {1'b0,s89[32]} + {1'b0,s88[32]};
assign {s97[34],s96[33]} = {1'b0,s90[33]} + {1'b0,s89[33]} + {1'b0,s88[33]};
assign {s97[35],s96[34]} = {1'b0,s90[34]} + {1'b0,s89[34]} + {1'b0,s88[34]};
assign {s97[36],s96[35]} = {1'b0,s90[35]} + {1'b0,s89[35]} + {1'b0,s88[35]};
assign {s97[37],s96[36]} = {1'b0,s90[36]} + {1'b0,s89[36]} + {1'b0,s88[36]};
assign {s97[38],s96[37]} = {1'b0,s90[37]} + {1'b0,s89[37]} + {1'b0,s88[37]};
assign {s97[39],s96[38]} = {1'b0,s90[38]} + {1'b0,s89[38]} + {1'b0,s88[38]};
assign {s97[40],s96[39]} = {1'b0,s90[39]} + {1'b0,s89[39]} + {1'b0,s88[39]};
assign {s97[41],s96[40]} = {1'b0,s90[40]} + {1'b0,s89[40]} + {1'b0,s88[40]};
assign {s97[42],s96[41]} = {1'b0,s90[41]} + {1'b0,s89[41]} + {1'b0,s88[41]};
assign {s97[43],s96[42]} = {1'b0,s90[42]} + {1'b0,s89[42]} + {1'b0,s88[42]};
assign {s97[44],s96[43]} = {1'b0,s90[43]} + {1'b0,s89[43]} + {1'b0,s88[43]};
assign {s97[45],s96[44]} = {1'b0,s90[44]} + {1'b0,s89[44]} + {1'b0,s88[44]};
assign {s97[46],s96[45]} = {1'b0,s90[45]} + {1'b0,s89[45]} + {1'b0,s88[45]};
assign {s97[47],s96[46]} = {1'b0,s90[46]} + {1'b0,s89[46]} + {1'b0,s88[46]};
assign {s97[48],s96[47]} = {1'b0,s90[47]} + {1'b0,s89[47]} + {1'b0,s88[47]};
assign {s97[49],s96[48]} = {1'b0,s90[48]} + {1'b0,s89[48]} + {1'b0,s88[48]};
assign {s97[50],s96[49]} = {1'b0,s90[49]} + {1'b0,s89[49]} + {1'b0,s88[49]};
assign {s97[51],s96[50]} = {1'b0,s90[50]} + {1'b0,s89[50]} + {1'b0,s88[50]};
assign {s97[52],s96[51]} = {1'b0,s90[51]} + {1'b0,s89[51]} + {1'b0,s88[51]};
assign {s97[53],s96[52]} = {1'b0,s90[52]} + {1'b0,s89[52]} + {1'b0,s88[52]};
assign {s97[54],s96[53]} = {1'b0,s90[53]} + {1'b0,s89[53]} + {1'b0,s88[53]};
assign {s97[55],s96[54]} = {1'b0,s90[54]} + {1'b0,s89[54]} + {1'b0,s88[54]};
assign {s97[56],s96[55]} = {1'b0,s90[55]} + {1'b0,s89[55]} + {1'b0,s88[55]};
assign {s97[57],s96[56]} = {1'b0,s90[56]} + {1'b0,s89[56]} + {1'b0,s88[56]};
assign {s97[58],s96[57]} = {1'b0,s90[57]} + {1'b0,s89[57]} + {1'b0,s88[57]};
assign {s97[59],s96[58]} = {1'b0,s90[58]} + {1'b0,s89[58]} + {1'b0,s88[58]};
assign {s97[60],s96[59]} = {1'b0,s90[59]} + {1'b0,s89[59]} + {1'b0,s88[59]};
assign {s97[61],s96[60]} = {1'b0,s90[60]} + {1'b0,s89[60]} + {1'b0,s88[60]};
assign {s97[62],s96[61]} = {1'b0,s90[61]} + {1'b0,s89[61]} + {1'b0,s88[61]};
assign {s97[63],s96[62]} = {1'b0,s90[62]} + {1'b0,s89[62]} + {1'b0,s88[62]};
assign {s97[64],s96[63]} = {1'b0,s90[63]} + {1'b0,s89[63]} + {1'b0,s88[63]};
assign {s97[65],s96[64]} = {1'b0,s90[64]} + {1'b0,s89[64]} + {1'b0,s88[64]};
assign {s97[66],s96[65]} = {1'b0,s90[65]} + {1'b0,s89[65]} + {1'b0,s88[65]};
assign {s97[67],s96[66]} = {1'b0,s90[66]} + {1'b0,s89[66]} + {1'b0,s88[66]};
assign {s99[8],s98[7]} = {1'b0,s91[7]};
assign {s99[9],s98[8]} = {1'b0,s91[8]};
assign {s99[10],s98[9]} = {1'b0,s91[9]};
assign {s99[11],s98[10]} = {1'b0,s91[10]};
assign {s99[12],s98[11]} = {1'b0,s91[11]};
assign {s99[13],s98[12]} = {1'b0,s91[12]};
assign {s99[14],s98[13]} = {1'b0,s91[13]};
assign {s99[15],s98[14]} = {1'b0,s91[14]};
assign {s99[16],s98[15]} = {1'b0,s91[15]};
assign {s99[17],s98[16]} = {1'b0,s91[16]};
assign {s99[18],s98[17]} = {1'b0,s91[17]};
assign {s99[19],s98[18]} = {1'b0,s91[18]};
assign {s99[20],s98[19]} = {1'b0,s92[19]} + {1'b0,s91[19]};
assign {s99[21],s98[20]} = {1'b0,s93[20]} + {1'b0,s92[20]} + {1'b0,s91[20]};
assign {s99[22],s98[21]} = {1'b0,s93[21]} + {1'b0,s92[21]} + {1'b0,s91[21]};
assign {s99[23],s98[22]} = {1'b0,s93[22]} + {1'b0,s92[22]} + {1'b0,s91[22]};
assign {s99[24],s98[23]} = {1'b0,s93[23]} + {1'b0,s92[23]} + {1'b0,s91[23]};
assign {s99[25],s98[24]} = {1'b0,s93[24]} + {1'b0,s92[24]} + {1'b0,s91[24]};
assign {s99[26],s98[25]} = {1'b0,s93[25]} + {1'b0,s92[25]} + {1'b0,s91[25]};
assign {s99[27],s98[26]} = {1'b0,s93[26]} + {1'b0,s92[26]} + {1'b0,s91[26]};
assign {s99[28],s98[27]} = {1'b0,s93[27]} + {1'b0,s92[27]} + {1'b0,s91[27]};
assign {s99[29],s98[28]} = {1'b0,s93[28]} + {1'b0,s92[28]} + {1'b0,s91[28]};
assign {s99[30],s98[29]} = {1'b0,s93[29]} + {1'b0,s92[29]} + {1'b0,s91[29]};
assign {s99[31],s98[30]} = {1'b0,s93[30]} + {1'b0,s92[30]} + {1'b0,s91[30]};
assign {s99[32],s98[31]} = {1'b0,s93[31]} + {1'b0,s92[31]} + {1'b0,s91[31]};
assign {s99[33],s98[32]} = {1'b0,s93[32]} + {1'b0,s92[32]} + {1'b0,s91[32]};
assign {s99[34],s98[33]} = {1'b0,s93[33]} + {1'b0,s92[33]} + {1'b0,s91[33]};
assign {s99[35],s98[34]} = {1'b0,s93[34]} + {1'b0,s92[34]} + {1'b0,s91[34]};
assign {s99[36],s98[35]} = {1'b0,s93[35]} + {1'b0,s92[35]} + {1'b0,s91[35]};
assign {s99[37],s98[36]} = {1'b0,s93[36]} + {1'b0,s92[36]} + {1'b0,s91[36]};
assign {s99[38],s98[37]} = {1'b0,s93[37]} + {1'b0,s92[37]} + {1'b0,s91[37]};
assign {s99[39],s98[38]} = {1'b0,s93[38]} + {1'b0,s92[38]} + {1'b0,s91[38]};
assign {s99[40],s98[39]} = {1'b0,s93[39]} + {1'b0,s92[39]} + {1'b0,s91[39]};
assign {s99[41],s98[40]} = {1'b0,s93[40]} + {1'b0,s92[40]} + {1'b0,s91[40]};
assign {s99[42],s98[41]} = {1'b0,s93[41]} + {1'b0,s92[41]} + {1'b0,s91[41]};
assign {s99[43],s98[42]} = {1'b0,s93[42]} + {1'b0,s92[42]} + {1'b0,s91[42]};
assign {s99[44],s98[43]} = {1'b0,s93[43]} + {1'b0,s92[43]} + {1'b0,s91[43]};
assign {s99[45],s98[44]} = {1'b0,s93[44]} + {1'b0,s92[44]} + {1'b0,s91[44]};
assign {s99[46],s98[45]} = {1'b0,s93[45]} + {1'b0,s92[45]} + {1'b0,s91[45]};
assign {s99[47],s98[46]} = {1'b0,s93[46]} + {1'b0,s92[46]} + {1'b0,s91[46]};
assign {s99[48],s98[47]} = {1'b0,s93[47]} + {1'b0,s92[47]} + {1'b0,s91[47]};
assign {s99[49],s98[48]} = {1'b0,s93[48]} + {1'b0,s92[48]} + {1'b0,s91[48]};
assign {s99[50],s98[49]} = {1'b0,s93[49]} + {1'b0,s92[49]} + {1'b0,s91[49]};
assign {s99[51],s98[50]} = {1'b0,s93[50]} + {1'b0,s92[50]} + {1'b0,s91[50]};
assign {s99[52],s98[51]} = {1'b0,s93[51]} + {1'b0,s92[51]} + {1'b0,s91[51]};
assign {s99[53],s98[52]} = {1'b0,s93[52]} + {1'b0,s92[52]} + {1'b0,s91[52]};
assign {s99[54],s98[53]} = {1'b0,s93[53]} + {1'b0,s92[53]} + {1'b0,s91[53]};
assign {s99[55],s98[54]} = {1'b0,s93[54]} + {1'b0,s92[54]} + {1'b0,s91[54]};
assign {s99[56],s98[55]} = {1'b0,s93[55]} + {1'b0,s92[55]} + {1'b0,s91[55]};
assign {s99[57],s98[56]} = {1'b0,s93[56]} + {1'b0,s92[56]} + {1'b0,s91[56]};
assign {s99[58],s98[57]} = {1'b0,s93[57]} + {1'b0,s92[57]} + {1'b0,s91[57]};
assign {s99[59],s98[58]} = {1'b0,s93[58]} + {1'b0,s92[58]} + {1'b0,s91[58]};
assign {s99[60],s98[59]} = {1'b0,s93[59]} + {1'b0,s92[59]} + {1'b0,s91[59]};
assign {s99[61],s98[60]} = {1'b0,s93[60]} + {1'b0,s92[60]} + {1'b0,s91[60]};
assign {s99[62],s98[61]} = {1'b0,s93[61]} + {1'b0,s92[61]} + {1'b0,s91[61]};
assign {s99[63],s98[62]} = {1'b0,s93[62]} + {1'b0,s92[62]} + {1'b0,s91[62]};
assign {s99[64],s98[63]} = {1'b0,s93[63]} + {1'b0,s92[63]} + {1'b0,s91[63]};
assign {s99[65],s98[64]} = {1'b0,s93[64]} + {1'b0,s92[64]} + {1'b0,s91[64]};
assign {s99[66],s98[65]} = {1'b0,s93[65]} + {1'b0,s92[65]} + {1'b0,s91[65]};
assign {s99[67],s98[66]} = {1'b0,s93[66]} + {1'b0,s92[66]} + {1'b0,s91[66]};
assign s100 = s94[(PPLEN - 1):28];
assign s101 = s95[(PPLEN - 1):32];
assign {s103[1],s102[0]} = {1'b0,s96[0]};
assign {s103[2],s102[1]} = {1'b0,s97[1]} + {1'b0,s96[1]};
assign {s103[3],s102[2]} = {1'b0,s97[2]} + {1'b0,s96[2]};
assign {s103[4],s102[3]} = {1'b0,s97[3]} + {1'b0,s96[3]};
assign {s103[5],s102[4]} = {1'b0,s97[4]} + {1'b0,s96[4]};
assign {s103[6],s102[5]} = {1'b0,s97[5]} + {1'b0,s96[5]};
assign {s103[7],s102[6]} = {1'b0,s97[6]} + {1'b0,s96[6]};
assign {s103[8],s102[7]} = {1'b0,s98[7]} + {1'b0,s97[7]} + {1'b0,s96[7]};
assign {s103[9],s102[8]} = {1'b0,s98[8]} + {1'b0,s97[8]} + {1'b0,s96[8]};
assign {s103[10],s102[9]} = {1'b0,s98[9]} + {1'b0,s97[9]} + {1'b0,s96[9]};
assign {s103[11],s102[10]} = {1'b0,s98[10]} + {1'b0,s97[10]} + {1'b0,s96[10]};
assign {s103[12],s102[11]} = {1'b0,s98[11]} + {1'b0,s97[11]} + {1'b0,s96[11]};
assign {s103[13],s102[12]} = {1'b0,s98[12]} + {1'b0,s97[12]} + {1'b0,s96[12]};
assign {s103[14],s102[13]} = {1'b0,s98[13]} + {1'b0,s97[13]} + {1'b0,s96[13]};
assign {s103[15],s102[14]} = {1'b0,s98[14]} + {1'b0,s97[14]} + {1'b0,s96[14]};
assign {s103[16],s102[15]} = {1'b0,s98[15]} + {1'b0,s97[15]} + {1'b0,s96[15]};
assign {s103[17],s102[16]} = {1'b0,s98[16]} + {1'b0,s97[16]} + {1'b0,s96[16]};
assign {s103[18],s102[17]} = {1'b0,s98[17]} + {1'b0,s97[17]} + {1'b0,s96[17]};
assign {s103[19],s102[18]} = {1'b0,s98[18]} + {1'b0,s97[18]} + {1'b0,s96[18]};
assign {s103[20],s102[19]} = {1'b0,s98[19]} + {1'b0,s97[19]} + {1'b0,s96[19]};
assign {s103[21],s102[20]} = {1'b0,s98[20]} + {1'b0,s97[20]} + {1'b0,s96[20]};
assign {s103[22],s102[21]} = {1'b0,s98[21]} + {1'b0,s97[21]} + {1'b0,s96[21]};
assign {s103[23],s102[22]} = {1'b0,s98[22]} + {1'b0,s97[22]} + {1'b0,s96[22]};
assign {s103[24],s102[23]} = {1'b0,s98[23]} + {1'b0,s97[23]} + {1'b0,s96[23]};
assign {s103[25],s102[24]} = {1'b0,s98[24]} + {1'b0,s97[24]} + {1'b0,s96[24]};
assign {s103[26],s102[25]} = {1'b0,s98[25]} + {1'b0,s97[25]} + {1'b0,s96[25]};
assign {s103[27],s102[26]} = {1'b0,s98[26]} + {1'b0,s97[26]} + {1'b0,s96[26]};
assign {s103[28],s102[27]} = {1'b0,s98[27]} + {1'b0,s97[27]} + {1'b0,s96[27]};
assign {s103[29],s102[28]} = {1'b0,s98[28]} + {1'b0,s97[28]} + {1'b0,s96[28]};
assign {s103[30],s102[29]} = {1'b0,s98[29]} + {1'b0,s97[29]} + {1'b0,s96[29]};
assign {s103[31],s102[30]} = {1'b0,s98[30]} + {1'b0,s97[30]} + {1'b0,s96[30]};
assign {s103[32],s102[31]} = {1'b0,s98[31]} + {1'b0,s97[31]} + {1'b0,s96[31]};
assign {s103[33],s102[32]} = {1'b0,s98[32]} + {1'b0,s97[32]} + {1'b0,s96[32]};
assign {s103[34],s102[33]} = {1'b0,s98[33]} + {1'b0,s97[33]} + {1'b0,s96[33]};
assign {s103[35],s102[34]} = {1'b0,s98[34]} + {1'b0,s97[34]} + {1'b0,s96[34]};
assign {s103[36],s102[35]} = {1'b0,s98[35]} + {1'b0,s97[35]} + {1'b0,s96[35]};
assign {s103[37],s102[36]} = {1'b0,s98[36]} + {1'b0,s97[36]} + {1'b0,s96[36]};
assign {s103[38],s102[37]} = {1'b0,s98[37]} + {1'b0,s97[37]} + {1'b0,s96[37]};
assign {s103[39],s102[38]} = {1'b0,s98[38]} + {1'b0,s97[38]} + {1'b0,s96[38]};
assign {s103[40],s102[39]} = {1'b0,s98[39]} + {1'b0,s97[39]} + {1'b0,s96[39]};
assign {s103[41],s102[40]} = {1'b0,s98[40]} + {1'b0,s97[40]} + {1'b0,s96[40]};
assign {s103[42],s102[41]} = {1'b0,s98[41]} + {1'b0,s97[41]} + {1'b0,s96[41]};
assign {s103[43],s102[42]} = {1'b0,s98[42]} + {1'b0,s97[42]} + {1'b0,s96[42]};
assign {s103[44],s102[43]} = {1'b0,s98[43]} + {1'b0,s97[43]} + {1'b0,s96[43]};
assign {s103[45],s102[44]} = {1'b0,s98[44]} + {1'b0,s97[44]} + {1'b0,s96[44]};
assign {s103[46],s102[45]} = {1'b0,s98[45]} + {1'b0,s97[45]} + {1'b0,s96[45]};
assign {s103[47],s102[46]} = {1'b0,s98[46]} + {1'b0,s97[46]} + {1'b0,s96[46]};
assign {s103[48],s102[47]} = {1'b0,s98[47]} + {1'b0,s97[47]} + {1'b0,s96[47]};
assign {s103[49],s102[48]} = {1'b0,s98[48]} + {1'b0,s97[48]} + {1'b0,s96[48]};
assign {s103[50],s102[49]} = {1'b0,s98[49]} + {1'b0,s97[49]} + {1'b0,s96[49]};
assign {s103[51],s102[50]} = {1'b0,s98[50]} + {1'b0,s97[50]} + {1'b0,s96[50]};
assign {s103[52],s102[51]} = {1'b0,s98[51]} + {1'b0,s97[51]} + {1'b0,s96[51]};
assign {s103[53],s102[52]} = {1'b0,s98[52]} + {1'b0,s97[52]} + {1'b0,s96[52]};
assign {s103[54],s102[53]} = {1'b0,s98[53]} + {1'b0,s97[53]} + {1'b0,s96[53]};
assign {s103[55],s102[54]} = {1'b0,s98[54]} + {1'b0,s97[54]} + {1'b0,s96[54]};
assign {s103[56],s102[55]} = {1'b0,s98[55]} + {1'b0,s97[55]} + {1'b0,s96[55]};
assign {s103[57],s102[56]} = {1'b0,s98[56]} + {1'b0,s97[56]} + {1'b0,s96[56]};
assign {s103[58],s102[57]} = {1'b0,s98[57]} + {1'b0,s97[57]} + {1'b0,s96[57]};
assign {s103[59],s102[58]} = {1'b0,s98[58]} + {1'b0,s97[58]} + {1'b0,s96[58]};
assign {s103[60],s102[59]} = {1'b0,s98[59]} + {1'b0,s97[59]} + {1'b0,s96[59]};
assign {s103[61],s102[60]} = {1'b0,s98[60]} + {1'b0,s97[60]} + {1'b0,s96[60]};
assign {s103[62],s102[61]} = {1'b0,s98[61]} + {1'b0,s97[61]} + {1'b0,s96[61]};
assign {s103[63],s102[62]} = {1'b0,s98[62]} + {1'b0,s97[62]} + {1'b0,s96[62]};
assign {s103[64],s102[63]} = {1'b0,s98[63]} + {1'b0,s97[63]} + {1'b0,s96[63]};
assign {s103[65],s102[64]} = {1'b0,s98[64]} + {1'b0,s97[64]} + {1'b0,s96[64]};
assign {s103[66],s102[65]} = {1'b0,s98[65]} + {1'b0,s97[65]} + {1'b0,s96[65]};
assign {s103[67],s102[66]} = {1'b0,s98[66]} + {1'b0,s97[66]} + {1'b0,s96[66]};
assign {s105[9],s104[8]} = {1'b0,s99[8]};
assign {s105[10],s104[9]} = {1'b0,s99[9]};
assign {s105[11],s104[10]} = {1'b0,s99[10]};
assign {s105[12],s104[11]} = {1'b0,s99[11]};
assign {s105[13],s104[12]} = {1'b0,s99[12]};
assign {s105[14],s104[13]} = {1'b0,s99[13]};
assign {s105[15],s104[14]} = {1'b0,s99[14]};
assign {s105[16],s104[15]} = {1'b0,s99[15]};
assign {s105[17],s104[16]} = {1'b0,s99[16]};
assign {s105[18],s104[17]} = {1'b0,s99[17]};
assign {s105[19],s104[18]} = {1'b0,s99[18]};
assign {s105[20],s104[19]} = {1'b0,s99[19]};
assign {s105[21],s104[20]} = {1'b0,s99[20]};
assign {s105[22],s104[21]} = {1'b0,s99[21]};
assign {s105[23],s104[22]} = {1'b0,s99[22]};
assign {s105[24],s104[23]} = {1'b0,s99[23]};
assign {s105[25],s104[24]} = {1'b0,s99[24]};
assign {s105[26],s104[25]} = {1'b0,s99[25]};
assign {s105[27],s104[26]} = {1'b0,s99[26]};
assign {s105[28],s104[27]} = {1'b0,s99[27]};
assign {s105[29],s104[28]} = {1'b0,s100[28]} + {1'b0,s99[28]};
assign {s105[30],s104[29]} = {1'b0,s100[29]} + {1'b0,s99[29]};
assign {s105[31],s104[30]} = {1'b0,s100[30]} + {1'b0,s99[30]};
assign {s105[32],s104[31]} = {1'b0,s100[31]} + {1'b0,s99[31]};
assign {s105[33],s104[32]} = {1'b0,s101[32]} + {1'b0,s100[32]} + {1'b0,s99[32]};
assign {s105[34],s104[33]} = {1'b0,s101[33]} + {1'b0,s100[33]} + {1'b0,s99[33]};
assign {s105[35],s104[34]} = {1'b0,s101[34]} + {1'b0,s100[34]} + {1'b0,s99[34]};
assign {s105[36],s104[35]} = {1'b0,s101[35]} + {1'b0,s100[35]} + {1'b0,s99[35]};
assign {s105[37],s104[36]} = {1'b0,s101[36]} + {1'b0,s100[36]} + {1'b0,s99[36]};
assign {s105[38],s104[37]} = {1'b0,s101[37]} + {1'b0,s100[37]} + {1'b0,s99[37]};
assign {s105[39],s104[38]} = {1'b0,s101[38]} + {1'b0,s100[38]} + {1'b0,s99[38]};
assign {s105[40],s104[39]} = {1'b0,s101[39]} + {1'b0,s100[39]} + {1'b0,s99[39]};
assign {s105[41],s104[40]} = {1'b0,s101[40]} + {1'b0,s100[40]} + {1'b0,s99[40]};
assign {s105[42],s104[41]} = {1'b0,s101[41]} + {1'b0,s100[41]} + {1'b0,s99[41]};
assign {s105[43],s104[42]} = {1'b0,s101[42]} + {1'b0,s100[42]} + {1'b0,s99[42]};
assign {s105[44],s104[43]} = {1'b0,s101[43]} + {1'b0,s100[43]} + {1'b0,s99[43]};
assign {s105[45],s104[44]} = {1'b0,s101[44]} + {1'b0,s100[44]} + {1'b0,s99[44]};
assign {s105[46],s104[45]} = {1'b0,s101[45]} + {1'b0,s100[45]} + {1'b0,s99[45]};
assign {s105[47],s104[46]} = {1'b0,s101[46]} + {1'b0,s100[46]} + {1'b0,s99[46]};
assign {s105[48],s104[47]} = {1'b0,s101[47]} + {1'b0,s100[47]} + {1'b0,s99[47]};
assign {s105[49],s104[48]} = {1'b0,s101[48]} + {1'b0,s100[48]} + {1'b0,s99[48]};
assign {s105[50],s104[49]} = {1'b0,s101[49]} + {1'b0,s100[49]} + {1'b0,s99[49]};
assign {s105[51],s104[50]} = {1'b0,s101[50]} + {1'b0,s100[50]} + {1'b0,s99[50]};
assign {s105[52],s104[51]} = {1'b0,s101[51]} + {1'b0,s100[51]} + {1'b0,s99[51]};
assign {s105[53],s104[52]} = {1'b0,s101[52]} + {1'b0,s100[52]} + {1'b0,s99[52]};
assign {s105[54],s104[53]} = {1'b0,s101[53]} + {1'b0,s100[53]} + {1'b0,s99[53]};
assign {s105[55],s104[54]} = {1'b0,s101[54]} + {1'b0,s100[54]} + {1'b0,s99[54]};
assign {s105[56],s104[55]} = {1'b0,s101[55]} + {1'b0,s100[55]} + {1'b0,s99[55]};
assign {s105[57],s104[56]} = {1'b0,s101[56]} + {1'b0,s100[56]} + {1'b0,s99[56]};
assign {s105[58],s104[57]} = {1'b0,s101[57]} + {1'b0,s100[57]} + {1'b0,s99[57]};
assign {s105[59],s104[58]} = {1'b0,s101[58]} + {1'b0,s100[58]} + {1'b0,s99[58]};
assign {s105[60],s104[59]} = {1'b0,s101[59]} + {1'b0,s100[59]} + {1'b0,s99[59]};
assign {s105[61],s104[60]} = {1'b0,s101[60]} + {1'b0,s100[60]} + {1'b0,s99[60]};
assign {s105[62],s104[61]} = {1'b0,s101[61]} + {1'b0,s100[61]} + {1'b0,s99[61]};
assign {s105[63],s104[62]} = {1'b0,s101[62]} + {1'b0,s100[62]} + {1'b0,s99[62]};
assign {s105[64],s104[63]} = {1'b0,s101[63]} + {1'b0,s100[63]} + {1'b0,s99[63]};
assign {s105[65],s104[64]} = {1'b0,s101[64]} + {1'b0,s100[64]} + {1'b0,s99[64]};
assign {s105[66],s104[65]} = {1'b0,s101[65]} + {1'b0,s100[65]} + {1'b0,s99[65]};
assign {s105[67],s104[66]} = {1'b0,s101[66]} + {1'b0,s100[66]} + {1'b0,s99[66]};
assign {s107[1],s106[0]} = {1'b0,s102[0]};
assign {s107[2],s106[1]} = {1'b0,s103[1]} + {1'b0,s102[1]};
assign {s107[3],s106[2]} = {1'b0,s103[2]} + {1'b0,s102[2]};
assign {s107[4],s106[3]} = {1'b0,s103[3]} + {1'b0,s102[3]};
assign {s107[5],s106[4]} = {1'b0,s103[4]} + {1'b0,s102[4]};
assign {s107[6],s106[5]} = {1'b0,s103[5]} + {1'b0,s102[5]};
assign {s107[7],s106[6]} = {1'b0,s103[6]} + {1'b0,s102[6]};
assign {s107[8],s106[7]} = {1'b0,s103[7]} + {1'b0,s102[7]};
assign {s107[9],s106[8]} = {1'b0,s104[8]} + {1'b0,s103[8]} + {1'b0,s102[8]};
assign {s107[10],s106[9]} = {1'b0,s104[9]} + {1'b0,s103[9]} + {1'b0,s102[9]};
assign {s107[11],s106[10]} = {1'b0,s104[10]} + {1'b0,s103[10]} + {1'b0,s102[10]};
assign {s107[12],s106[11]} = {1'b0,s104[11]} + {1'b0,s103[11]} + {1'b0,s102[11]};
assign {s107[13],s106[12]} = {1'b0,s104[12]} + {1'b0,s103[12]} + {1'b0,s102[12]};
assign {s107[14],s106[13]} = {1'b0,s104[13]} + {1'b0,s103[13]} + {1'b0,s102[13]};
assign {s107[15],s106[14]} = {1'b0,s104[14]} + {1'b0,s103[14]} + {1'b0,s102[14]};
assign {s107[16],s106[15]} = {1'b0,s104[15]} + {1'b0,s103[15]} + {1'b0,s102[15]};
assign {s107[17],s106[16]} = {1'b0,s104[16]} + {1'b0,s103[16]} + {1'b0,s102[16]};
assign {s107[18],s106[17]} = {1'b0,s104[17]} + {1'b0,s103[17]} + {1'b0,s102[17]};
assign {s107[19],s106[18]} = {1'b0,s104[18]} + {1'b0,s103[18]} + {1'b0,s102[18]};
assign {s107[20],s106[19]} = {1'b0,s104[19]} + {1'b0,s103[19]} + {1'b0,s102[19]};
assign {s107[21],s106[20]} = {1'b0,s104[20]} + {1'b0,s103[20]} + {1'b0,s102[20]};
assign {s107[22],s106[21]} = {1'b0,s104[21]} + {1'b0,s103[21]} + {1'b0,s102[21]};
assign {s107[23],s106[22]} = {1'b0,s104[22]} + {1'b0,s103[22]} + {1'b0,s102[22]};
assign {s107[24],s106[23]} = {1'b0,s104[23]} + {1'b0,s103[23]} + {1'b0,s102[23]};
assign {s107[25],s106[24]} = {1'b0,s104[24]} + {1'b0,s103[24]} + {1'b0,s102[24]};
assign {s107[26],s106[25]} = {1'b0,s104[25]} + {1'b0,s103[25]} + {1'b0,s102[25]};
assign {s107[27],s106[26]} = {1'b0,s104[26]} + {1'b0,s103[26]} + {1'b0,s102[26]};
assign {s107[28],s106[27]} = {1'b0,s104[27]} + {1'b0,s103[27]} + {1'b0,s102[27]};
assign {s107[29],s106[28]} = {1'b0,s104[28]} + {1'b0,s103[28]} + {1'b0,s102[28]};
assign {s107[30],s106[29]} = {1'b0,s104[29]} + {1'b0,s103[29]} + {1'b0,s102[29]};
assign {s107[31],s106[30]} = {1'b0,s104[30]} + {1'b0,s103[30]} + {1'b0,s102[30]};
assign {s107[32],s106[31]} = {1'b0,s104[31]} + {1'b0,s103[31]} + {1'b0,s102[31]};
assign {s107[33],s106[32]} = {1'b0,s104[32]} + {1'b0,s103[32]} + {1'b0,s102[32]};
assign {s107[34],s106[33]} = {1'b0,s104[33]} + {1'b0,s103[33]} + {1'b0,s102[33]};
assign {s107[35],s106[34]} = {1'b0,s104[34]} + {1'b0,s103[34]} + {1'b0,s102[34]};
assign {s107[36],s106[35]} = {1'b0,s104[35]} + {1'b0,s103[35]} + {1'b0,s102[35]};
assign {s107[37],s106[36]} = {1'b0,s104[36]} + {1'b0,s103[36]} + {1'b0,s102[36]};
assign {s107[38],s106[37]} = {1'b0,s104[37]} + {1'b0,s103[37]} + {1'b0,s102[37]};
assign {s107[39],s106[38]} = {1'b0,s104[38]} + {1'b0,s103[38]} + {1'b0,s102[38]};
assign {s107[40],s106[39]} = {1'b0,s104[39]} + {1'b0,s103[39]} + {1'b0,s102[39]};
assign {s107[41],s106[40]} = {1'b0,s104[40]} + {1'b0,s103[40]} + {1'b0,s102[40]};
assign {s107[42],s106[41]} = {1'b0,s104[41]} + {1'b0,s103[41]} + {1'b0,s102[41]};
assign {s107[43],s106[42]} = {1'b0,s104[42]} + {1'b0,s103[42]} + {1'b0,s102[42]};
assign {s107[44],s106[43]} = {1'b0,s104[43]} + {1'b0,s103[43]} + {1'b0,s102[43]};
assign {s107[45],s106[44]} = {1'b0,s104[44]} + {1'b0,s103[44]} + {1'b0,s102[44]};
assign {s107[46],s106[45]} = {1'b0,s104[45]} + {1'b0,s103[45]} + {1'b0,s102[45]};
assign {s107[47],s106[46]} = {1'b0,s104[46]} + {1'b0,s103[46]} + {1'b0,s102[46]};
assign {s107[48],s106[47]} = {1'b0,s104[47]} + {1'b0,s103[47]} + {1'b0,s102[47]};
assign {s107[49],s106[48]} = {1'b0,s104[48]} + {1'b0,s103[48]} + {1'b0,s102[48]};
assign {s107[50],s106[49]} = {1'b0,s104[49]} + {1'b0,s103[49]} + {1'b0,s102[49]};
assign {s107[51],s106[50]} = {1'b0,s104[50]} + {1'b0,s103[50]} + {1'b0,s102[50]};
assign {s107[52],s106[51]} = {1'b0,s104[51]} + {1'b0,s103[51]} + {1'b0,s102[51]};
assign {s107[53],s106[52]} = {1'b0,s104[52]} + {1'b0,s103[52]} + {1'b0,s102[52]};
assign {s107[54],s106[53]} = {1'b0,s104[53]} + {1'b0,s103[53]} + {1'b0,s102[53]};
assign {s107[55],s106[54]} = {1'b0,s104[54]} + {1'b0,s103[54]} + {1'b0,s102[54]};
assign {s107[56],s106[55]} = {1'b0,s104[55]} + {1'b0,s103[55]} + {1'b0,s102[55]};
assign {s107[57],s106[56]} = {1'b0,s104[56]} + {1'b0,s103[56]} + {1'b0,s102[56]};
assign {s107[58],s106[57]} = {1'b0,s104[57]} + {1'b0,s103[57]} + {1'b0,s102[57]};
assign {s107[59],s106[58]} = {1'b0,s104[58]} + {1'b0,s103[58]} + {1'b0,s102[58]};
assign {s107[60],s106[59]} = {1'b0,s104[59]} + {1'b0,s103[59]} + {1'b0,s102[59]};
assign {s107[61],s106[60]} = {1'b0,s104[60]} + {1'b0,s103[60]} + {1'b0,s102[60]};
assign {s107[62],s106[61]} = {1'b0,s104[61]} + {1'b0,s103[61]} + {1'b0,s102[61]};
assign {s107[63],s106[62]} = {1'b0,s104[62]} + {1'b0,s103[62]} + {1'b0,s102[62]};
assign {s107[64],s106[63]} = {1'b0,s104[63]} + {1'b0,s103[63]} + {1'b0,s102[63]};
assign {s107[65],s106[64]} = {1'b0,s104[64]} + {1'b0,s103[64]} + {1'b0,s102[64]};
assign {s107[66],s106[65]} = {1'b0,s104[65]} + {1'b0,s103[65]} + {1'b0,s102[65]};
assign {s107[67],s106[66]} = {1'b0,s104[66]} + {1'b0,s103[66]} + {1'b0,s102[66]};
assign s108 = s105[(PPLEN - 1):9];
assign {s110[1],s109[0]} = {1'b0,s106[0]};
assign {s110[2],s109[1]} = {1'b0,s107[1]} + {1'b0,s106[1]};
assign {s110[3],s109[2]} = {1'b0,s107[2]} + {1'b0,s106[2]};
assign {s110[4],s109[3]} = {1'b0,s107[3]} + {1'b0,s106[3]};
assign {s110[5],s109[4]} = {1'b0,s107[4]} + {1'b0,s106[4]};
assign {s110[6],s109[5]} = {1'b0,s107[5]} + {1'b0,s106[5]};
assign {s110[7],s109[6]} = {1'b0,s107[6]} + {1'b0,s106[6]};
assign {s110[8],s109[7]} = {1'b0,s107[7]} + {1'b0,s106[7]};
assign {s110[9],s109[8]} = {1'b0,s107[8]} + {1'b0,s106[8]};
assign {s110[10],s109[9]} = {1'b0,s108[9]} + {1'b0,s107[9]} + {1'b0,s106[9]};
assign {s110[11],s109[10]} = {1'b0,s108[10]} + {1'b0,s107[10]} + {1'b0,s106[10]};
assign {s110[12],s109[11]} = {1'b0,s108[11]} + {1'b0,s107[11]} + {1'b0,s106[11]};
assign {s110[13],s109[12]} = {1'b0,s108[12]} + {1'b0,s107[12]} + {1'b0,s106[12]};
assign {s110[14],s109[13]} = {1'b0,s108[13]} + {1'b0,s107[13]} + {1'b0,s106[13]};
assign {s110[15],s109[14]} = {1'b0,s108[14]} + {1'b0,s107[14]} + {1'b0,s106[14]};
assign {s110[16],s109[15]} = {1'b0,s108[15]} + {1'b0,s107[15]} + {1'b0,s106[15]};
assign {s110[17],s109[16]} = {1'b0,s108[16]} + {1'b0,s107[16]} + {1'b0,s106[16]};
assign {s110[18],s109[17]} = {1'b0,s108[17]} + {1'b0,s107[17]} + {1'b0,s106[17]};
assign {s110[19],s109[18]} = {1'b0,s108[18]} + {1'b0,s107[18]} + {1'b0,s106[18]};
assign {s110[20],s109[19]} = {1'b0,s108[19]} + {1'b0,s107[19]} + {1'b0,s106[19]};
assign {s110[21],s109[20]} = {1'b0,s108[20]} + {1'b0,s107[20]} + {1'b0,s106[20]};
assign {s110[22],s109[21]} = {1'b0,s108[21]} + {1'b0,s107[21]} + {1'b0,s106[21]};
assign {s110[23],s109[22]} = {1'b0,s108[22]} + {1'b0,s107[22]} + {1'b0,s106[22]};
assign {s110[24],s109[23]} = {1'b0,s108[23]} + {1'b0,s107[23]} + {1'b0,s106[23]};
assign {s110[25],s109[24]} = {1'b0,s108[24]} + {1'b0,s107[24]} + {1'b0,s106[24]};
assign {s110[26],s109[25]} = {1'b0,s108[25]} + {1'b0,s107[25]} + {1'b0,s106[25]};
assign {s110[27],s109[26]} = {1'b0,s108[26]} + {1'b0,s107[26]} + {1'b0,s106[26]};
assign {s110[28],s109[27]} = {1'b0,s108[27]} + {1'b0,s107[27]} + {1'b0,s106[27]};
assign {s110[29],s109[28]} = {1'b0,s108[28]} + {1'b0,s107[28]} + {1'b0,s106[28]};
assign {s110[30],s109[29]} = {1'b0,s108[29]} + {1'b0,s107[29]} + {1'b0,s106[29]};
assign {s110[31],s109[30]} = {1'b0,s108[30]} + {1'b0,s107[30]} + {1'b0,s106[30]};
assign {s110[32],s109[31]} = {1'b0,s108[31]} + {1'b0,s107[31]} + {1'b0,s106[31]};
assign {s110[33],s109[32]} = {1'b0,s108[32]} + {1'b0,s107[32]} + {1'b0,s106[32]};
assign {s110[34],s109[33]} = {1'b0,s108[33]} + {1'b0,s107[33]} + {1'b0,s106[33]};
assign {s110[35],s109[34]} = {1'b0,s108[34]} + {1'b0,s107[34]} + {1'b0,s106[34]};
assign {s110[36],s109[35]} = {1'b0,s108[35]} + {1'b0,s107[35]} + {1'b0,s106[35]};
assign {s110[37],s109[36]} = {1'b0,s108[36]} + {1'b0,s107[36]} + {1'b0,s106[36]};
assign {s110[38],s109[37]} = {1'b0,s108[37]} + {1'b0,s107[37]} + {1'b0,s106[37]};
assign {s110[39],s109[38]} = {1'b0,s108[38]} + {1'b0,s107[38]} + {1'b0,s106[38]};
assign {s110[40],s109[39]} = {1'b0,s108[39]} + {1'b0,s107[39]} + {1'b0,s106[39]};
assign {s110[41],s109[40]} = {1'b0,s108[40]} + {1'b0,s107[40]} + {1'b0,s106[40]};
assign {s110[42],s109[41]} = {1'b0,s108[41]} + {1'b0,s107[41]} + {1'b0,s106[41]};
assign {s110[43],s109[42]} = {1'b0,s108[42]} + {1'b0,s107[42]} + {1'b0,s106[42]};
assign {s110[44],s109[43]} = {1'b0,s108[43]} + {1'b0,s107[43]} + {1'b0,s106[43]};
assign {s110[45],s109[44]} = {1'b0,s108[44]} + {1'b0,s107[44]} + {1'b0,s106[44]};
assign {s110[46],s109[45]} = {1'b0,s108[45]} + {1'b0,s107[45]} + {1'b0,s106[45]};
assign {s110[47],s109[46]} = {1'b0,s108[46]} + {1'b0,s107[46]} + {1'b0,s106[46]};
assign {s110[48],s109[47]} = {1'b0,s108[47]} + {1'b0,s107[47]} + {1'b0,s106[47]};
assign {s110[49],s109[48]} = {1'b0,s108[48]} + {1'b0,s107[48]} + {1'b0,s106[48]};
assign {s110[50],s109[49]} = {1'b0,s108[49]} + {1'b0,s107[49]} + {1'b0,s106[49]};
assign {s110[51],s109[50]} = {1'b0,s108[50]} + {1'b0,s107[50]} + {1'b0,s106[50]};
assign {s110[52],s109[51]} = {1'b0,s108[51]} + {1'b0,s107[51]} + {1'b0,s106[51]};
assign {s110[53],s109[52]} = {1'b0,s108[52]} + {1'b0,s107[52]} + {1'b0,s106[52]};
assign {s110[54],s109[53]} = {1'b0,s108[53]} + {1'b0,s107[53]} + {1'b0,s106[53]};
assign {s110[55],s109[54]} = {1'b0,s108[54]} + {1'b0,s107[54]} + {1'b0,s106[54]};
assign {s110[56],s109[55]} = {1'b0,s108[55]} + {1'b0,s107[55]} + {1'b0,s106[55]};
assign {s110[57],s109[56]} = {1'b0,s108[56]} + {1'b0,s107[56]} + {1'b0,s106[56]};
assign {s110[58],s109[57]} = {1'b0,s108[57]} + {1'b0,s107[57]} + {1'b0,s106[57]};
assign {s110[59],s109[58]} = {1'b0,s108[58]} + {1'b0,s107[58]} + {1'b0,s106[58]};
assign {s110[60],s109[59]} = {1'b0,s108[59]} + {1'b0,s107[59]} + {1'b0,s106[59]};
assign {s110[61],s109[60]} = {1'b0,s108[60]} + {1'b0,s107[60]} + {1'b0,s106[60]};
assign {s110[62],s109[61]} = {1'b0,s108[61]} + {1'b0,s107[61]} + {1'b0,s106[61]};
assign {s110[63],s109[62]} = {1'b0,s108[62]} + {1'b0,s107[62]} + {1'b0,s106[62]};
assign {s110[64],s109[63]} = {1'b0,s108[63]} + {1'b0,s107[63]} + {1'b0,s106[63]};
assign {s110[65],s109[64]} = {1'b0,s108[64]} + {1'b0,s107[64]} + {1'b0,s106[64]};
assign {s110[66],s109[65]} = {1'b0,s108[65]} + {1'b0,s107[65]} + {1'b0,s106[65]};
assign {s110[67],s109[66]} = {1'b0,s108[66]} + {1'b0,s107[66]} + {1'b0,s106[66]};
assign mul_wt_sum = s109[PPLEN - 1:0];
assign mul_wt_cout = {s110[PPLEN - 1:1],1'b0};
endmodule

