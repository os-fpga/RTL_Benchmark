library ieee;
use ieee.std_logic_1164.all;


entity top is
	 port(A: in std_logic_vector(127 downto 0);
	  P: out std_logic_vector(6 downto 0);
	  F: out std_logic);
 end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977: std_logic;

begin

w0 <= not A(125) and A(127);
w1 <= A(126) and A(127);
w2 <= A(126) and not w1;
w3 <= A(125) and not w2;
w4 <= not w0 and not w3;
w5 <= not A(123) and not w4;
w6 <= not A(124) and not w2;
w7 <= A(124) and not w4;
w8 <= not w6 and not w7;
w9 <= A(123) and not w8;
w10 <= not w5 and not w9;
w11 <= not A(121) and not w10;
w12 <= not A(122) and not w8;
w13 <= A(122) and not w10;
w14 <= not w12 and not w13;
w15 <= A(121) and not w14;
w16 <= not w11 and not w15;
w17 <= not A(119) and not w16;
w18 <= not A(120) and not w14;
w19 <= A(120) and not w16;
w20 <= not w18 and not w19;
w21 <= A(119) and not w20;
w22 <= not w17 and not w21;
w23 <= not A(117) and not w22;
w24 <= not A(118) and not w20;
w25 <= A(118) and not w22;
w26 <= not w24 and not w25;
w27 <= A(117) and not w26;
w28 <= not w23 and not w27;
w29 <= not A(115) and not w28;
w30 <= not A(116) and not w26;
w31 <= A(116) and not w28;
w32 <= not w30 and not w31;
w33 <= A(115) and not w32;
w34 <= not w29 and not w33;
w35 <= not A(113) and not w34;
w36 <= not A(114) and not w32;
w37 <= A(114) and not w34;
w38 <= not w36 and not w37;
w39 <= A(113) and not w38;
w40 <= not w35 and not w39;
w41 <= not A(111) and not w40;
w42 <= not A(112) and not w38;
w43 <= A(112) and not w40;
w44 <= not w42 and not w43;
w45 <= A(111) and not w44;
w46 <= not w41 and not w45;
w47 <= not A(109) and not w46;
w48 <= not A(110) and not w44;
w49 <= A(110) and not w46;
w50 <= not w48 and not w49;
w51 <= A(109) and not w50;
w52 <= not w47 and not w51;
w53 <= not A(107) and not w52;
w54 <= not A(108) and not w50;
w55 <= A(108) and not w52;
w56 <= not w54 and not w55;
w57 <= A(107) and not w56;
w58 <= not w53 and not w57;
w59 <= not A(105) and not w58;
w60 <= not A(106) and not w56;
w61 <= A(106) and not w58;
w62 <= not w60 and not w61;
w63 <= A(105) and not w62;
w64 <= not w59 and not w63;
w65 <= not A(103) and not w64;
w66 <= not A(104) and not w62;
w67 <= A(104) and not w64;
w68 <= not w66 and not w67;
w69 <= A(103) and not w68;
w70 <= not w65 and not w69;
w71 <= not A(101) and not w70;
w72 <= not A(102) and not w68;
w73 <= A(102) and not w70;
w74 <= not w72 and not w73;
w75 <= A(101) and not w74;
w76 <= not w71 and not w75;
w77 <= not A(99) and not w76;
w78 <= not A(100) and not w74;
w79 <= A(100) and not w76;
w80 <= not w78 and not w79;
w81 <= A(99) and not w80;
w82 <= not w77 and not w81;
w83 <= not A(97) and not w82;
w84 <= not A(98) and not w80;
w85 <= A(98) and not w82;
w86 <= not w84 and not w85;
w87 <= A(97) and not w86;
w88 <= not w83 and not w87;
w89 <= not A(95) and not w88;
w90 <= not A(96) and not w86;
w91 <= A(96) and not w88;
w92 <= not w90 and not w91;
w93 <= A(95) and not w92;
w94 <= not w89 and not w93;
w95 <= not A(93) and not w94;
w96 <= not A(94) and not w92;
w97 <= A(94) and not w94;
w98 <= not w96 and not w97;
w99 <= A(93) and not w98;
w100 <= not w95 and not w99;
w101 <= not A(91) and not w100;
w102 <= not A(92) and not w98;
w103 <= A(92) and not w100;
w104 <= not w102 and not w103;
w105 <= A(91) and not w104;
w106 <= not w101 and not w105;
w107 <= not A(89) and not w106;
w108 <= not A(90) and not w104;
w109 <= A(90) and not w106;
w110 <= not w108 and not w109;
w111 <= A(89) and not w110;
w112 <= not w107 and not w111;
w113 <= not A(87) and not w112;
w114 <= not A(88) and not w110;
w115 <= A(88) and not w112;
w116 <= not w114 and not w115;
w117 <= A(87) and not w116;
w118 <= not w113 and not w117;
w119 <= not A(85) and not w118;
w120 <= not A(86) and not w116;
w121 <= A(86) and not w118;
w122 <= not w120 and not w121;
w123 <= A(85) and not w122;
w124 <= not w119 and not w123;
w125 <= not A(83) and not w124;
w126 <= not A(84) and not w122;
w127 <= A(84) and not w124;
w128 <= not w126 and not w127;
w129 <= A(83) and not w128;
w130 <= not w125 and not w129;
w131 <= not A(81) and not w130;
w132 <= not A(82) and not w128;
w133 <= A(82) and not w130;
w134 <= not w132 and not w133;
w135 <= A(81) and not w134;
w136 <= not w131 and not w135;
w137 <= not A(79) and not w136;
w138 <= not A(80) and not w134;
w139 <= A(80) and not w136;
w140 <= not w138 and not w139;
w141 <= A(79) and not w140;
w142 <= not w137 and not w141;
w143 <= not A(77) and not w142;
w144 <= not A(78) and not w140;
w145 <= A(78) and not w142;
w146 <= not w144 and not w145;
w147 <= A(77) and not w146;
w148 <= not w143 and not w147;
w149 <= not A(75) and not w148;
w150 <= not A(76) and not w146;
w151 <= A(76) and not w148;
w152 <= not w150 and not w151;
w153 <= A(75) and not w152;
w154 <= not w149 and not w153;
w155 <= not A(73) and not w154;
w156 <= not A(74) and not w152;
w157 <= A(74) and not w154;
w158 <= not w156 and not w157;
w159 <= A(73) and not w158;
w160 <= not w155 and not w159;
w161 <= not A(71) and not w160;
w162 <= not A(72) and not w158;
w163 <= A(72) and not w160;
w164 <= not w162 and not w163;
w165 <= A(71) and not w164;
w166 <= not w161 and not w165;
w167 <= not A(69) and not w166;
w168 <= not A(70) and not w164;
w169 <= A(70) and not w166;
w170 <= not w168 and not w169;
w171 <= A(69) and not w170;
w172 <= not w167 and not w171;
w173 <= not A(67) and not w172;
w174 <= not A(68) and not w170;
w175 <= A(68) and not w172;
w176 <= not w174 and not w175;
w177 <= A(67) and not w176;
w178 <= not w173 and not w177;
w179 <= not A(65) and not w178;
w180 <= not A(66) and not w176;
w181 <= A(66) and not w178;
w182 <= not w180 and not w181;
w183 <= A(65) and not w182;
w184 <= not w179 and not w183;
w185 <= not A(63) and not w184;
w186 <= not A(64) and not w182;
w187 <= A(64) and not w184;
w188 <= not w186 and not w187;
w189 <= A(63) and not w188;
w190 <= not w185 and not w189;
w191 <= not A(61) and not w190;
w192 <= not A(62) and not w188;
w193 <= A(62) and not w190;
w194 <= not w192 and not w193;
w195 <= A(61) and not w194;
w196 <= not w191 and not w195;
w197 <= not A(59) and not w196;
w198 <= not A(60) and not w194;
w199 <= A(60) and not w196;
w200 <= not w198 and not w199;
w201 <= A(59) and not w200;
w202 <= not w197 and not w201;
w203 <= not A(57) and not w202;
w204 <= not A(58) and not w200;
w205 <= A(58) and not w202;
w206 <= not w204 and not w205;
w207 <= A(57) and not w206;
w208 <= not w203 and not w207;
w209 <= not A(55) and not w208;
w210 <= not A(56) and not w206;
w211 <= A(56) and not w208;
w212 <= not w210 and not w211;
w213 <= A(55) and not w212;
w214 <= not w209 and not w213;
w215 <= not A(53) and not w214;
w216 <= not A(54) and not w212;
w217 <= A(54) and not w214;
w218 <= not w216 and not w217;
w219 <= A(53) and not w218;
w220 <= not w215 and not w219;
w221 <= not A(51) and not w220;
w222 <= not A(52) and not w218;
w223 <= A(52) and not w220;
w224 <= not w222 and not w223;
w225 <= A(51) and not w224;
w226 <= not w221 and not w225;
w227 <= not A(49) and not w226;
w228 <= not A(50) and not w224;
w229 <= A(50) and not w226;
w230 <= not w228 and not w229;
w231 <= A(49) and not w230;
w232 <= not w227 and not w231;
w233 <= not A(47) and not w232;
w234 <= not A(48) and not w230;
w235 <= A(48) and not w232;
w236 <= not w234 and not w235;
w237 <= A(47) and not w236;
w238 <= not w233 and not w237;
w239 <= not A(45) and not w238;
w240 <= not A(46) and not w236;
w241 <= A(46) and not w238;
w242 <= not w240 and not w241;
w243 <= A(45) and not w242;
w244 <= not w239 and not w243;
w245 <= not A(43) and not w244;
w246 <= not A(44) and not w242;
w247 <= A(44) and not w244;
w248 <= not w246 and not w247;
w249 <= A(43) and not w248;
w250 <= not w245 and not w249;
w251 <= not A(41) and not w250;
w252 <= not A(42) and not w248;
w253 <= A(42) and not w250;
w254 <= not w252 and not w253;
w255 <= A(41) and not w254;
w256 <= not w251 and not w255;
w257 <= not A(39) and not w256;
w258 <= not A(40) and not w254;
w259 <= A(40) and not w256;
w260 <= not w258 and not w259;
w261 <= A(39) and not w260;
w262 <= not w257 and not w261;
w263 <= not A(37) and not w262;
w264 <= not A(38) and not w260;
w265 <= A(38) and not w262;
w266 <= not w264 and not w265;
w267 <= A(37) and not w266;
w268 <= not w263 and not w267;
w269 <= not A(35) and not w268;
w270 <= not A(36) and not w266;
w271 <= A(36) and not w268;
w272 <= not w270 and not w271;
w273 <= A(35) and not w272;
w274 <= not w269 and not w273;
w275 <= not A(33) and not w274;
w276 <= not A(34) and not w272;
w277 <= A(34) and not w274;
w278 <= not w276 and not w277;
w279 <= A(33) and not w278;
w280 <= not w275 and not w279;
w281 <= not A(31) and not w280;
w282 <= not A(32) and not w278;
w283 <= A(32) and not w280;
w284 <= not w282 and not w283;
w285 <= A(31) and not w284;
w286 <= not w281 and not w285;
w287 <= not A(29) and not w286;
w288 <= not A(30) and not w284;
w289 <= A(30) and not w286;
w290 <= not w288 and not w289;
w291 <= A(29) and not w290;
w292 <= not w287 and not w291;
w293 <= not A(27) and not w292;
w294 <= not A(28) and not w290;
w295 <= A(28) and not w292;
w296 <= not w294 and not w295;
w297 <= A(27) and not w296;
w298 <= not w293 and not w297;
w299 <= not A(25) and not w298;
w300 <= not A(26) and not w296;
w301 <= A(26) and not w298;
w302 <= not w300 and not w301;
w303 <= A(25) and not w302;
w304 <= not w299 and not w303;
w305 <= not A(23) and not w304;
w306 <= not A(24) and not w302;
w307 <= A(24) and not w304;
w308 <= not w306 and not w307;
w309 <= A(23) and not w308;
w310 <= not w305 and not w309;
w311 <= not A(21) and not w310;
w312 <= not A(22) and not w308;
w313 <= A(22) and not w310;
w314 <= not w312 and not w313;
w315 <= A(21) and not w314;
w316 <= not w311 and not w315;
w317 <= not A(19) and not w316;
w318 <= not A(20) and not w314;
w319 <= A(20) and not w316;
w320 <= not w318 and not w319;
w321 <= A(19) and not w320;
w322 <= not w317 and not w321;
w323 <= not A(17) and not w322;
w324 <= not A(18) and not w320;
w325 <= A(18) and not w322;
w326 <= not w324 and not w325;
w327 <= A(17) and not w326;
w328 <= not w323 and not w327;
w329 <= not A(15) and not w328;
w330 <= not A(16) and not w326;
w331 <= A(16) and not w328;
w332 <= not w330 and not w331;
w333 <= A(15) and not w332;
w334 <= not w329 and not w333;
w335 <= not A(13) and not w334;
w336 <= not A(14) and not w332;
w337 <= A(14) and not w334;
w338 <= not w336 and not w337;
w339 <= A(13) and not w338;
w340 <= not w335 and not w339;
w341 <= not A(11) and not w340;
w342 <= not A(12) and not w338;
w343 <= A(12) and not w340;
w344 <= not w342 and not w343;
w345 <= A(11) and not w344;
w346 <= not w341 and not w345;
w347 <= not A(9) and not w346;
w348 <= not A(10) and not w344;
w349 <= A(10) and not w346;
w350 <= not w348 and not w349;
w351 <= A(9) and not w350;
w352 <= not w347 and not w351;
w353 <= not A(7) and not w352;
w354 <= not A(8) and not w350;
w355 <= A(8) and not w352;
w356 <= not w354 and not w355;
w357 <= A(7) and not w356;
w358 <= not w353 and not w357;
w359 <= not A(5) and not w358;
w360 <= not A(6) and not w356;
w361 <= A(6) and not w358;
w362 <= not w360 and not w361;
w363 <= A(5) and not w362;
w364 <= not w359 and not w363;
w365 <= not A(3) and not w364;
w366 <= not A(4) and not w362;
w367 <= A(4) and not w364;
w368 <= not w366 and not w367;
w369 <= A(3) and not w368;
w370 <= not w365 and not w369;
w371 <= A(1) and not A(2);
w372 <= w370 and not w371;
w373 <= w368 and w371;
w374 <= not w372 and not w373;
w375 <= not A(126) and A(127);
w376 <= not A(126) and not w375;
w377 <= not A(124) and not A(125);
w378 <= not A(122) and not A(123);
w379 <= A(121) and w378;
w380 <= w377 and not w379;
w381 <= w376 and not w380;
w382 <= not A(120) and not w381;
w383 <= w377 and not w378;
w384 <= w376 and not w383;
w385 <= A(120) and not w384;
w386 <= not w382 and not w385;
w387 <= not A(118) and not A(119);
w388 <= w386 and not w387;
w389 <= w384 and w387;
w390 <= not w388 and not w389;
w391 <= not A(116) and not A(117);
w392 <= w390 and not w391;
w393 <= not w386 and w391;
w394 <= not w392 and not w393;
w395 <= not A(114) and not A(115);
w396 <= w394 and not w395;
w397 <= not w390 and w395;
w398 <= not w396 and not w397;
w399 <= not A(112) and not A(113);
w400 <= w398 and not w399;
w401 <= not w394 and w399;
w402 <= not w400 and not w401;
w403 <= not A(110) and not A(111);
w404 <= w402 and not w403;
w405 <= not w398 and w403;
w406 <= not w404 and not w405;
w407 <= not A(108) and not A(109);
w408 <= w406 and not w407;
w409 <= not w402 and w407;
w410 <= not w408 and not w409;
w411 <= not A(106) and not A(107);
w412 <= w410 and not w411;
w413 <= not w406 and w411;
w414 <= not w412 and not w413;
w415 <= not A(104) and not A(105);
w416 <= w414 and not w415;
w417 <= not w410 and w415;
w418 <= not w416 and not w417;
w419 <= not A(102) and not A(103);
w420 <= w418 and not w419;
w421 <= not w414 and w419;
w422 <= not w420 and not w421;
w423 <= not A(100) and not A(101);
w424 <= w422 and not w423;
w425 <= not w418 and w423;
w426 <= not w424 and not w425;
w427 <= not A(98) and not A(99);
w428 <= w426 and not w427;
w429 <= not w422 and w427;
w430 <= not w428 and not w429;
w431 <= not A(96) and not A(97);
w432 <= w430 and not w431;
w433 <= not w426 and w431;
w434 <= not w432 and not w433;
w435 <= not A(94) and not A(95);
w436 <= w434 and not w435;
w437 <= not w430 and w435;
w438 <= not w436 and not w437;
w439 <= not A(92) and not A(93);
w440 <= w438 and not w439;
w441 <= not w434 and w439;
w442 <= not w440 and not w441;
w443 <= not A(90) and not A(91);
w444 <= w442 and not w443;
w445 <= not w438 and w443;
w446 <= not w444 and not w445;
w447 <= not A(88) and not A(89);
w448 <= w446 and not w447;
w449 <= not w442 and w447;
w450 <= not w448 and not w449;
w451 <= not A(86) and not A(87);
w452 <= w450 and not w451;
w453 <= not w446 and w451;
w454 <= not w452 and not w453;
w455 <= not A(84) and not A(85);
w456 <= w454 and not w455;
w457 <= not w450 and w455;
w458 <= not w456 and not w457;
w459 <= not A(82) and not A(83);
w460 <= w458 and not w459;
w461 <= not w454 and w459;
w462 <= not w460 and not w461;
w463 <= not A(80) and not A(81);
w464 <= w462 and not w463;
w465 <= not w458 and w463;
w466 <= not w464 and not w465;
w467 <= not A(78) and not A(79);
w468 <= w466 and not w467;
w469 <= not w462 and w467;
w470 <= not w468 and not w469;
w471 <= not A(76) and not A(77);
w472 <= w470 and not w471;
w473 <= not w466 and w471;
w474 <= not w472 and not w473;
w475 <= not A(74) and not A(75);
w476 <= w474 and not w475;
w477 <= not w470 and w475;
w478 <= not w476 and not w477;
w479 <= not A(72) and not A(73);
w480 <= w478 and not w479;
w481 <= not w474 and w479;
w482 <= not w480 and not w481;
w483 <= not A(70) and not A(71);
w484 <= w482 and not w483;
w485 <= not w478 and w483;
w486 <= not w484 and not w485;
w487 <= not A(68) and not A(69);
w488 <= w486 and not w487;
w489 <= not w482 and w487;
w490 <= not w488 and not w489;
w491 <= not A(66) and not A(67);
w492 <= w490 and not w491;
w493 <= not w486 and w491;
w494 <= not w492 and not w493;
w495 <= not A(64) and not A(65);
w496 <= w494 and not w495;
w497 <= not w490 and w495;
w498 <= not w496 and not w497;
w499 <= not A(62) and not A(63);
w500 <= w498 and not w499;
w501 <= not w494 and w499;
w502 <= not w500 and not w501;
w503 <= not A(60) and not A(61);
w504 <= w502 and not w503;
w505 <= not w498 and w503;
w506 <= not w504 and not w505;
w507 <= not A(58) and not A(59);
w508 <= w506 and not w507;
w509 <= not w502 and w507;
w510 <= not w508 and not w509;
w511 <= not A(56) and not A(57);
w512 <= w510 and not w511;
w513 <= not w506 and w511;
w514 <= not w512 and not w513;
w515 <= not A(54) and not A(55);
w516 <= w514 and not w515;
w517 <= not w510 and w515;
w518 <= not w516 and not w517;
w519 <= not A(52) and not A(53);
w520 <= w518 and not w519;
w521 <= not w514 and w519;
w522 <= not w520 and not w521;
w523 <= not A(50) and not A(51);
w524 <= w522 and not w523;
w525 <= not w518 and w523;
w526 <= not w524 and not w525;
w527 <= not A(48) and not A(49);
w528 <= w526 and not w527;
w529 <= not w522 and w527;
w530 <= not w528 and not w529;
w531 <= not A(46) and not A(47);
w532 <= w530 and not w531;
w533 <= not w526 and w531;
w534 <= not w532 and not w533;
w535 <= not A(44) and not A(45);
w536 <= w534 and not w535;
w537 <= not w530 and w535;
w538 <= not w536 and not w537;
w539 <= not A(42) and not A(43);
w540 <= w538 and not w539;
w541 <= not w534 and w539;
w542 <= not w540 and not w541;
w543 <= not A(40) and not A(41);
w544 <= w542 and not w543;
w545 <= not w538 and w543;
w546 <= not w544 and not w545;
w547 <= not A(38) and not A(39);
w548 <= w546 and not w547;
w549 <= not w542 and w547;
w550 <= not w548 and not w549;
w551 <= not A(36) and not A(37);
w552 <= w550 and not w551;
w553 <= not w546 and w551;
w554 <= not w552 and not w553;
w555 <= not A(34) and not A(35);
w556 <= w554 and not w555;
w557 <= not w550 and w555;
w558 <= not w556 and not w557;
w559 <= not A(32) and not A(33);
w560 <= w558 and not w559;
w561 <= not w554 and w559;
w562 <= not w560 and not w561;
w563 <= not A(30) and not A(31);
w564 <= w562 and not w563;
w565 <= not w558 and w563;
w566 <= not w564 and not w565;
w567 <= not A(28) and not A(29);
w568 <= w566 and not w567;
w569 <= not w562 and w567;
w570 <= not w568 and not w569;
w571 <= not A(26) and not A(27);
w572 <= w570 and not w571;
w573 <= not w566 and w571;
w574 <= not w572 and not w573;
w575 <= not A(24) and not A(25);
w576 <= w574 and not w575;
w577 <= not w570 and w575;
w578 <= not w576 and not w577;
w579 <= not A(22) and not A(23);
w580 <= w578 and not w579;
w581 <= not w574 and w579;
w582 <= not w580 and not w581;
w583 <= not A(20) and not A(21);
w584 <= w582 and not w583;
w585 <= not w578 and w583;
w586 <= not w584 and not w585;
w587 <= not A(18) and not A(19);
w588 <= w586 and not w587;
w589 <= not w582 and w587;
w590 <= not w588 and not w589;
w591 <= not A(16) and not A(17);
w592 <= w590 and not w591;
w593 <= not w586 and w591;
w594 <= not w592 and not w593;
w595 <= not A(14) and not A(15);
w596 <= w594 and not w595;
w597 <= not w590 and w595;
w598 <= not w596 and not w597;
w599 <= not A(12) and not A(13);
w600 <= w598 and not w599;
w601 <= not w594 and w599;
w602 <= not w600 and not w601;
w603 <= not A(10) and not A(11);
w604 <= w602 and not w603;
w605 <= not w598 and w603;
w606 <= not w604 and not w605;
w607 <= not A(8) and not A(9);
w608 <= w606 and not w607;
w609 <= not w602 and w607;
w610 <= not w608 and not w609;
w611 <= not A(6) and not A(7);
w612 <= w610 and not w611;
w613 <= not w606 and w611;
w614 <= not w612 and not w613;
w615 <= not A(4) and not A(5);
w616 <= w614 and not w615;
w617 <= not w610 and w615;
w618 <= not w616 and not w617;
w619 <= not A(2) and not A(3);
w620 <= w618 and not w619;
w621 <= not w614 and w619;
w622 <= not w620 and not w621;
w623 <= w376 and w377;
w624 <= not A(120) and not A(121);
w625 <= w378 and w624;
w626 <= not A(117) and w387;
w627 <= not A(116) and w626;
w628 <= w625 and not w627;
w629 <= w623 and not w628;
w630 <= not A(113) and not A(114);
w631 <= not A(112) and w630;
w632 <= w629 and not w631;
w633 <= A(115) and w627;
w634 <= w625 and not w633;
w635 <= w623 and not w634;
w636 <= w631 and w635;
w637 <= not w632 and not w636;
w638 <= not A(109) and w403;
w639 <= not A(108) and w638;
w640 <= w637 and not w639;
w641 <= not w629 and w639;
w642 <= not w640 and not w641;
w643 <= not A(105) and w411;
w644 <= not A(104) and w643;
w645 <= w642 and not w644;
w646 <= not w637 and w644;
w647 <= not w645 and not w646;
w648 <= not A(101) and w419;
w649 <= not A(100) and w648;
w650 <= w647 and not w649;
w651 <= not w642 and w649;
w652 <= not w650 and not w651;
w653 <= not A(97) and w427;
w654 <= not A(96) and w653;
w655 <= w652 and not w654;
w656 <= not w647 and w654;
w657 <= not w655 and not w656;
w658 <= not A(93) and w435;
w659 <= not A(92) and w658;
w660 <= w657 and not w659;
w661 <= not w652 and w659;
w662 <= not w660 and not w661;
w663 <= not A(89) and w443;
w664 <= not A(88) and w663;
w665 <= w662 and not w664;
w666 <= not w657 and w664;
w667 <= not w665 and not w666;
w668 <= not A(85) and w451;
w669 <= not A(84) and w668;
w670 <= w667 and not w669;
w671 <= not w662 and w669;
w672 <= not w670 and not w671;
w673 <= not A(81) and w459;
w674 <= not A(80) and w673;
w675 <= w672 and not w674;
w676 <= not w667 and w674;
w677 <= not w675 and not w676;
w678 <= not A(77) and w467;
w679 <= not A(76) and w678;
w680 <= w677 and not w679;
w681 <= not w672 and w679;
w682 <= not w680 and not w681;
w683 <= not A(73) and w475;
w684 <= not A(72) and w683;
w685 <= w682 and not w684;
w686 <= not w677 and w684;
w687 <= not w685 and not w686;
w688 <= not A(69) and w483;
w689 <= not A(68) and w688;
w690 <= w687 and not w689;
w691 <= not w682 and w689;
w692 <= not w690 and not w691;
w693 <= not A(65) and w491;
w694 <= not A(64) and w693;
w695 <= w692 and not w694;
w696 <= not w687 and w694;
w697 <= not w695 and not w696;
w698 <= not A(61) and w499;
w699 <= not A(60) and w698;
w700 <= w697 and not w699;
w701 <= not w692 and w699;
w702 <= not w700 and not w701;
w703 <= not A(57) and w507;
w704 <= not A(56) and w703;
w705 <= w702 and not w704;
w706 <= not w697 and w704;
w707 <= not w705 and not w706;
w708 <= not A(53) and w515;
w709 <= not A(52) and w708;
w710 <= w707 and not w709;
w711 <= not w702 and w709;
w712 <= not w710 and not w711;
w713 <= not A(49) and w523;
w714 <= not A(48) and w713;
w715 <= w712 and not w714;
w716 <= not w707 and w714;
w717 <= not w715 and not w716;
w718 <= not A(45) and w531;
w719 <= not A(44) and w718;
w720 <= w717 and not w719;
w721 <= not w712 and w719;
w722 <= not w720 and not w721;
w723 <= not A(41) and w539;
w724 <= not A(40) and w723;
w725 <= w722 and not w724;
w726 <= not w717 and w724;
w727 <= not w725 and not w726;
w728 <= not A(37) and w547;
w729 <= not A(36) and w728;
w730 <= w727 and not w729;
w731 <= not w722 and w729;
w732 <= not w730 and not w731;
w733 <= not A(33) and w555;
w734 <= not A(32) and w733;
w735 <= w732 and not w734;
w736 <= not w727 and w734;
w737 <= not w735 and not w736;
w738 <= not A(29) and w563;
w739 <= not A(28) and w738;
w740 <= w737 and not w739;
w741 <= not w732 and w739;
w742 <= not w740 and not w741;
w743 <= not A(25) and w571;
w744 <= not A(24) and w743;
w745 <= w742 and not w744;
w746 <= not w737 and w744;
w747 <= not w745 and not w746;
w748 <= not A(21) and w579;
w749 <= not A(20) and w748;
w750 <= w747 and not w749;
w751 <= not w742 and w749;
w752 <= not w750 and not w751;
w753 <= not A(17) and w587;
w754 <= not A(16) and w753;
w755 <= w752 and not w754;
w756 <= not w747 and w754;
w757 <= not w755 and not w756;
w758 <= not A(13) and w595;
w759 <= not A(12) and w758;
w760 <= w757 and not w759;
w761 <= not w752 and w759;
w762 <= not w760 and not w761;
w763 <= not A(9) and w603;
w764 <= not A(8) and w763;
w765 <= w762 and not w764;
w766 <= not w757 and w764;
w767 <= not w765 and not w766;
w768 <= not A(5) and w611;
w769 <= not A(4) and w768;
w770 <= w767 and not w769;
w771 <= not w762 and w769;
w772 <= not w770 and not w771;
w773 <= w623 and w625;
w774 <= not A(113) and w395;
w775 <= not A(112) and w627;
w776 <= w774 and w775;
w777 <= not A(107) and w639;
w778 <= not A(106) and w777;
w779 <= not A(105) and w778;
w780 <= not A(104) and w779;
w781 <= w776 and not w780;
w782 <= w773 and not w781;
w783 <= not A(101) and not A(102);
w784 <= not A(100) and w783;
w785 <= not A(99) and w784;
w786 <= not A(98) and w785;
w787 <= not A(97) and w786;
w788 <= not A(96) and w787;
w789 <= w782 and not w788;
w790 <= A(103) and w780;
w791 <= w776 and not w790;
w792 <= w773 and not w791;
w793 <= w788 and w792;
w794 <= not w789 and not w793;
w795 <= not A(91) and w659;
w796 <= not A(90) and w795;
w797 <= not A(89) and w796;
w798 <= not A(88) and w797;
w799 <= w794 and not w798;
w800 <= not w782 and w798;
w801 <= not w799 and not w800;
w802 <= not A(83) and w669;
w803 <= not A(82) and w802;
w804 <= not A(81) and w803;
w805 <= not A(80) and w804;
w806 <= w801 and not w805;
w807 <= not w794 and w805;
w808 <= not w806 and not w807;
w809 <= not A(75) and w679;
w810 <= not A(74) and w809;
w811 <= not A(73) and w810;
w812 <= not A(72) and w811;
w813 <= w808 and not w812;
w814 <= not w801 and w812;
w815 <= not w813 and not w814;
w816 <= not A(67) and w689;
w817 <= not A(66) and w816;
w818 <= not A(65) and w817;
w819 <= not A(64) and w818;
w820 <= w815 and not w819;
w821 <= not w808 and w819;
w822 <= not w820 and not w821;
w823 <= not A(59) and w699;
w824 <= not A(58) and w823;
w825 <= not A(57) and w824;
w826 <= not A(56) and w825;
w827 <= w822 and not w826;
w828 <= not w815 and w826;
w829 <= not w827 and not w828;
w830 <= not A(51) and w709;
w831 <= not A(50) and w830;
w832 <= not A(49) and w831;
w833 <= not A(48) and w832;
w834 <= w829 and not w833;
w835 <= not w822 and w833;
w836 <= not w834 and not w835;
w837 <= not A(43) and w719;
w838 <= not A(42) and w837;
w839 <= not A(41) and w838;
w840 <= not A(40) and w839;
w841 <= w836 and not w840;
w842 <= not w829 and w840;
w843 <= not w841 and not w842;
w844 <= not A(35) and w729;
w845 <= not A(34) and w844;
w846 <= not A(33) and w845;
w847 <= not A(32) and w846;
w848 <= w843 and not w847;
w849 <= not w836 and w847;
w850 <= not w848 and not w849;
w851 <= not A(27) and w739;
w852 <= not A(26) and w851;
w853 <= not A(25) and w852;
w854 <= not A(24) and w853;
w855 <= w850 and not w854;
w856 <= not w843 and w854;
w857 <= not w855 and not w856;
w858 <= not A(19) and w749;
w859 <= not A(18) and w858;
w860 <= not A(17) and w859;
w861 <= not A(16) and w860;
w862 <= w857 and not w861;
w863 <= not w850 and w861;
w864 <= not w862 and not w863;
w865 <= not A(11) and w759;
w866 <= not A(10) and w865;
w867 <= not A(9) and w866;
w868 <= not A(8) and w867;
w869 <= w864 and not w868;
w870 <= not w857 and w868;
w871 <= not w869 and not w870;
w872 <= w773 and w776;
w873 <= not A(99) and w649;
w874 <= not A(98) and w780;
w875 <= not A(97) and w874;
w876 <= not A(96) and w875;
w877 <= w873 and w876;
w878 <= not A(87) and w798;
w879 <= not A(86) and w878;
w880 <= not A(85) and w879;
w881 <= not A(84) and w880;
w882 <= not A(83) and w881;
w883 <= not A(82) and w882;
w884 <= not A(81) and w883;
w885 <= not A(80) and w884;
w886 <= w877 and not w885;
w887 <= w872 and not w886;
w888 <= not A(77) and not A(78);
w889 <= not A(76) and w888;
w890 <= not A(75) and w889;
w891 <= not A(74) and w890;
w892 <= not A(73) and w891;
w893 <= not A(72) and w892;
w894 <= not A(71) and w893;
w895 <= not A(70) and w894;
w896 <= not A(69) and w895;
w897 <= not A(68) and w896;
w898 <= not A(67) and w897;
w899 <= not A(66) and w898;
w900 <= not A(65) and w899;
w901 <= not A(64) and w900;
w902 <= w887 and not w901;
w903 <= A(79) and w885;
w904 <= w877 and not w903;
w905 <= w872 and not w904;
w906 <= w901 and w905;
w907 <= not w902 and not w906;
w908 <= not A(55) and w826;
w909 <= not A(54) and w908;
w910 <= not A(53) and w909;
w911 <= not A(52) and w910;
w912 <= not A(51) and w911;
w913 <= not A(50) and w912;
w914 <= not A(49) and w913;
w915 <= not A(48) and w914;
w916 <= w907 and not w915;
w917 <= not w887 and w915;
w918 <= not w916 and not w917;
w919 <= not A(39) and w840;
w920 <= not A(38) and w919;
w921 <= not A(37) and w920;
w922 <= not A(36) and w921;
w923 <= not A(35) and w922;
w924 <= not A(34) and w923;
w925 <= not A(33) and w924;
w926 <= not A(32) and w925;
w927 <= w918 and not w926;
w928 <= not w907 and w926;
w929 <= not w927 and not w928;
w930 <= not A(23) and w854;
w931 <= not A(22) and w930;
w932 <= not A(21) and w931;
w933 <= not A(20) and w932;
w934 <= not A(19) and w933;
w935 <= not A(18) and w934;
w936 <= not A(17) and w935;
w937 <= not A(16) and w936;
w938 <= w929 and not w937;
w939 <= not w918 and w937;
w940 <= not w938 and not w939;
w941 <= w872 and w877;
w942 <= not A(71) and w812;
w943 <= not A(70) and w885;
w944 <= not A(69) and w943;
w945 <= not A(68) and w944;
w946 <= not A(67) and w945;
w947 <= not A(66) and w946;
w948 <= not A(65) and w947;
w949 <= not A(64) and w948;
w950 <= w942 and w949;
w951 <= not A(47) and w915;
w952 <= not A(46) and w951;
w953 <= not A(45) and w952;
w954 <= not A(44) and w953;
w955 <= not A(43) and w954;
w956 <= not A(42) and w955;
w957 <= not A(41) and w956;
w958 <= not A(40) and w957;
w959 <= not A(39) and w958;
w960 <= not A(38) and w959;
w961 <= not A(37) and w960;
w962 <= not A(36) and w961;
w963 <= not A(35) and w962;
w964 <= not A(34) and w963;
w965 <= not A(33) and w964;
w966 <= not A(32) and w965;
w967 <= w950 and not w966;
w968 <= w941 and not w967;
w969 <= w941 and w950;
w970 <= not A(0) and w969;
w971 <= w868 and w970;
w972 <= not A(3) and w971;
w973 <= not A(2) and w972;
w974 <= w937 and w966;
w975 <= w769 and w974;
w976 <= not A(1) and w975;
w977 <= w973 and w976;
one <= '1';
P(0) <= w374;-- level 250
P(1) <= w622;-- level 124
P(2) <= not w772;-- level 62
P(3) <= not w871;-- level 34
P(4) <= not w940;-- level 26
P(5) <= not w968;-- level 33
P(6) <= not w969;-- level 24
F <= not w977;-- level 35
end Behavioral;