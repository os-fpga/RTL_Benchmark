module BUFG (
   input wire I,
   output wire O
   );

   assign O = I;
   
endmodule