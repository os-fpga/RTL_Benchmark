`ifdef SAMPLE_AE350_SMU_CONFIG_VH
`else
`define SAMPLE_AE350_SMU_CONFIG_VH


`endif // SAMPLE_AE350_SMU_CONFIG_VH

