// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: rca_monitor.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Tue Mar 19 21:50:30 2019
//=============================================================================
// Description: Monitor for rca
//=============================================================================

`ifndef RCA_MONITOR_SV
`define RCA_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file rca.tpl

class rca_monitor extends uvm_monitor;

  `uvm_component_utils(rca_monitor)

  virtual rca_if vif;

  uvm_analysis_port #(trans) analysis_port;

  trans m_trans;

  extern function new(string name, uvm_component parent);

  // Methods build_phase, run_phase, and do_mon generated by setting monitor_inc in file rca.tpl
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file rca.tpl

endclass : rca_monitor 


function rca_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


function void rca_monitor::build_phase(uvm_phase phase);
endfunction : build_phase


task rca_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = trans::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/rca_monitor_inc.sv
task rca_monitor::do_mon;
  forever @(posedge vif.clk)
    begin
	  m_trans.input1 = vif.a;
	  m_trans.input2 = vif.b;
	  m_trans.carryinput = vif.ci;
	  m_trans.carryoutput = vif.co;
	  m_trans.sum = vif.s;
	  analysis_port.write(m_trans);
	  `uvm_info(get_type_name(),$sformatf("a(%0d) + b(%0d) + ci(%0d) = co(%0d) and s(%0d)", vif.a, vif.b, vif.ci, vif.co, vif.s), UVM_MEDIUM);
    end
endtask// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file rca.tpl

`endif // RCA_MONITOR_SV

