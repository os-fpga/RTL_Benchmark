`ifndef _REG_MAP_VH_
`define _REG_MAP_VH_
localparam REG_USTATUS  = 12'h000;
localparam REG_NONE     = REG_USTATUS;
localparam REG_SSTATUS  = 12'h100;
localparam REG_SATP     = 12'h180;

localparam REG_MSTATUS  = 12'h300;
localparam REG_MISA     = 12'h301;
localparam REG_MSCRATCH = 12'h340;

localparam REG_MMSC_CFG = 12'hfc2;

localparam REG_DCSR     = 12'h7b0;
localparam REG_DPC      = 12'h7b1;
localparam REG_DSCRATCH0= 12'h7b2;
localparam REG_DSCRATCH1= 12'h7b3;
localparam REG_TSELECT  = 12'h7a0;
localparam REG_TDATA1   = 12'h7a1;
localparam REG_TDATA2   = 12'h7a2;
localparam REG_TDATA3   = 12'h7a3;
localparam REG_TINFO    = 12'h7a4;
localparam REG_TCONTROL = 12'h7a5;

localparam REG_VSTART   = 12'h008;
localparam REG_VXSAT    = 12'h009;
localparam REG_VXRM     = 12'h00A;
localparam REG_VCSR     = 12'h00F;
localparam REG_VL       = 12'hC20;
localparam REG_VTYPE    = 12'hC21;
localparam REG_VLENB    = 12'hC22;

localparam REG_CYCLE	= 12'hb00;
localparam REG_CYCLEH	= 12'hb80;
localparam REG_INSTRET	= 12'hb02;
localparam REG_INSTRETH	= 12'hb82;
localparam REG_MCOUNTERMASK_M = 12'h7d1;
localparam REG_MCOUNTERMASK_S = 12'h7d2;
localparam REG_MCOUNTERMASK_U = 12'h7d3;

localparam GPR_X0	= 5'd0;
localparam GPR_X1	= 5'd1;
localparam GPR_X2	= 5'd2;
localparam GPR_X3	= 5'd3;
localparam GPR_X4	= 5'd4;
localparam GPR_X5	= 5'd5;
localparam GPR_X6	= 5'd6;
localparam GPR_X7	= 5'd7;
localparam GPR_X8	= 5'd8;
localparam GPR_X9	= 5'd9;
localparam GPR_X10	= 5'd10;
localparam GPR_X11	= 5'd11;
localparam GPR_X12	= 5'd12;
localparam GPR_X13	= 5'd13;
localparam GPR_X14	= 5'd14;
localparam GPR_X15	= 5'd15;
localparam GPR_X16	= 5'd16;
localparam GPR_X17	= 5'd17;
localparam GPR_X18	= 5'd18;
localparam GPR_X19	= 5'd19;
localparam GPR_X20	= 5'd20;
localparam GPR_X21	= 5'd21;
localparam GPR_X22	= 5'd22;
localparam GPR_X23	= 5'd23;
localparam GPR_X24	= 5'd24;
localparam GPR_X25	= 5'd25;
localparam GPR_X26	= 5'd26;
localparam GPR_X27	= 5'd27;
localparam GPR_X28	= 5'd28;
localparam GPR_X29	= 5'd29;
localparam GPR_X30	= 5'd30;
localparam GPR_X31	= 5'd31;

localparam FPR_F0	= 5'd0;
localparam FPR_F1	= 5'd1;
localparam FPR_F2	= 5'd2;
localparam FPR_F3	= 5'd3;
localparam FPR_F4	= 5'd4;
localparam FPR_F5	= 5'd5;
localparam FPR_F6	= 5'd6;
localparam FPR_F7	= 5'd7;
localparam FPR_F8	= 5'd8;
localparam FPR_F9	= 5'd9;
localparam FPR_F10	= 5'd10;
localparam FPR_F11	= 5'd11;
localparam FPR_F12	= 5'd12;
localparam FPR_F13	= 5'd13;
localparam FPR_F14	= 5'd14;
localparam FPR_F15	= 5'd15;
localparam FPR_F16	= 5'd16;
localparam FPR_F17	= 5'd17;
localparam FPR_F18	= 5'd18;
localparam FPR_F19	= 5'd19;
localparam FPR_F20	= 5'd20;
localparam FPR_F21	= 5'd21;
localparam FPR_F22	= 5'd22;
localparam FPR_F23	= 5'd23;
localparam FPR_F24	= 5'd24;
localparam FPR_F25	= 5'd25;
localparam FPR_F26	= 5'd26;
localparam FPR_F27	= 5'd27;
localparam FPR_F28	= 5'd28;
localparam FPR_F29	= 5'd29;
localparam FPR_F30	= 5'd30;
localparam FPR_F31	= 5'd31;

localparam GPR_ZERO	= 5'd0;
localparam GPR_RA	= 5'd1;
localparam GPR_SP	= 5'd2;
localparam GPR_GP	= 5'd3;
localparam GPR_TP	= 5'd4;
localparam GPR_T0	= 5'd5;
localparam GPR_T1	= 5'd6;
localparam GPR_T2	= 5'd7;
localparam GPR_S0	= 5'd8;
localparam GPR_S1	= 5'd9;
localparam GPR_A0	= 5'd10;
localparam GPR_A1	= 5'd11;
localparam GPR_A2	= 5'd12;
localparam GPR_A3	= 5'd13;
localparam GPR_A4	= 5'd14;
localparam GPR_A5	= 5'd15;
localparam GPR_A6	= 5'd16;
localparam GPR_A7	= 5'd17;
localparam GPR_S2	= 5'd18;
localparam GPR_S3	= 5'd19;
localparam GPR_S4	= 5'd20;
localparam GPR_S5	= 5'd21;
localparam GPR_S6	= 5'd22;
localparam GPR_S7	= 5'd23;
localparam GPR_S8	= 5'd24;
localparam GPR_S9	= 5'd25;
localparam GPR_S10	= 5'd26;
localparam GPR_S11	= 5'd27;
localparam GPR_T3	= 5'd28;
localparam GPR_T4	= 5'd29;
localparam GPR_T5	= 5'd30;
localparam GPR_T6	= 5'd31;

localparam FPR_FT0	= 5'd0;
localparam FPR_FT1	= 5'd1;
localparam FPR_FT2	= 5'd2;
localparam FPR_FT3	= 5'd3;
localparam FPR_FT4	= 5'd4;
localparam FPR_FT5	= 5'd5;
localparam FPR_FT6	= 5'd6;
localparam FPR_FT7	= 5'd7;
localparam FPR_FS0	= 5'd8;
localparam FPR_FS1	= 5'd9;
localparam FPR_FA0	= 5'd10;
localparam FPR_FA1	= 5'd11;
localparam FPR_FA2	= 5'd12;
localparam FPR_FA3	= 5'd13;
localparam FPR_FA4	= 5'd14;
localparam FPR_FA5	= 5'd15;
localparam FPR_FA6	= 5'd16;
localparam FPR_FA7	= 5'd17;
localparam FPR_FS2	= 5'd18;
localparam FPR_FS3	= 5'd19;
localparam FPR_FS4	= 5'd20;
localparam FPR_FS5	= 5'd21;
localparam FPR_FS6	= 5'd22;
localparam FPR_FS7	= 5'd23;
localparam FPR_FS8	= 5'd24;
localparam FPR_FS9	= 5'd25;
localparam FPR_FS10	= 5'd26;
localparam FPR_FS11	= 5'd27;
localparam FPR_FT8	= 5'd28;
localparam FPR_FT9	= 5'd29;
localparam FPR_FT10	= 5'd30;
localparam FPR_FT11	= 5'd31;
`endif

