----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Istvan Nagy, buenos@freemail.hu
-- 
-- Create Date:    15:58:13 05/30/2010 
-- Design Name: 
-- Module Name:    s6bfip_memory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
-- This memory controller was generated for the Hynix H5PS5162FFR-S6C memory
--  chip, but based on the Elpida EDE5116AJBG chip parameters in the MIG-tool.
--  The memory data rate was specified as 500Mt/s, using 250MHz reference clock.
--  The refclk is expected to be as a single ended on-board signal, so here
--  we have to generate is with a PLL and route it out to the PCB then back to 
--  the MCB. If it is possible, then try to use internal routing using bufpll-mcb.
--
-- Refclk: from PLL. The PLL is normally driven by an external pin.
--  That pin is connected to an OBUFDS, driven by BUFPLL. we can conenct the input of
--  the PLL to a BUFG, running from one of the on-chip clocks.
-- The entity memc3_infrastructure contains the PLL.
--   It has: 
--     sys_clk -> sys_clk_ibufg -> PLL[(CLKIN1)=>(div=1)(CLKOUT0)] -> clk_2x_0 -> BUFPLL_MCB
--   It also contains a IBUFG/IBUFGDS for the sys_clk, that has to be removed, and this has
--   to be added instead: sys_clk_ibufg <= sys_clk;
--   Connect c3_sys_clk to the on-chip 25MHz clock (x25m_clk) in this file.
--   The PLL multiplier has to be changed, to multiply the 25MHz to 500MHz, by 20.
--    CLKFBOUT_MULT      => 20,
--
-- MCB user guide (ug388) CLOCKING notes:
-- ==============================
--The MCB requires three basic types of clocks:
-- - MCB system clocks determine the operating frequency of the memory controller and
--physical interface to the external memory device.
-- - Calibration clock determines the operating frequency of the calibration logic.
-- - User clocks determine the operating frequency of the User Interface ports. These
--clocks can be completely asynchronous to the system and calibration clocks. The
--Command and Data Path FIFOs handle the necessary clock domain transfer from the
--User Interface to the internal controller logic.
--
--It must be driven by the I/O clock network (BUFPLL_MCB). The I/O clock network is
--designed for significantly higher frequencies than the global clock network, allowing
--memory interfaces to operate at up to 800 Mb/s.
--
--To create the desired system clock frequency on the I/O clock network, an external clock
--source drives one of the PLLs in the center column of the device. The external clock
--frequency is not critical as long as the PLL can synthesize the desired MCB system clocks
--from it.
--The PLL generates two system clock outputs, sysclk_2x and sysclk_2x_180, that are twice
--the frequency of the desired memory clock (for example, for a 800 Mb/s DDR2 interface
--with a memory clock equal to 400 MHz, the system clocks are set to 800 MHz) and 180
--degrees out of phase from each other. Only two clock lines are available on each side of the
--device to drive the I/O clock network from the PLLs. The pair of system clocks uses these
--two clock lines to connect to the MCBs on the left or right side of the device. Thus for
--devices with four MCBs, the two MCBs on the same side of the device must share the same
--system clock pair and therefore must run at the same data rate, although the memory
--standard implemented can be different. DCMs do not have access to the I/O clock network
--and cannot, therefore, be used to drive MCBs.
--When the pair of system clocks reaches the I/O clock network, they are rebuffered by a
--BUFPLL_MCB driver. This driver also creates clock enable strobes required by the MCB:
--pll_ce_0 and pll_ce_90.
--
--The calibration related clock, mcb_drp_clk, must be generated by the PLL and must be
--phase-synchronized (i.e., in phase) with the sysclk_2x domain.The calibration clock rate is
--limited by normal static timing analysis, with a typical achievable frequency of 100 MHz.
--In general, a calibration clock frequency of at least 50 MHz should be used to allow the
--MCB to complete calibration operations in a reasonable period of time.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;


entity s6bfip_memory is
    Port (--FPGA_PINS (EXTERNAL):
			  mcb3_dram_dq        : inout  std_logic_vector(15 downto 0);
			  mcb3_dram_a         : out std_logic_vector(12 downto 0);
			  mcb3_dram_ba        : out std_logic_vector(1 downto 0);
			  mcb3_dram_ras_n     : out std_logic;
			  mcb3_dram_cas_n     : out std_logic;
			  mcb3_dram_we_n      : out std_logic;
			  mcb3_dram_odt       : out std_logic;
			  mcb3_dram_cke       : out std_logic;
			  mcb3_dram_dm        : out std_logic;
			  mcb3_dram_udqs      : inout  std_logic;
			  mcb3_dram_udqs_n    : inout  std_logic;
			  mcb3_rzq            : inout  std_logic;
			  mcb3_zio            : inout  std_logic;
			  mcb3_dram_udm       : out std_logic;
			  mcb3_dram_dqs       : inout  std_logic;
			  mcb3_dram_dqs_n     : inout  std_logic;
			  mcb3_dram_ck        : out std_logic;
			  mcb3_dram_ck_n      : out std_logic;	
			  --ONCHIP PORTS:
			  --channel-0
			  channel0_wb_data_i : in std_logic_vector(31 downto 0); 
			  channel0_wb_data_o : out std_logic_vector(31 downto 0);
			  channel0_wb_addr_i : in std_logic_vector(25 downto 0);
			  channel0_wb_cyc_i : in std_logic;
			  channel0_wb_stb_i : in std_logic;
			  channel0_wb_wr_i : in std_logic;
			  channel0_wb_ack_o : out std_logic;
			  channel0_wb_clk_i : in std_logic; 	
			  channel0_wb_sel_i : in std_logic_vector(3 downto 0);
			  --channel-1
			  channel1_wb_data_i : in std_logic_vector(31 downto 0); 
			  channel1_wb_data_o : out std_logic_vector(31 downto 0);
			  channel1_wb_addr_i : in std_logic_vector(25 downto 0);
			  channel1_wb_cyc_i : in std_logic;
			  channel1_wb_stb_i : in std_logic;
			  channel1_wb_wr_i : in std_logic;
			  channel1_wb_ack_o : out std_logic;
			  channel1_wb_clk_i : in std_logic; 
			  channel1_wb_sel_i : in std_logic_vector(3 downto 0);
			  --channel-2
			  channel2_wb_data_i : in std_logic_vector(31 downto 0); 
			  channel2_wb_data_o : out std_logic_vector(31 downto 0);
			  channel2_wb_addr_i : in std_logic_vector(25 downto 0);
			  channel2_wb_cyc_i : in std_logic;
			  channel2_wb_stb_i : in std_logic;
			  channel2_wb_wr_i : in std_logic;
			  channel2_wb_ack_o : out std_logic;
			  channel2_wb_clk_i : in std_logic; 
			  channel2_wb_sel_i : in std_logic_vector(3 downto 0);
			  --channel-3
			  channel3_wb_data_i : in std_logic_vector(31 downto 0); 
			  channel3_wb_data_o : out std_logic_vector(31 downto 0);
			  channel3_wb_addr_i : in std_logic_vector(25 downto 0);
			  channel3_wb_cyc_i : in std_logic;
			  channel3_wb_stb_i : in std_logic;
			  channel3_wb_wr_i : in std_logic;
			  channel3_wb_ack_o : out std_logic;
			  channel3_wb_clk_i : in std_logic; 
			  channel3_wb_sel_i : in std_logic_vector(3 downto 0);
			  --System signals:
			  x25m_clk : in std_logic; 
			  reset : in std_logic 
			 );
end s6bfip_memory;

architecture Behavioral of s6bfip_memory is

   -- Internal Signals ------------------------------------------------------------
	--SIGNAL dummy : std_logic_vector(15 downto 0);	--write data bus
	SIGNAL c3_sys_clk :  std_logic;
	SIGNAL c3_sys_rst_n :  std_logic;
	SIGNAL c3_p0_cmd_clk :  std_logic;
	SIGNAL c3_p0_cmd_en :  std_logic;
	SIGNAL c3_p0_cmd_instr :  std_logic_vector(2 downto 0);
	SIGNAL c3_p0_cmd_bl :  std_logic_vector(5 downto 0);
	SIGNAL c3_p0_cmd_byte_addr :  std_logic_vector(29 downto 0);
	SIGNAL c3_p0_wr_clk :  std_logic;
	SIGNAL c3_p0_wr_en :  std_logic;
	SIGNAL c3_p0_wr_mask :  std_logic_vector(3 downto 0);
	SIGNAL c3_p0_wr_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p0_rd_clk :  std_logic;
	SIGNAL c3_p0_rd_en :  std_logic;
	SIGNAL c3_p1_cmd_clk :  std_logic;
	SIGNAL c3_p1_cmd_en :  std_logic;
	SIGNAL c3_p1_cmd_instr :  std_logic_vector(2 downto 0);
	SIGNAL c3_p1_cmd_bl :  std_logic_vector(5 downto 0);
	SIGNAL c3_p1_cmd_byte_addr :  std_logic_vector(29 downto 0);
	SIGNAL c3_p1_wr_clk :  std_logic;
	SIGNAL c3_p1_wr_en :  std_logic;
	SIGNAL c3_p1_wr_mask :  std_logic_vector(3 downto 0);
	SIGNAL c3_p1_wr_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p1_rd_clk :  std_logic;
	SIGNAL c3_p1_rd_en :  std_logic;
	SIGNAL c3_p2_cmd_clk :  std_logic;
	SIGNAL c3_p2_cmd_en :  std_logic;
	SIGNAL c3_p2_cmd_instr :  std_logic_vector(2 downto 0);
	SIGNAL c3_p2_cmd_bl :  std_logic_vector(5 downto 0);
	SIGNAL c3_p2_cmd_byte_addr :  std_logic_vector(29 downto 0);
	SIGNAL c3_p2_wr_clk :  std_logic;
	SIGNAL c3_p2_wr_en :  std_logic;
	SIGNAL c3_p2_wr_mask :  std_logic_vector(3 downto 0);
	SIGNAL c3_p2_wr_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p2_rd_clk :  std_logic;
	SIGNAL c3_p2_rd_en :  std_logic;
	SIGNAL c3_p3_cmd_clk :  std_logic;
	SIGNAL c3_p3_cmd_en :  std_logic;
	SIGNAL c3_p3_cmd_instr :  std_logic_vector(2 downto 0);
	SIGNAL c3_p3_cmd_bl :  std_logic_vector(5 downto 0);
	SIGNAL c3_p3_cmd_byte_addr :  std_logic_vector(29 downto 0);
	SIGNAL c3_p3_wr_clk :  std_logic;
	SIGNAL c3_p3_wr_en :  std_logic;
	SIGNAL c3_p3_wr_mask :  std_logic_vector(3 downto 0);
	SIGNAL c3_p3_wr_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p3_rd_clk :  std_logic;
	SIGNAL c3_p3_rd_en :  std_logic;    
	SIGNAL c3_calib_done :  std_logic;
	SIGNAL c3_clk0 :  std_logic;
	SIGNAL c3_rst0 :  std_logic;
	SIGNAL c3_p0_cmd_empty :  std_logic;
	SIGNAL c3_p0_cmd_full :  std_logic;
	SIGNAL c3_p0_wr_full :  std_logic;
	SIGNAL c3_p0_wr_empty :  std_logic;
	SIGNAL c3_p0_wr_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p0_wr_underrun :  std_logic;
	SIGNAL c3_p0_wr_error :  std_logic;
	SIGNAL c3_p0_rd_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p0_rd_full :  std_logic;
	SIGNAL c3_p0_rd_empty :  std_logic;
	SIGNAL c3_p0_rd_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p0_rd_overflow :  std_logic;
	SIGNAL c3_p0_rd_error :  std_logic;
	SIGNAL c3_p1_cmd_empty :  std_logic;
	SIGNAL c3_p1_cmd_full :  std_logic;
	SIGNAL c3_p1_wr_full :  std_logic;
	SIGNAL c3_p1_wr_empty :  std_logic;
	SIGNAL c3_p1_wr_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p1_wr_underrun :  std_logic;
	SIGNAL c3_p1_wr_error :  std_logic;
	SIGNAL c3_p1_rd_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p1_rd_full :  std_logic;
	SIGNAL c3_p1_rd_empty :  std_logic;
	SIGNAL c3_p1_rd_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p1_rd_overflow :  std_logic;
	SIGNAL c3_p1_rd_error :  std_logic;
	SIGNAL c3_p2_cmd_empty :  std_logic;
	SIGNAL c3_p2_cmd_full :  std_logic;
	SIGNAL c3_p2_wr_full :  std_logic;
	SIGNAL c3_p2_wr_empty :  std_logic;
	SIGNAL c3_p2_wr_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p2_wr_underrun :  std_logic;
	SIGNAL c3_p2_wr_error :  std_logic;
	SIGNAL c3_p2_rd_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p2_rd_full :  std_logic;
	SIGNAL c3_p2_rd_empty :  std_logic;
	SIGNAL c3_p2_rd_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p2_rd_overflow :  std_logic;
	SIGNAL c3_p2_rd_error :  std_logic;
	SIGNAL c3_p3_cmd_empty :  std_logic;
	SIGNAL c3_p3_cmd_full :  std_logic;
	SIGNAL c3_p3_wr_full :  std_logic;
	SIGNAL c3_p3_wr_empty :  std_logic;
	SIGNAL c3_p3_wr_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p3_wr_underrun :  std_logic;
	SIGNAL c3_p3_wr_error :  std_logic;
	SIGNAL c3_p3_rd_data :  std_logic_vector(31 downto 0);
	SIGNAL c3_p3_rd_full :  std_logic;
	SIGNAL c3_p3_rd_empty :  std_logic;
	SIGNAL c3_p3_rd_count :  std_logic_vector(6 downto 0);
	SIGNAL c3_p3_rd_overflow :  std_logic;
	SIGNAL c3_p3_rd_error :  std_logic;
	
	SIGNAL channel0_wb_state :  std_logic_vector(3 downto 0);
	SIGNAL channel1_wb_state :  std_logic_vector(3 downto 0);
	SIGNAL channel2_wb_state :  std_logic_vector(3 downto 0);
	SIGNAL channel3_wb_state :  std_logic_vector(3 downto 0);
	SIGNAL channel0_wb_cyc_i_delayed :  std_logic;
	SIGNAL channel1_wb_cyc_i_delayed :  std_logic;
	SIGNAL channel2_wb_cyc_i_delayed :  std_logic;
	SIGNAL channel3_wb_cyc_i_delayed :  std_logic;
	SIGNAL c3_p0_wr_en_delayed :  std_logic;
	SIGNAL c3_p1_wr_en_delayed :  std_logic;
	SIGNAL c3_p2_wr_en_delayed :  std_logic;
	SIGNAL c3_p3_wr_en_delayed :  std_logic;
	



	-- COMPONENT DECLARATIONS (introducing the IPs) --------------------------------

	COMPONENT memco
	PORT(
		c3_sys_clk : IN std_logic;
		c3_sys_rst_n : IN std_logic;
		c3_p0_cmd_clk : IN std_logic;
		c3_p0_cmd_en : IN std_logic;
		c3_p0_cmd_instr : IN std_logic_vector(2 downto 0);
		c3_p0_cmd_bl : IN std_logic_vector(5 downto 0);
		c3_p0_cmd_byte_addr : IN std_logic_vector(29 downto 0);
		c3_p0_wr_clk : IN std_logic;
		c3_p0_wr_en : IN std_logic;
		c3_p0_wr_mask : IN std_logic_vector(3 downto 0);
		c3_p0_wr_data : IN std_logic_vector(31 downto 0);
		c3_p0_rd_clk : IN std_logic;
		c3_p0_rd_en : IN std_logic;
		c3_p1_cmd_clk : IN std_logic;
		c3_p1_cmd_en : IN std_logic;
		c3_p1_cmd_instr : IN std_logic_vector(2 downto 0);
		c3_p1_cmd_bl : IN std_logic_vector(5 downto 0);
		c3_p1_cmd_byte_addr : IN std_logic_vector(29 downto 0);
		c3_p1_wr_clk : IN std_logic;
		c3_p1_wr_en : IN std_logic;
		c3_p1_wr_mask : IN std_logic_vector(3 downto 0);
		c3_p1_wr_data : IN std_logic_vector(31 downto 0);
		c3_p1_rd_clk : IN std_logic;
		c3_p1_rd_en : IN std_logic;
		c3_p2_cmd_clk : IN std_logic;
		c3_p2_cmd_en : IN std_logic;
		c3_p2_cmd_instr : IN std_logic_vector(2 downto 0);
		c3_p2_cmd_bl : IN std_logic_vector(5 downto 0);
		c3_p2_cmd_byte_addr : IN std_logic_vector(29 downto 0);
		c3_p2_wr_clk : IN std_logic;
		c3_p2_wr_en : IN std_logic;
		c3_p2_wr_mask : IN std_logic_vector(3 downto 0);
		c3_p2_wr_data : IN std_logic_vector(31 downto 0);
		c3_p2_rd_clk : IN std_logic;
		c3_p2_rd_en : IN std_logic;
		c3_p3_cmd_clk : IN std_logic;
		c3_p3_cmd_en : IN std_logic;
		c3_p3_cmd_instr : IN std_logic_vector(2 downto 0);
		c3_p3_cmd_bl : IN std_logic_vector(5 downto 0);
		c3_p3_cmd_byte_addr : IN std_logic_vector(29 downto 0);
		c3_p3_wr_clk : IN std_logic;
		c3_p3_wr_en : IN std_logic;
		c3_p3_wr_mask : IN std_logic_vector(3 downto 0);
		c3_p3_wr_data : IN std_logic_vector(31 downto 0);
		c3_p3_rd_clk : IN std_logic;
		c3_p3_rd_en : IN std_logic;    
		mcb3_dram_dq : INOUT std_logic_vector(15 downto 0);
		mcb3_dram_udqs : INOUT std_logic;
		mcb3_dram_udqs_n : INOUT std_logic;
		mcb3_rzq : INOUT std_logic;
		mcb3_zio : INOUT std_logic;
		mcb3_dram_dqs : INOUT std_logic;
		mcb3_dram_dqs_n : INOUT std_logic;      
		mcb3_dram_a : OUT std_logic_vector(12 downto 0);
		mcb3_dram_ba : OUT std_logic_vector(1 downto 0);
		mcb3_dram_ras_n : OUT std_logic;
		mcb3_dram_cas_n : OUT std_logic;
		mcb3_dram_we_n : OUT std_logic;
		mcb3_dram_odt : OUT std_logic;
		mcb3_dram_cke : OUT std_logic;
		mcb3_dram_dm : OUT std_logic;
		mcb3_dram_udm : OUT std_logic;
		c3_calib_done : OUT std_logic;
		c3_clk0 : OUT std_logic;
		c3_rst0 : OUT std_logic;
		mcb3_dram_ck : OUT std_logic;
		mcb3_dram_ck_n : OUT std_logic;
		c3_p0_cmd_empty : OUT std_logic;
		c3_p0_cmd_full : OUT std_logic;
		c3_p0_wr_full : OUT std_logic;
		c3_p0_wr_empty : OUT std_logic;
		c3_p0_wr_count : OUT std_logic_vector(6 downto 0);
		c3_p0_wr_underrun : OUT std_logic;
		c3_p0_wr_error : OUT std_logic;
		c3_p0_rd_data : OUT std_logic_vector(31 downto 0);
		c3_p0_rd_full : OUT std_logic;
		c3_p0_rd_empty : OUT std_logic;
		c3_p0_rd_count : OUT std_logic_vector(6 downto 0);
		c3_p0_rd_overflow : OUT std_logic;
		c3_p0_rd_error : OUT std_logic;
		c3_p1_cmd_empty : OUT std_logic;
		c3_p1_cmd_full : OUT std_logic;
		c3_p1_wr_full : OUT std_logic;
		c3_p1_wr_empty : OUT std_logic;
		c3_p1_wr_count : OUT std_logic_vector(6 downto 0);
		c3_p1_wr_underrun : OUT std_logic;
		c3_p1_wr_error : OUT std_logic;
		c3_p1_rd_data : OUT std_logic_vector(31 downto 0);
		c3_p1_rd_full : OUT std_logic;
		c3_p1_rd_empty : OUT std_logic;
		c3_p1_rd_count : OUT std_logic_vector(6 downto 0);
		c3_p1_rd_overflow : OUT std_logic;
		c3_p1_rd_error : OUT std_logic;
		c3_p2_cmd_empty : OUT std_logic;
		c3_p2_cmd_full : OUT std_logic;
		c3_p2_wr_full : OUT std_logic;
		c3_p2_wr_empty : OUT std_logic;
		c3_p2_wr_count : OUT std_logic_vector(6 downto 0);
		c3_p2_wr_underrun : OUT std_logic;
		c3_p2_wr_error : OUT std_logic;
		c3_p2_rd_data : OUT std_logic_vector(31 downto 0);
		c3_p2_rd_full : OUT std_logic;
		c3_p2_rd_empty : OUT std_logic;
		c3_p2_rd_count : OUT std_logic_vector(6 downto 0);
		c3_p2_rd_overflow : OUT std_logic;
		c3_p2_rd_error : OUT std_logic;
		c3_p3_cmd_empty : OUT std_logic;
		c3_p3_cmd_full : OUT std_logic;
		c3_p3_wr_full : OUT std_logic;
		c3_p3_wr_empty : OUT std_logic;
		c3_p3_wr_count : OUT std_logic_vector(6 downto 0);
		c3_p3_wr_underrun : OUT std_logic;
		c3_p3_wr_error : OUT std_logic;
		c3_p3_rd_data : OUT std_logic_vector(31 downto 0);
		c3_p3_rd_full : OUT std_logic;
		c3_p3_rd_empty : OUT std_logic;
		c3_p3_rd_count : OUT std_logic_vector(6 downto 0);
		c3_p3_rd_overflow : OUT std_logic;
		c3_p3_rd_error : OUT std_logic
		);
	END COMPONENT;







---- ------- SYNTHESIS ATTRIBUTES: --------------------------------------------------
--attribute keep_hierarchy : string; 
--attribute keep_hierarchy of s6bfip_memory: entity is "yes"; 






-- --------ARCHITECTURE BODY BEGINS -----------------------------------------------
begin




	-- COMPONENT INSTALLATIONS (connecting the IPs to local signals) ---------------
	

Inst_memco:	memco  PORT MAP(	
	mcb3_dram_dq	=>  mcb3_dram_dq,
	mcb3_dram_a	=>  mcb3_dram_a,
	mcb3_dram_ba	=>  mcb3_dram_ba,
	mcb3_dram_ras_n	=>  mcb3_dram_ras_n,
	mcb3_dram_cas_n	=>  mcb3_dram_cas_n,
	mcb3_dram_we_n	=>  mcb3_dram_we_n,
	mcb3_dram_odt	=>  mcb3_dram_odt,
	mcb3_dram_cke	=>  mcb3_dram_cke,
	mcb3_dram_dm	=>  mcb3_dram_dm,
	mcb3_dram_udqs	=>  mcb3_dram_udqs,
	mcb3_dram_udqs_n	=>  mcb3_dram_udqs_n,
	mcb3_rzq	=>  mcb3_rzq,
	mcb3_zio	=>  mcb3_zio,
	mcb3_dram_udm	=>  mcb3_dram_udm,
	c3_sys_clk	=>  c3_sys_clk,
	c3_sys_rst_n	=>  c3_sys_rst_n,
	c3_calib_done	=>  c3_calib_done,
	c3_clk0	=>  c3_clk0,
	c3_rst0	=>  c3_rst0,
	mcb3_dram_dqs	=>  mcb3_dram_dqs,
	mcb3_dram_dqs_n	=>  mcb3_dram_dqs_n,
	mcb3_dram_ck	=>  mcb3_dram_ck,
	mcb3_dram_ck_n	=>  mcb3_dram_ck_n,
	c3_p0_cmd_clk	=>  c3_p0_cmd_clk,
	c3_p0_cmd_en	=>  c3_p0_cmd_en,
	c3_p0_cmd_instr	=>  c3_p0_cmd_instr,
	c3_p0_cmd_bl	=>  c3_p0_cmd_bl,
	c3_p0_cmd_byte_addr	=>  c3_p0_cmd_byte_addr,
	c3_p0_cmd_empty	=>  c3_p0_cmd_empty,
	c3_p0_cmd_full	=>  c3_p0_cmd_full,
	c3_p0_wr_clk	=>  c3_p0_wr_clk,
	c3_p0_wr_en	=>  c3_p0_wr_en,
	c3_p0_wr_mask	=>  c3_p0_wr_mask,
	c3_p0_wr_data	=>  c3_p0_wr_data,
	c3_p0_wr_full	=>  c3_p0_wr_full,
	c3_p0_wr_empty	=>  c3_p0_wr_empty,
	c3_p0_wr_count	=>  c3_p0_wr_count,
	c3_p0_wr_underrun	=>  c3_p0_wr_underrun,
	c3_p0_wr_error	=>  c3_p0_wr_error,
	c3_p0_rd_clk	=>  c3_p0_rd_clk,
	c3_p0_rd_en	=>  c3_p0_rd_en,
	c3_p0_rd_data	=>  c3_p0_rd_data,
	c3_p0_rd_full	=>  c3_p0_rd_full,
	c3_p0_rd_empty	=>  c3_p0_rd_empty,
	c3_p0_rd_count	=>  c3_p0_rd_count,
	c3_p0_rd_overflow	=>  c3_p0_rd_overflow,
	c3_p0_rd_error	=>  c3_p0_rd_error,
	c3_p1_cmd_clk	=>  c3_p1_cmd_clk,
	c3_p1_cmd_en	=>  c3_p1_cmd_en,
	c3_p1_cmd_instr	=>  c3_p1_cmd_instr,
	c3_p1_cmd_bl	=>  c3_p1_cmd_bl,
	c3_p1_cmd_byte_addr	=>  c3_p1_cmd_byte_addr,
	c3_p1_cmd_empty	=>  c3_p1_cmd_empty,
	c3_p1_cmd_full	=>  c3_p1_cmd_full,
	c3_p1_wr_clk	=>  c3_p1_wr_clk,
	c3_p1_wr_en	=>  c3_p1_wr_en,
	c3_p1_wr_mask	=>  c3_p1_wr_mask,
	c3_p1_wr_data	=>  c3_p1_wr_data,
	c3_p1_wr_full	=>  c3_p1_wr_full,
	c3_p1_wr_empty	=>  c3_p1_wr_empty,
	c3_p1_wr_count	=>  c3_p1_wr_count,
	c3_p1_wr_underrun	=>  c3_p1_wr_underrun,
	c3_p1_wr_error	=>  c3_p1_wr_error,
	c3_p1_rd_clk	=>  c3_p1_rd_clk,
	c3_p1_rd_en	=>  c3_p1_rd_en,
	c3_p1_rd_data	=>  c3_p1_rd_data,
	c3_p1_rd_full	=>  c3_p1_rd_full,
	c3_p1_rd_empty	=>  c3_p1_rd_empty,
	c3_p1_rd_count	=>  c3_p1_rd_count,
	c3_p1_rd_overflow	=>  c3_p1_rd_overflow,
	c3_p1_rd_error	=>  c3_p1_rd_error,
	c3_p2_cmd_clk	=>  c3_p2_cmd_clk,
	c3_p2_cmd_en	=>  c3_p2_cmd_en,
	c3_p2_cmd_instr	=>  c3_p2_cmd_instr,
	c3_p2_cmd_bl	=>  c3_p2_cmd_bl,
	c3_p2_cmd_byte_addr	=>  c3_p2_cmd_byte_addr,
	c3_p2_cmd_empty	=>  c3_p2_cmd_empty,
	c3_p2_cmd_full	=>  c3_p2_cmd_full,
	c3_p2_wr_clk	=>  c3_p2_wr_clk,
	c3_p2_wr_en	=>  c3_p2_wr_en,
	c3_p2_wr_mask	=>  c3_p2_wr_mask,
	c3_p2_wr_data	=>  c3_p2_wr_data,
	c3_p2_wr_full	=>  c3_p2_wr_full,
	c3_p2_wr_empty	=>  c3_p2_wr_empty,
	c3_p2_wr_count	=>  c3_p2_wr_count,
	c3_p2_wr_underrun	=>  c3_p2_wr_underrun,
	c3_p2_wr_error	=>  c3_p2_wr_error,
	c3_p2_rd_clk	=>  c3_p2_rd_clk,
	c3_p2_rd_en	=>  c3_p2_rd_en,
	c3_p2_rd_data	=>  c3_p2_rd_data,
	c3_p2_rd_full	=>  c3_p2_rd_full,
	c3_p2_rd_empty	=>  c3_p2_rd_empty,
	c3_p2_rd_count	=>  c3_p2_rd_count,
	c3_p2_rd_overflow	=>  c3_p2_rd_overflow,
	c3_p2_rd_error	=>  c3_p2_rd_error,
	c3_p3_cmd_clk	=>  c3_p3_cmd_clk,
	c3_p3_cmd_en	=>  c3_p3_cmd_en,
	c3_p3_cmd_instr	=>  c3_p3_cmd_instr,
	c3_p3_cmd_bl	=>  c3_p3_cmd_bl,
	c3_p3_cmd_byte_addr	=>  c3_p3_cmd_byte_addr,
	c3_p3_cmd_empty	=>  c3_p3_cmd_empty,
	c3_p3_cmd_full	=>  c3_p3_cmd_full,
	c3_p3_wr_clk	=>  c3_p3_wr_clk,
	c3_p3_wr_en	=>  c3_p3_wr_en,
	c3_p3_wr_mask	=>  c3_p3_wr_mask,
	c3_p3_wr_data	=>  c3_p3_wr_data,
	c3_p3_wr_full	=>  c3_p3_wr_full,
	c3_p3_wr_empty	=>  c3_p3_wr_empty,
	c3_p3_wr_count	=>  c3_p3_wr_count,
	c3_p3_wr_underrun	=>  c3_p3_wr_underrun,
	c3_p3_wr_error	=>  c3_p3_wr_error,
	c3_p3_rd_clk	=>  c3_p3_rd_clk,
	c3_p3_rd_en	=>  c3_p3_rd_en,
	c3_p3_rd_data	=>  c3_p3_rd_data,
	c3_p3_rd_full	=>  c3_p3_rd_full,
	c3_p3_rd_empty	=>  c3_p3_rd_empty,
	c3_p3_rd_count	=>  c3_p3_rd_count,
	c3_p3_rd_overflow	=>  c3_p3_rd_overflow,
	c3_p3_rd_error	=>  c3_p3_rd_error  
	);  






	-- MAIN LOGIC: -----------------------------------------------------------------

	c3_sys_clk <= x25m_clk;
	c3_sys_rst_n <= reset;

	--unused ports on mem controller: 
	-- <= c3_clk0;
	-- <= c3_rst0;
	-- <= c3_calib_done;



	-- Statemachine / GlueLogic for the PORT-0.--------------------------------
	--This is the glue between the wishbone bus and the Memco-IP.
    process (reset, channel0_wb_clk_i, channel0_wb_cyc_i, channel0_wb_state,
				channel0_wb_wr_i, c3_p0_cmd_full, c3_p0_wr_full, c3_p0_rd_data, c3_p0_cmd_full, c3_p0_wr_full,
				c3_p0_rd_empty, c3_p0_wr_en_delayed, c3_p0_wr_en) 
    begin
    if (reset='1') then 
       channel0_wb_state (3 downto 0) <= "0000";
		 channel0_wb_ack_o <= '0';
		 c3_p0_rd_en <= '0';
		 channel0_wb_data_o <= (OTHERS => '0');
    else
      if (channel0_wb_clk_i'event and channel0_wb_clk_i = '1') then
		
           --generating the delayed wb_cyc value
			  channel0_wb_cyc_i_delayed <= channel0_wb_cyc_i;
			  c3_p0_wr_en_delayed <= c3_p0_wr_en;
					 
			  --State machine:
			  case ( channel0_wb_state ) is

					 --********** IDLE STATE  **********
                when "0000" =>   --state 0        
                    if (channel0_wb_cyc_i ='1' and channel0_wb_wr_i='1' and  c3_p0_cmd_full='0' and c3_p0_wr_full='0') then --write
						    channel0_wb_state <= "0001";
							 c3_p0_wr_en <= '1'; --data is already valid, latch it
						  elsif (channel0_wb_cyc_i ='1' and channel0_wb_wr_i='0' and c3_p0_cmd_full='0') then --read
						    channel0_wb_state <= "0010";
							 c3_p0_cmd_en <= '1';
						  end if;
						  channel0_wb_ack_o <= '0';
						  c3_p0_rd_en <= '0';

                --********** Write STATE ********** 
                when "0001" =>   --state 1
                    if (c3_p0_wr_en='0' and c3_p0_wr_en_delayed='0') then --2clk delay
						    c3_p0_cmd_en <= '1';
							 channel0_wb_state <= "0011"; 
						  end if;
						  c3_p0_wr_en <= '0';
                --* Write complete *
                when "0011" =>   --state 3
                    c3_p0_cmd_en <= '0';
						  channel0_wb_ack_o <= '1';
						  channel0_wb_state <= "0100";  --back to idle
					  
                --********** Read STATE **********     				 
                when "0010" =>   --state 2
                    c3_p0_cmd_en <= '0';
						  if (c3_p0_rd_empty='0') then --if RD FIFO has read data returned
						    c3_p0_rd_en <= '1';
							 channel0_wb_state <= "0100"; --to idle
							 channel0_wb_data_o <= c3_p0_rd_data; --latch and hold the data
							 channel0_wb_ack_o <= '1'; --signal acknowledge for one clk
						  end if;

                --********** "wait for end of wb cycle" STATE **********
                when "0100" =>   --state 4
                    channel0_wb_state <= "0000"; --to idle
						  channel0_wb_ack_o <= '0';
						  c3_p0_rd_en <= '0';
						  
                when others => --error
                      channel0_wb_state <= "0000"; --back to idle
							 
            end case;  
				
       end if; --clocking       
    end if; --reset/non-reset
    end process;
	 
	 --Asynchronous (non-delayed) assigments:
	 c3_p0_rd_clk <= channel0_wb_clk_i;
	 c3_p0_wr_clk <= channel0_wb_clk_i;
	 c3_p0_cmd_clk <= channel0_wb_clk_i;
	 c3_p0_cmd_byte_addr(29 downto 26) <= "0000";
	 c3_p0_cmd_byte_addr(25 downto 2) <= channel0_wb_addr_i (25 downto 2);
	 c3_p0_cmd_byte_addr(1 downto 0) <= "00";
	 c3_p0_cmd_instr (2 downto 1) <= "00";
	 c3_p0_cmd_instr (0) <= not channel0_wb_wr_i;
	 c3_p0_cmd_bl (5 downto 0) <= "000000"; --always single accesses, no multy-dw bursts.
	 c3_p0_wr_data <= channel0_wb_data_i; 
	 c3_p0_wr_mask(0) <= not channel0_wb_sel_i(0);
	 c3_p0_wr_mask(1) <= not channel0_wb_sel_i(1);
	 c3_p0_wr_mask(2) <= not channel0_wb_sel_i(2);
	 c3_p0_wr_mask(3) <= not channel0_wb_sel_i(3);
	 







	-- Statemachine / GlueLogic for the PORT-1.--------------------------------
	--This is the glue between the wishbone bus and the Memco-IP.
    process (reset, channel1_wb_clk_i, channel1_wb_cyc_i, channel1_wb_state,
				channel1_wb_wr_i, c3_p1_cmd_full, c3_p1_wr_full, c3_p1_rd_data,  c3_p1_cmd_full, c3_p1_wr_full,
				c3_p1_rd_empty, c3_p1_wr_en_delayed, c3_p1_wr_en) 
    begin
    if (reset='1') then 
       channel1_wb_state (3 downto 0) <= "0000";
		 channel1_wb_ack_o <= '0';
		 c3_p1_rd_en <= '0';
		 channel1_wb_data_o <= (OTHERS => '0');
    else
      if (channel1_wb_clk_i'event and channel1_wb_clk_i = '1') then
		
           --generating the delayed wb_cyc value
			  channel1_wb_cyc_i_delayed <= channel1_wb_cyc_i;
			  c3_p1_wr_en_delayed <= c3_p1_wr_en;
					 
			  --State machine:
			  case ( channel1_wb_state ) is

					 --********** IDLE STATE  **********
                when "0000" =>   --state 0        
                    if (channel1_wb_cyc_i ='1' and channel1_wb_wr_i='1' and  c3_p1_cmd_full='0' and c3_p1_wr_full='0') then --write
						    channel1_wb_state <= "0001";
							 c3_p1_wr_en <= '1'; --data is already valid, latch it
						  elsif (channel1_wb_cyc_i ='1' and channel1_wb_wr_i='0' and c3_p1_cmd_full='0') then --read
						    channel1_wb_state <= "0010";
							 c3_p1_cmd_en <= '1';
						  end if;
						  channel1_wb_ack_o <= '0';
						  c3_p1_rd_en <= '0';

                --********** Write STATE ********** 
                when "0001" =>   --state 1
                    if (c3_p1_wr_en='0' and c3_p1_wr_en_delayed='0') then --2clk delay
						    c3_p1_cmd_en <= '1';
							 channel1_wb_state <= "0011"; 
						  end if;
						  c3_p1_wr_en <= '0';
                --* Write complete *
                when "0011" =>   --state 3
                    c3_p1_cmd_en <= '0';
						  channel1_wb_ack_o <= '1';
						  channel1_wb_state <= "0100";  --back to idle
					  
                --********** Read STATE **********     				 
                when "0010" =>   --state 2
                    c3_p1_cmd_en <= '0';
						  if (c3_p1_rd_empty='0') then --if RD FIFO has read data returned
						    c3_p1_rd_en <= '1';
							 channel1_wb_state <= "0100"; --back to idle
							 channel1_wb_data_o <= c3_p1_rd_data; --latch and hold the data
							 channel1_wb_ack_o <= '1'; --signal acknowledge for one clk
						  end if;

                --********** "wait for end of wb cycle" STATE **********
                when "0100" =>   --state 4
                    channel1_wb_state <= "0000"; --to idle
						  channel1_wb_ack_o <= '0';
						  c3_p1_rd_en <= '0';
						  
                when others => --error
                      channel1_wb_state <= "0000"; --back to idle
            end case;  
				
       end if; --clocking       
    end if; --reset/non-reset
    end process;
	 
	 --Asynchronous (non-delayed) assigments:
	 c3_p1_rd_clk <= channel1_wb_clk_i;
	 c3_p1_wr_clk <= channel1_wb_clk_i;
	 c3_p1_cmd_clk <= channel1_wb_clk_i;
	 c3_p1_cmd_byte_addr(29 downto 26) <= "0000";
	 c3_p1_cmd_byte_addr(25 downto 2) <= channel1_wb_addr_i (25 downto 2);
	 c3_p1_cmd_byte_addr(1 downto 0) <= "00";
	 c3_p1_cmd_instr (2 downto 1) <= "00";
	 c3_p1_cmd_instr (0) <= not channel1_wb_wr_i;
	 c3_p1_cmd_bl (5 downto 0) <= "000000"; --always single accesses, no multy-dw bursts.
	 c3_p1_wr_data <= channel1_wb_data_i; 
	 c3_p1_wr_mask(0) <= not channel1_wb_sel_i(0);
	 c3_p1_wr_mask(1) <= not channel1_wb_sel_i(1);
	 c3_p1_wr_mask(2) <= not channel1_wb_sel_i(2);
	 c3_p1_wr_mask(3) <= not channel1_wb_sel_i(3);










	-- Statemachine / GlueLogic for the PORT-2.--------------------------------
	--This is the glue between the wishbone bus and the Memco-IP.
    process (reset, channel2_wb_clk_i, channel2_wb_cyc_i, channel2_wb_state,
				channel2_wb_wr_i, c3_p2_cmd_full, c3_p2_wr_full, c3_p2_rd_data, c3_p2_cmd_full, c3_p2_wr_full,
				c3_p2_rd_empty, c3_p2_wr_en_delayed, c3_p2_wr_en) 
    begin
    if (reset='1') then 
       channel2_wb_state (3 downto 0) <= "0000";
		 channel2_wb_ack_o <= '0';
		 c3_p2_rd_en <= '0';
		 channel2_wb_data_o <= (OTHERS => '0');
    else
      if (channel2_wb_clk_i'event and channel2_wb_clk_i = '1') then
		
           --generating the delayed wb_cyc value
			  channel2_wb_cyc_i_delayed <= channel2_wb_cyc_i;
			  c3_p2_wr_en_delayed <= c3_p2_wr_en;
					 
			  --State machine:
			  case ( channel2_wb_state ) is

					 --********** IDLE STATE  **********
                when "0000" =>   --state 0        
                    if (channel2_wb_cyc_i ='1' and channel2_wb_wr_i='1' and  c3_p2_cmd_full='0' and c3_p2_wr_full='0') then --write
						    channel2_wb_state <= "0001";
							 c3_p2_wr_en <= '1'; --data is already valid, latch it
						  elsif (channel2_wb_cyc_i ='1' and channel2_wb_wr_i='0' and c3_p2_cmd_full='0') then --read
						    channel2_wb_state <= "0010";
							 c3_p2_cmd_en <= '1';
						  end if;
						  channel2_wb_ack_o <= '0';
						  c3_p2_rd_en <= '0';

                --********** Write STATE ********** 
                when "0001" =>   --state 1
                    if (c3_p2_wr_en='0' and c3_p2_wr_en_delayed='0') then --2clk delay
						    c3_p2_cmd_en <= '1';
							 channel2_wb_state <= "0011"; 
						  end if;
						  c3_p2_wr_en <= '0';
                --* Write complete *
                when "0011" =>   --state 3
                    c3_p2_cmd_en <= '0';
						  channel2_wb_ack_o <= '1';
						  channel2_wb_state <= "0100";  --back to idle
					  
                --********** Read STATE **********     				 
                when "0010" =>   --state 2
                    c3_p2_cmd_en <= '0';
						  if (c3_p2_rd_empty='0') then --if RD FIFO has read data returned
						    c3_p2_rd_en <= '1';
							 channel2_wb_state <= "0100"; --to idle
							 channel2_wb_data_o <= c3_p2_rd_data; --latch and hold the data
							 channel2_wb_ack_o <= '1'; --signal acknowledge for one clk
						  end if;

                --********** "wait for end of wb cycle" STATE **********
                when "0100" =>   --state 4
                    channel2_wb_state <= "0000"; --to idle
						  channel2_wb_ack_o <= '0';
						  c3_p2_rd_en <= '0';

                when others => --error
                      channel2_wb_state <= "0000"; --back to idle
            end case;  
				
       end if; --clocking       
    end if; --reset/non-reset
    end process;
	 
	 --Asynchronous (non-delayed) assigments:
	 c3_p2_rd_clk <= channel2_wb_clk_i;
	 c3_p2_wr_clk <= channel2_wb_clk_i;
	 c3_p2_cmd_clk <= channel2_wb_clk_i;
	 c3_p2_cmd_byte_addr(29 downto 26) <= "0000";
	 c3_p2_cmd_byte_addr(25 downto 2) <= channel2_wb_addr_i (25 downto 2);
	 c3_p2_cmd_byte_addr(1 downto 0) <= "00";
	 c3_p2_cmd_instr (2 downto 1) <= "00";
	 c3_p2_cmd_instr (0) <= not channel2_wb_wr_i;
	 c3_p2_cmd_bl (5 downto 0) <= "000000"; --always single accesses, no multy-dw bursts.
	 c3_p2_wr_data <= channel2_wb_data_i; 
	 c3_p2_wr_mask(0) <= not channel2_wb_sel_i(0);
	 c3_p2_wr_mask(1) <= not channel2_wb_sel_i(1);
	 c3_p2_wr_mask(2) <= not channel2_wb_sel_i(2);
	 c3_p2_wr_mask(3) <= not channel2_wb_sel_i(3);











	-- Statemachine / GlueLogic for the PORT-3.--------------------------------
	--This is the glue between the wishbone bus and the Memco-IP.
    process (reset, channel3_wb_clk_i, channel3_wb_cyc_i, channel3_wb_state,
				channel3_wb_wr_i, c3_p3_cmd_full, c3_p3_wr_full, c3_p3_rd_data, c3_p3_cmd_full, c3_p3_wr_full,
				c3_p3_rd_empty, c3_p3_wr_en_delayed, c3_p3_wr_en) 
    begin
    if (reset='1') then 
       channel3_wb_state (3 downto 0) <= "0000";
		 channel3_wb_ack_o <= '0';
		 c3_p3_rd_en <= '0';
		 channel3_wb_data_o <= (OTHERS => '0');
    else
      if (channel3_wb_clk_i'event and channel3_wb_clk_i = '1') then
		
           --generating the delayed wb_cyc value
			  channel3_wb_cyc_i_delayed <= channel3_wb_cyc_i;
			  c3_p3_wr_en_delayed <= c3_p3_wr_en;
					 
			  --State machine:
			  case ( channel3_wb_state ) is

					 --********** IDLE STATE  **********
                when "0000" =>   --state 0        
                    if (channel3_wb_cyc_i ='1' and channel3_wb_wr_i='1' and  c3_p3_cmd_full='0' and c3_p3_wr_full='0') then --write
						    channel3_wb_state <= "0001";
							 c3_p3_wr_en <= '1'; --data is already valid, latch it
						  elsif (channel3_wb_cyc_i ='1' and channel3_wb_wr_i='0' and c3_p3_cmd_full='0') then --read
						    channel3_wb_state <= "0010";
							 c3_p3_cmd_en <= '1';
						  end if;
						  channel3_wb_ack_o <= '0';
						  c3_p3_rd_en <= '0';

                --********** Write STATE ********** 
                when "0001" =>   --state 1
                    if (c3_p3_wr_en='0' and c3_p3_wr_en_delayed='0') then --2clk delay
						    c3_p3_cmd_en <= '1';
							 channel3_wb_state <= "0011"; 
						  end if;
						  c3_p3_wr_en <= '0';
                --* Write complete *
                when "0011" =>   --state 3
                    c3_p3_cmd_en <= '0';
						  channel3_wb_ack_o <= '1';
						  channel3_wb_state <= "0100";  --back to idle
					  
                --********** Read STATE **********     				 
                when "0010" =>   --state 2
                    c3_p3_cmd_en <= '0';
						  if (c3_p3_rd_empty='0') then --if RD FIFO has read data returned
						    c3_p3_rd_en <= '1';
							 channel3_wb_state <= "0100"; --to idle
							 channel3_wb_data_o <= c3_p3_rd_data; --latch and hold the data
							 channel3_wb_ack_o <= '1'; --signal acknowledge for one clk
						  end if;

                --********** "wait for end of wb cycle" STATE **********
                when "0100" =>   --state 4
                    channel3_wb_state <= "0000"; --to idle
						  channel3_wb_ack_o <= '0';
						  c3_p3_rd_en <= '0';

                when others => --error
                      channel3_wb_state <= "0000"; --back to idle
            end case;  
				
       end if; --clocking       
    end if; --reset/non-reset
    end process;
	 
	 --Asynchronous (non-delayed) assigments:
	 c3_p3_rd_clk <= channel3_wb_clk_i;
	 c3_p3_wr_clk <= channel3_wb_clk_i;
	 c3_p3_cmd_clk <= channel3_wb_clk_i;
	 c3_p3_cmd_byte_addr(29 downto 26) <= "0000";
	 c3_p3_cmd_byte_addr(25 downto 2) <= channel3_wb_addr_i (25 downto 2);
	 c3_p3_cmd_byte_addr(1 downto 0) <= "00";
	 c3_p3_cmd_instr (2 downto 1) <= "00";
	 c3_p3_cmd_instr (0) <= not channel3_wb_wr_i;
	 c3_p3_cmd_bl (5 downto 0) <= "000000"; --always single accesses, no multy-dw bursts.
	 c3_p3_wr_data <= channel3_wb_data_i; 
	 c3_p3_wr_mask(0) <= not channel3_wb_sel_i(0);
	 c3_p3_wr_mask(1) <= not channel3_wb_sel_i(1);
	 c3_p3_wr_mask(2) <= not channel3_wb_sel_i(2);
	 c3_p3_wr_mask(3) <= not channel3_wb_sel_i(3);














-- -------- END OF FILE -----------------------------------------------------------
end Behavioral;
